
module blink(clk, stdin_valid_in, stdin_in, stdout_ready_in, stdin_ready_out, stdout_valid_out, stdout_out);
  input [0:0] stdin_valid_in;
  input [31:0] stdin_in;
  input [0:0] stdout_ready_in;
  input [0:0] clk;
  output [0:0] stdin_ready_out;
  output [0:0] stdout_valid_out;
  output [31:0] stdout_out;
  wire [0:0] exp_223;
  wire [0:0] exp_206;
  wire [0:0] exp_214;
  wire [0:0] exp_5;
  wire [0:0] exp_228;
  wire [0:0] exp_575;
  wire [0:0] exp_512;
  wire [0:0] exp_377;
  wire [6:0] exp_362;
  wire [31:0] exp_360;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [10:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_242;
  wire [32:0] exp_845;
  wire [0:0] exp_841;
  wire [0:0] exp_537;
  wire [0:0] exp_515;
  wire [0:0] exp_373;
  wire [6:0] exp_372;
  wire [0:0] exp_375;
  wire [6:0] exp_374;
  wire [0:0] exp_536;
  wire [0:0] exp_381;
  wire [6:0] exp_380;
  wire [0:0] exp_535;
  wire [0:0] exp_534;
  wire [0:0] exp_533;
  wire [2:0] exp_363;
  wire [0:0] exp_532;
  wire [0:0] exp_516;
  wire [31:0] exp_352;
  wire [31:0] exp_290;
  wire [0:0] exp_286;
  wire [4:0] exp_266;
  wire [0:0] exp_285;
  wire [0:0] exp_289;
  wire [31:0] exp_282;
  wire [0:0] exp_263;
  wire [0:0] exp_836;
  wire [0:0] exp_835;
  wire [0:0] exp_834;
  wire [0:0] exp_833;
  wire [4:0] exp_245;
  wire [4:0] exp_828;
  wire [0:0] exp_827;
  wire [0:0] exp_419;
  wire [0:0] exp_418;
  wire [0:0] exp_417;
  wire [0:0] exp_416;
  wire [0:0] exp_415;
  wire [0:0] exp_414;
  wire [0:0] exp_365;
  wire [4:0] exp_364;
  wire [0:0] exp_367;
  wire [5:0] exp_366;
  wire [0:0] exp_369;
  wire [5:0] exp_368;
  wire [0:0] exp_371;
  wire [4:0] exp_370;
  wire [0:0] exp_822;
  wire [0:0] exp_821;
  wire [0:0] exp_607;
  wire [0:0] exp_581;
  wire [0:0] exp_579;
  wire [6:0] exp_577;
  wire [5:0] exp_578;
  wire [0:0] exp_580;
  wire [0:0] exp_606;
  wire [2:0] exp_576;
  wire [0:0] exp_820;
  wire [0:0] exp_818;
  wire [0:0] exp_811;
  wire [2:0] exp_726;
  wire [2:0] exp_733;
  wire [0:0] exp_728;
  wire [2:0] exp_727;
  wire [0:0] exp_732;
  wire [2:0] exp_730;
  wire [0:0] exp_729;
  wire [0:0] exp_731;
  wire [0:0] exp_722;
  wire [0:0] exp_721;
  wire [0:0] exp_720;
  wire [2:0] exp_810;
  wire [0:0] exp_819;
  wire [0:0] exp_629;
  wire [5:0] exp_613;
  wire [5:0] exp_620;
  wire [0:0] exp_615;
  wire [5:0] exp_614;
  wire [0:0] exp_619;
  wire [5:0] exp_617;
  wire [0:0] exp_616;
  wire [0:0] exp_618;
  wire [5:0] exp_628;
  wire [0:0] exp_240;
  wire [0:0] exp_239;
  wire [0:0] exp_237;
  wire [0:0] exp_236;
  wire [0:0] exp_234;
  wire [0:0] exp_235;
  wire [0:0] exp_233;
  wire [0:0] exp_846;
  wire [0:0] exp_232;
  wire [0:0] exp_231;
  wire [0:0] exp_850;
  wire [0:0] exp_849;
  wire [0:0] exp_848;
  wire [0:0] exp_847;
  wire [0:0] exp_227;
  wire [0:0] exp_218;
  wire [0:0] exp_213;
  wire [0:0] exp_210;
  wire [31:0] exp_1;
  wire [31:0] exp_224;
  wire [31:0] exp_431;
  wire [31:0] exp_430;
  wire [31:0] exp_429;
  wire [31:0] exp_428;
  wire [11:0] exp_427;
  wire [11:0] exp_426;
  wire [11:0] exp_425;
  wire [0:0] exp_379;
  wire [5:0] exp_378;
  wire [0:0] exp_424;
  wire [11:0] exp_420;
  wire [11:0] exp_423;
  wire [6:0] exp_421;
  wire [4:0] exp_422;
  wire [31:0] exp_209;
  wire [0:0] exp_212;
  wire [31:0] exp_211;
  wire [0:0] exp_217;
  wire [0:0] exp_196;
  wire [0:0] exp_191;
  wire [0:0] exp_188;
  wire [31:0] exp_187;
  wire [0:0] exp_190;
  wire [31:0] exp_189;
  wire [0:0] exp_195;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [31:0] exp_146;
  wire [0:0] exp_149;
  wire [31:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [12:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_229;
  wire [0:0] exp_514;
  wire [0:0] exp_513;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_176;
  wire [0:0] exp_183;
  wire [0:0] exp_198;
  wire [0:0] exp_205;
  wire [0:0] exp_221;
  wire [0:0] exp_824;
  wire [0:0] exp_823;
  wire [0:0] exp_238;
  wire [0:0] exp_281;
  wire [31:0] exp_253;
  wire [0:0] exp_252;
  wire [1:0] exp_261;
  wire [4:0] exp_248;
  wire [0:0] exp_251;
  wire [0:0] exp_830;
  wire [0:0] exp_829;
  wire [4:0] exp_247;
  wire [31:0] exp_249;
  wire [31:0] exp_826;
  wire [0:0] exp_825;
  wire [31:0] exp_462;
  wire [0:0] exp_461;
  wire [31:0] exp_413;
  wire [2:0] exp_356;
  wire [2:0] exp_347;
  wire [0:0] exp_344;
  wire [0:0] exp_278;
  wire [6:0] exp_268;
  wire [6:0] exp_277;
  wire [0:0] exp_280;
  wire [6:0] exp_279;
  wire [0:0] exp_346;
  wire [2:0] exp_334;
  wire [0:0] exp_276;
  wire [4:0] exp_275;
  wire [0:0] exp_333;
  wire [2:0] exp_321;
  wire [0:0] exp_274;
  wire [5:0] exp_273;
  wire [0:0] exp_320;
  wire [2:0] exp_270;
  wire [0:0] exp_319;
  wire [0:0] exp_332;
  wire [0:0] exp_345;
  wire [0:0] exp_351;
  wire [0:0] exp_412;
  wire [31:0] exp_392;
  wire [0:0] exp_358;
  wire [0:0] exp_350;
  wire [0:0] exp_336;
  wire [0:0] exp_323;
  wire [0:0] exp_309;
  wire [0:0] exp_307;
  wire [0:0] exp_308;
  wire [0:0] exp_272;
  wire [4:0] exp_271;
  wire [0:0] exp_322;
  wire [0:0] exp_335;
  wire [0:0] exp_349;
  wire [0:0] exp_348;
  wire [0:0] exp_391;
  wire [31:0] exp_389;
  wire [31:0] exp_354;
  wire [31:0] exp_340;
  wire [0:0] exp_337;
  wire [0:0] exp_339;
  wire [31:0] exp_329;
  wire [0:0] exp_328;
  wire [31:0] exp_315;
  wire [0:0] exp_314;
  wire [31:0] exp_313;
  wire [31:0] exp_311;
  wire [19:0] exp_310;
  wire [3:0] exp_312;
  wire [31:0] exp_327;
  wire [31:0] exp_325;
  wire [19:0] exp_324;
  wire [3:0] exp_326;
  wire [31:0] exp_338;
  wire [31:0] exp_355;
  wire [31:0] exp_343;
  wire [0:0] exp_341;
  wire [0:0] exp_342;
  wire [31:0] exp_331;
  wire [0:0] exp_330;
  wire [31:0] exp_318;
  wire [0:0] exp_317;
  wire [31:0] exp_302;
  wire [0:0] exp_301;
  wire [31:0] exp_296;
  wire [0:0] exp_292;
  wire [4:0] exp_267;
  wire [0:0] exp_291;
  wire [0:0] exp_295;
  wire [31:0] exp_284;
  wire [0:0] exp_264;
  wire [0:0] exp_840;
  wire [0:0] exp_839;
  wire [0:0] exp_838;
  wire [0:0] exp_837;
  wire [4:0] exp_246;
  wire [0:0] exp_283;
  wire [31:0] exp_260;
  wire [0:0] exp_259;
  wire [1:0] exp_262;
  wire [4:0] exp_255;
  wire [0:0] exp_258;
  wire [0:0] exp_832;
  wire [0:0] exp_831;
  wire [4:0] exp_254;
  wire [31:0] exp_256;
  wire [31:0] exp_265;
  wire [31:0] exp_294;
  wire [0:0] exp_293;
  wire [31:0] exp_300;
  wire [31:0] exp_297;
  wire [31:0] exp_299;
  wire [11:0] exp_298;
  wire [31:0] exp_316;
  wire [31:0] exp_244;
  wire [0:0] exp_243;
  wire [31:0] exp_390;
  wire [31:0] exp_394;
  wire [31:0] exp_393;
  wire [5:0] exp_388;
  wire [5:0] exp_387;
  wire [5:0] exp_386;
  wire [4:0] exp_357;
  wire [4:0] exp_306;
  wire [0:0] exp_305;
  wire [4:0] exp_304;
  wire [4:0] exp_269;
  wire [31:0] exp_410;
  wire [1:0] exp_396;
  wire [0:0] exp_395;
  wire [31:0] exp_411;
  wire [1:0] exp_402;
  wire [0:0] exp_401;
  wire [31:0] exp_398;
  wire [31:0] exp_397;
  wire [31:0] exp_400;
  wire [31:0] exp_399;
  wire [31:0] exp_403;
  wire [31:0] exp_407;
  wire [32:0] exp_406;
  wire [32:0] exp_404;
  wire [0:0] exp_385;
  wire [0:0] exp_359;
  wire [0:0] exp_303;
  wire [0:0] exp_384;
  wire [0:0] exp_383;
  wire [0:0] exp_382;
  wire [32:0] exp_405;
  wire [31:0] exp_408;
  wire [31:0] exp_409;
  wire [31:0] exp_460;
  wire [0:0] exp_459;
  wire [31:0] exp_450;
  wire [7:0] exp_449;
  wire [7:0] exp_448;
  wire [7:0] exp_443;
  wire [1:0] exp_434;
  wire [1:0] exp_433;
  wire [1:0] exp_432;
  wire [0:0] exp_442;
  wire [7:0] exp_438;
  wire [31:0] exp_226;
  wire [31:0] exp_216;
  wire [0:0] exp_215;
  wire [31:0] exp_194;
  wire [0:0] exp_193;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [10:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_230;
  wire [3:0] exp_511;
  wire [0:0] exp_510;
  wire [3:0] exp_498;
  wire [3:0] exp_494;
  wire [1:0] exp_497;
  wire [1:0] exp_496;
  wire [1:0] exp_495;
  wire [3:0] exp_503;
  wire [3:0] exp_499;
  wire [0:0] exp_502;
  wire [0:0] exp_501;
  wire [0:0] exp_500;
  wire [3:0] exp_504;
  wire [3:0] exp_505;
  wire [3:0] exp_506;
  wire [3:0] exp_507;
  wire [3:0] exp_508;
  wire [3:0] exp_509;
  wire [10:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_225;
  wire [31:0] exp_493;
  wire [0:0] exp_492;
  wire [31:0] exp_480;
  wire [0:0] exp_479;
  wire [31:0] exp_466;
  wire [7:0] exp_465;
  wire [7:0] exp_464;
  wire [7:0] exp_463;
  wire [31:0] exp_353;
  wire [31:0] exp_474;
  wire [3:0] exp_473;
  wire [31:0] exp_476;
  wire [4:0] exp_475;
  wire [31:0] exp_478;
  wire [4:0] exp_477;
  wire [31:0] exp_484;
  wire [0:0] exp_437;
  wire [0:0] exp_436;
  wire [0:0] exp_435;
  wire [0:0] exp_483;
  wire [31:0] exp_470;
  wire [15:0] exp_469;
  wire [15:0] exp_468;
  wire [15:0] exp_467;
  wire [31:0] exp_482;
  wire [4:0] exp_481;
  wire [31:0] exp_486;
  wire [31:0] exp_485;
  wire [31:0] exp_472;
  wire [31:0] exp_471;
  wire [31:0] exp_487;
  wire [31:0] exp_488;
  wire [31:0] exp_489;
  wire [31:0] exp_490;
  wire [31:0] exp_491;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [10:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [10:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [10:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [10:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [10:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [10:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [10:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [10:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [10:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [10:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [10:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [10:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_179;
  wire [0:0] exp_177;
  wire [31:0] exp_139;
  wire [0:0] exp_178;
  wire [31:0] exp_157;
  wire [31:0] exp_164;
  wire [0:0] exp_159;
  wire [31:0] exp_158;
  wire [0:0] exp_163;
  wire [31:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [31:0] exp_167;
  wire [31:0] exp_174;
  wire [0:0] exp_169;
  wire [31:0] exp_168;
  wire [0:0] exp_173;
  wire [31:0] exp_171;
  wire [0:0] exp_170;
  wire [0:0] exp_172;
  wire [0:0] exp_166;
  wire [0:0] exp_165;
  wire [31:0] exp_182;
  wire [31:0] exp_201;
  wire [31:0] exp_204;
  wire [31:0] exp_219;
  wire [7:0] exp_439;
  wire [7:0] exp_440;
  wire [7:0] exp_441;
  wire [31:0] exp_453;
  wire [15:0] exp_452;
  wire [15:0] exp_451;
  wire [15:0] exp_447;
  wire [0:0] exp_446;
  wire [15:0] exp_444;
  wire [15:0] exp_445;
  wire [31:0] exp_454;
  wire [31:0] exp_455;
  wire [31:0] exp_456;
  wire [31:0] exp_457;
  wire [31:0] exp_458;
  wire [31:0] exp_817;
  wire [0:0] exp_816;
  wire [31:0] exp_813;
  wire [0:0] exp_584;
  wire [0:0] exp_583;
  wire [0:0] exp_582;
  wire [0:0] exp_812;
  wire [31:0] exp_808;
  wire [63:0] exp_807;
  wire [0:0] exp_804;
  wire [0:0] exp_787;
  wire [0:0] exp_764;
  wire [0:0] exp_761;
  wire [0:0] exp_759;
  wire [0:0] exp_741;
  wire [0:0] exp_740;
  wire [0:0] exp_739;
  wire [31:0] exp_737;
  wire [0:0] exp_736;
  wire [0:0] exp_735;
  wire [0:0] exp_724;
  wire [0:0] exp_723;
  wire [0:0] exp_587;
  wire [0:0] exp_586;
  wire [0:0] exp_585;
  wire [0:0] exp_590;
  wire [0:0] exp_589;
  wire [1:0] exp_588;
  wire [0:0] exp_760;
  wire [0:0] exp_744;
  wire [0:0] exp_743;
  wire [0:0] exp_742;
  wire [31:0] exp_738;
  wire [0:0] exp_725;
  wire [0:0] exp_746;
  wire [0:0] exp_745;
  wire [0:0] exp_766;
  wire [1:0] exp_765;
  wire [0:0] exp_789;
  wire [1:0] exp_788;
  wire [0:0] exp_806;
  wire [63:0] exp_803;
  wire [63:0] exp_802;
  wire [63:0] exp_798;
  wire [63:0] exp_794;
  wire [63:0] exp_790;
  wire [31:0] exp_783;
  wire [31:0] exp_770;
  wire [31:0] exp_768;
  wire [15:0] exp_767;
  wire [31:0] exp_762;
  wire [31:0] exp_752;
  wire [31:0] exp_751;
  wire [31:0] exp_750;
  wire [0:0] exp_747;
  wire [0:0] exp_749;
  wire [31:0] exp_748;
  wire [15:0] exp_769;
  wire [31:0] exp_763;
  wire [31:0] exp_758;
  wire [31:0] exp_757;
  wire [31:0] exp_756;
  wire [0:0] exp_753;
  wire [0:0] exp_755;
  wire [31:0] exp_754;
  wire [63:0] exp_793;
  wire [63:0] exp_791;
  wire [31:0] exp_784;
  wire [31:0] exp_774;
  wire [31:0] exp_772;
  wire [15:0] exp_771;
  wire [15:0] exp_773;
  wire [4:0] exp_792;
  wire [63:0] exp_797;
  wire [63:0] exp_795;
  wire [31:0] exp_785;
  wire [31:0] exp_778;
  wire [31:0] exp_776;
  wire [15:0] exp_775;
  wire [15:0] exp_777;
  wire [4:0] exp_796;
  wire [63:0] exp_801;
  wire [63:0] exp_799;
  wire [31:0] exp_786;
  wire [31:0] exp_782;
  wire [31:0] exp_780;
  wire [15:0] exp_779;
  wire [15:0] exp_781;
  wire [5:0] exp_800;
  wire [63:0] exp_805;
  wire [31:0] exp_809;
  wire [31:0] exp_815;
  wire [0:0] exp_608;
  wire [0:0] exp_814;
  wire [31:0] exp_718;
  wire [31:0] exp_712;
  wire [0:0] exp_708;
  wire [0:0] exp_707;
  wire [31:0] exp_656;
  wire [31:0] exp_653;
  wire [31:0] exp_652;
  wire [31:0] exp_651;
  wire [0:0] exp_648;
  wire [0:0] exp_639;
  wire [0:0] exp_638;
  wire [0:0] exp_637;
  wire [31:0] exp_633;
  wire [0:0] exp_631;
  wire [0:0] exp_630;
  wire [0:0] exp_610;
  wire [0:0] exp_609;
  wire [0:0] exp_650;
  wire [31:0] exp_649;
  wire [0:0] exp_641;
  wire [0:0] exp_640;
  wire [0:0] exp_706;
  wire [0:0] exp_711;
  wire [31:0] exp_699;
  wire [31:0] exp_698;
  wire [31:0] exp_697;
  wire [0:0] exp_694;
  wire [0:0] exp_658;
  wire [0:0] exp_654;
  wire [0:0] exp_636;
  wire [0:0] exp_635;
  wire [0:0] exp_634;
  wire [31:0] exp_632;
  wire [0:0] exp_696;
  wire [31:0] exp_692;
  wire [31:0] exp_662;
  wire [31:0] exp_689;
  wire [0:0] exp_623;
  wire [1:0] exp_622;
  wire [0:0] exp_688;
  wire [31:0] exp_681;
  wire [0:0] exp_671;
  wire [0:0] exp_670;
  wire [32:0] exp_669;
  wire [32:0] exp_668;
  wire [32:0] exp_667;
  wire [31:0] exp_665;
  wire [31:0] exp_660;
  wire [32:0] exp_686;
  wire [0:0] exp_685;
  wire [32:0] exp_673;
  wire [0:0] exp_672;
  wire [0:0] exp_684;
  wire [0:0] exp_659;
  wire [0:0] exp_666;
  wire [31:0] exp_664;
  wire [31:0] exp_691;
  wire [0:0] exp_690;
  wire [31:0] exp_683;
  wire [0:0] exp_682;
  wire [31:0] exp_655;
  wire [31:0] exp_647;
  wire [31:0] exp_646;
  wire [31:0] exp_645;
  wire [0:0] exp_642;
  wire [0:0] exp_644;
  wire [31:0] exp_643;
  wire [0:0] exp_663;
  wire [0:0] exp_680;
  wire [31:0] exp_675;
  wire [0:0] exp_674;
  wire [31:0] exp_679;
  wire [31:0] exp_677;
  wire [0:0] exp_676;
  wire [0:0] exp_678;
  wire [0:0] exp_687;
  wire [0:0] exp_661;
  wire [0:0] exp_625;
  wire [5:0] exp_624;
  wire [31:0] exp_695;
  wire [31:0] exp_710;
  wire [0:0] exp_709;
  wire [0:0] exp_627;
  wire [5:0] exp_626;
  wire [31:0] exp_719;
  wire [31:0] exp_717;
  wire [0:0] exp_715;
  wire [0:0] exp_714;
  wire [0:0] exp_713;
  wire [0:0] exp_716;
  wire [31:0] exp_705;
  wire [31:0] exp_704;
  wire [31:0] exp_703;
  wire [0:0] exp_700;
  wire [0:0] exp_657;
  wire [0:0] exp_702;
  wire [31:0] exp_693;
  wire [31:0] exp_701;
  wire [31:0] exp_288;
  wire [0:0] exp_287;
  wire [0:0] exp_517;
  wire [0:0] exp_530;
  wire [0:0] exp_531;
  wire [0:0] exp_518;
  wire [0:0] exp_519;
  wire [0:0] exp_524;
  wire [31:0] exp_521;
  wire [31:0] exp_520;
  wire [31:0] exp_523;
  wire [31:0] exp_522;
  wire [0:0] exp_529;
  wire [31:0] exp_526;
  wire [31:0] exp_525;
  wire [31:0] exp_528;
  wire [31:0] exp_527;
  wire [0:0] exp_844;
  wire [31:0] exp_843;
  wire [2:0] exp_842;
  wire [32:0] exp_574;
  wire [0:0] exp_573;
  wire [31:0] exp_564;
  wire [31:0] exp_563;
  wire [0:0] exp_562;
  wire [31:0] exp_549;
  wire [12:0] exp_548;
  wire [12:0] exp_547;
  wire [12:0] exp_546;
  wire [11:0] exp_545;
  wire [7:0] exp_544;
  wire [1:0] exp_543;
  wire [0:0] exp_538;
  wire [0:0] exp_539;
  wire [5:0] exp_540;
  wire [3:0] exp_541;
  wire [0:0] exp_542;
  wire [31:0] exp_561;
  wire [20:0] exp_560;
  wire [20:0] exp_559;
  wire [20:0] exp_558;
  wire [19:0] exp_557;
  wire [9:0] exp_556;
  wire [8:0] exp_555;
  wire [0:0] exp_550;
  wire [7:0] exp_551;
  wire [0:0] exp_552;
  wire [9:0] exp_553;
  wire [0:0] exp_554;
  wire [31:0] exp_361;
  wire [32:0] exp_572;
  wire [32:0] exp_571;
  wire [31:0] exp_569;
  wire [31:0] exp_568;
  wire [11:0] exp_567;
  wire [11:0] exp_566;
  wire [11:0] exp_565;
  wire [32:0] exp_570;
  wire [0:0] exp_241;
  wire [0:0] exp_80;
  wire [10:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_376;
  wire [0:0] exp_222;
  wire [0:0] exp_207;
  wire [0:0] exp_200;
  wire [0:0] exp_184;
  wire [0:0] exp_192;
  wire [0:0] exp_185;
  wire [31:0] exp_181;

  assign exp_223 = exp_206 & exp_222;
  assign exp_206 = exp_214;
  assign exp_214 = exp_5 & exp_213;
  assign exp_5 = exp_228;
  assign exp_228 = exp_575;
  assign exp_575 = exp_512 & exp_240;
  assign exp_512 = exp_377 | exp_379;
  assign exp_377 = exp_362 == exp_376;
  assign exp_362 = exp_360[6:0];

      reg [31:0] exp_360_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_360_reg <= exp_96;
        end
      end
      assign exp_360 = exp_360_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_242;

      reg [31:0] exp_242_reg = 0;
      always@(posedge clk) begin
        if (exp_241) begin
          exp_242_reg <= exp_845;
        end
      end
      assign exp_242 = exp_242_reg;
    
  reg [32:0] exp_845_reg;
  always@(*) begin
    case (exp_841)
      0:exp_845_reg <= exp_843;
      1:exp_845_reg <= exp_574;
      default:exp_845_reg <= exp_844;
    endcase
  end
  assign exp_845 = exp_845_reg;
  assign exp_841 = exp_537 & exp_240;
  assign exp_537 = exp_515 | exp_536;
  assign exp_515 = exp_373 | exp_375;
  assign exp_373 = exp_362 == exp_372;
  assign exp_372 = 111;
  assign exp_375 = exp_362 == exp_374;
  assign exp_374 = 103;

  reg [0:0] exp_536_reg;
  always@(*) begin
    case (exp_381)
      0:exp_536_reg <= exp_534;
      1:exp_536_reg <= exp_533;
      default:exp_536_reg <= exp_535;
    endcase
  end
  assign exp_536 = exp_536_reg;
  assign exp_381 = exp_362 == exp_380;
  assign exp_380 = 99;
  assign exp_535 = 0;
  assign exp_534 = 0;

  reg [0:0] exp_533_reg;
  always@(*) begin
    case (exp_363)
      0:exp_533_reg <= exp_516;
      1:exp_533_reg <= exp_517;
      2:exp_533_reg <= exp_530;
      3:exp_533_reg <= exp_531;
      4:exp_533_reg <= exp_518;
      5:exp_533_reg <= exp_519;
      6:exp_533_reg <= exp_524;
      7:exp_533_reg <= exp_529;
      default:exp_533_reg <= exp_532;
    endcase
  end
  assign exp_533 = exp_533_reg;
  assign exp_363 = exp_360[14:12];
  assign exp_532 = 0;
  assign exp_516 = exp_352 == exp_353;

      reg [31:0] exp_352_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_352_reg <= exp_290;
        end
      end
      assign exp_352 = exp_352_reg;
    
  reg [31:0] exp_290_reg;
  always@(*) begin
    case (exp_286)
      0:exp_290_reg <= exp_282;
      1:exp_290_reg <= exp_288;
      default:exp_290_reg <= exp_289;
    endcase
  end
  assign exp_290 = exp_290_reg;
  assign exp_286 = exp_266 == exp_285;
  assign exp_266 = exp_96[19:15];
  assign exp_285 = 0;
  assign exp_289 = 0;

  reg [31:0] exp_282_reg;
  always@(*) begin
    case (exp_263)
      0:exp_282_reg <= exp_253;
      1:exp_282_reg <= exp_265;
      default:exp_282_reg <= exp_281;
    endcase
  end
  assign exp_282 = exp_282_reg;
  assign exp_263 = exp_836;
  assign exp_836 = exp_835 & exp_232;
  assign exp_835 = exp_834 & exp_240;
  assign exp_834 = exp_833 & exp_827;
  assign exp_833 = exp_245 == exp_828;
  assign exp_245 = exp_96[19:15];
  assign exp_828 = exp_360[11:7];
  assign exp_827 = exp_419 | exp_822;
  assign exp_419 = exp_418 | exp_377;
  assign exp_418 = exp_417 | exp_371;
  assign exp_417 = exp_416 | exp_369;
  assign exp_416 = exp_415 | exp_375;
  assign exp_415 = exp_414 | exp_373;
  assign exp_414 = exp_365 | exp_367;
  assign exp_365 = exp_362 == exp_364;
  assign exp_364 = 19;
  assign exp_367 = exp_362 == exp_366;
  assign exp_366 = 51;
  assign exp_369 = exp_362 == exp_368;
  assign exp_368 = 55;
  assign exp_371 = exp_362 == exp_370;
  assign exp_370 = 23;
  assign exp_822 = exp_821 & exp_581;

  reg [0:0] exp_821_reg;
  always@(*) begin
    case (exp_607)
      0:exp_821_reg <= exp_818;
      1:exp_821_reg <= exp_819;
      default:exp_821_reg <= exp_820;
    endcase
  end
  assign exp_821 = exp_821_reg;
  assign exp_607 = exp_581 & exp_606;
  assign exp_581 = exp_579 & exp_580;
  assign exp_579 = exp_577 == exp_578;
  assign exp_577 = exp_360[6:0];
  assign exp_578 = 51;
  assign exp_580 = exp_360[25:25];
  assign exp_606 = exp_576[2:2];
  assign exp_576 = exp_360[14:12];
  assign exp_820 = 0;
  assign exp_818 = exp_811 & exp_581;
  assign exp_811 = exp_726 == exp_810;

      reg [2:0] exp_726_reg = 0;
      always@(posedge clk) begin
        if (exp_722) begin
          exp_726_reg <= exp_733;
        end
      end
      assign exp_726 = exp_726_reg;
    
  reg [2:0] exp_733_reg;
  always@(*) begin
    case (exp_728)
      0:exp_733_reg <= exp_730;
      1:exp_733_reg <= exp_731;
      default:exp_733_reg <= exp_732;
    endcase
  end
  assign exp_733 = exp_733_reg;
  assign exp_728 = exp_726 == exp_727;
  assign exp_727 = 4;
  assign exp_732 = 0;
  assign exp_730 = exp_726 + exp_729;
  assign exp_729 = 1;
  assign exp_731 = 0;
  assign exp_722 = exp_581 & exp_721;
  assign exp_721 = ~exp_720;
  assign exp_720 = exp_576[2:2];
  assign exp_810 = 4;
  assign exp_819 = exp_629 & exp_581;
  assign exp_629 = exp_613 == exp_628;

      reg [5:0] exp_613_reg = 0;
      always@(posedge clk) begin
        if (exp_607) begin
          exp_613_reg <= exp_620;
        end
      end
      assign exp_613 = exp_613_reg;
    
  reg [5:0] exp_620_reg;
  always@(*) begin
    case (exp_615)
      0:exp_620_reg <= exp_617;
      1:exp_620_reg <= exp_618;
      default:exp_620_reg <= exp_619;
    endcase
  end
  assign exp_620 = exp_620_reg;
  assign exp_615 = exp_613 == exp_614;
  assign exp_614 = 37;
  assign exp_619 = 0;
  assign exp_617 = exp_613 + exp_616;
  assign exp_616 = 1;
  assign exp_618 = 0;
  assign exp_628 = 37;

      reg [0:0] exp_240_reg = 0;
      always@(posedge clk) begin
        if (exp_232) begin
          exp_240_reg <= exp_239;
        end
      end
      assign exp_240 = exp_240_reg;
      assign exp_239 = exp_237 & exp_238;

      reg [0:0] exp_237_reg = 0;
      always@(posedge clk) begin
        if (exp_232) begin
          exp_237_reg <= exp_236;
        end
      end
      assign exp_237 = exp_237_reg;
      assign exp_236 = exp_234 & exp_235;
  assign exp_234 = 1;
  assign exp_235 = ~exp_233;
  assign exp_233 = exp_846;
  assign exp_846 = exp_240 & exp_537;
  assign exp_232 = ~exp_231;
  assign exp_231 = exp_850;
  assign exp_850 = exp_240 & exp_849;
  assign exp_849 = exp_848 | exp_824;
  assign exp_848 = exp_228 & exp_847;
  assign exp_847 = ~exp_227;
  assign exp_227 = exp_218;

  reg [0:0] exp_218_reg;
  always@(*) begin
    case (exp_213)
      0:exp_218_reg <= exp_196;
      1:exp_218_reg <= exp_205;
      default:exp_218_reg <= exp_217;
    endcase
  end
  assign exp_218 = exp_218_reg;
  assign exp_213 = exp_210 & exp_212;
  assign exp_210 = exp_1 >= exp_209;
  assign exp_1 = exp_224;
  assign exp_224 = exp_431;
  assign exp_431 = exp_430 + exp_429;
  assign exp_430 = 0;
  assign exp_429 = exp_352 + exp_428;
  assign exp_428 = $signed(exp_427);
  assign exp_427 = exp_426 + exp_425;
  assign exp_426 = 0;

  reg [11:0] exp_425_reg;
  always@(*) begin
    case (exp_379)
      0:exp_425_reg <= exp_420;
      1:exp_425_reg <= exp_423;
      default:exp_425_reg <= exp_424;
    endcase
  end
  assign exp_425 = exp_425_reg;
  assign exp_379 = exp_362 == exp_378;
  assign exp_378 = 35;
  assign exp_424 = 0;
  assign exp_420 = exp_360[31:20];
  assign exp_423 = {exp_421, exp_422};  assign exp_421 = exp_360[31:25];
  assign exp_422 = exp_360[11:7];
  assign exp_209 = 2147483664;
  assign exp_212 = exp_1 <= exp_211;
  assign exp_211 = 2147483664;
  assign exp_217 = 0;

  reg [0:0] exp_196_reg;
  always@(*) begin
    case (exp_191)
      0:exp_196_reg <= exp_155;
      1:exp_196_reg <= exp_183;
      default:exp_196_reg <= exp_195;
    endcase
  end
  assign exp_196 = exp_196_reg;
  assign exp_191 = exp_188 & exp_190;
  assign exp_188 = exp_1 >= exp_187;
  assign exp_187 = 2147483656;
  assign exp_190 = exp_1 <= exp_189;
  assign exp_189 = 2147483656;
  assign exp_195 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 2147483648;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 2147483652;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 8188;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_229;
  assign exp_229 = exp_514;
  assign exp_514 = exp_513 + exp_379;
  assign exp_513 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_176;
  assign exp_176 = 1;
  assign exp_183 = exp_198;
  assign exp_198 = stdout_ready_in;
  assign exp_205 = exp_221;
  assign exp_221 = stdin_valid_in;
  assign exp_824 = exp_581 & exp_823;
  assign exp_823 = ~exp_821;
  assign exp_238 = ~exp_233;
  assign exp_281 = 0;

  //Create RAM
  reg [31:0] exp_253_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_251) begin
      exp_253_ram[exp_247] <= exp_249;
    end
  end
  assign exp_253 = exp_253_ram[exp_248];
  assign exp_252 = exp_261;
  assign exp_261 = 1;
  assign exp_248 = exp_245;
  assign exp_251 = exp_830;
  assign exp_830 = exp_829 & exp_232;
  assign exp_829 = exp_827 & exp_240;
  assign exp_247 = exp_828;
  assign exp_249 = exp_826;

  reg [31:0] exp_826_reg;
  always@(*) begin
    case (exp_822)
      0:exp_826_reg <= exp_462;
      1:exp_826_reg <= exp_817;
      default:exp_826_reg <= exp_825;
    endcase
  end
  assign exp_826 = exp_826_reg;
  assign exp_825 = 0;

  reg [31:0] exp_462_reg;
  always@(*) begin
    case (exp_377)
      0:exp_462_reg <= exp_413;
      1:exp_462_reg <= exp_460;
      default:exp_462_reg <= exp_461;
    endcase
  end
  assign exp_462 = exp_462_reg;
  assign exp_461 = 0;

  reg [31:0] exp_413_reg;
  always@(*) begin
    case (exp_356)
      0:exp_413_reg <= exp_392;
      1:exp_413_reg <= exp_394;
      2:exp_413_reg <= exp_410;
      3:exp_413_reg <= exp_411;
      4:exp_413_reg <= exp_403;
      5:exp_413_reg <= exp_407;
      6:exp_413_reg <= exp_408;
      7:exp_413_reg <= exp_409;
      default:exp_413_reg <= exp_412;
    endcase
  end
  assign exp_413 = exp_413_reg;

      reg [2:0] exp_356_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_356_reg <= exp_347;
        end
      end
      assign exp_356 = exp_356_reg;
    
  reg [2:0] exp_347_reg;
  always@(*) begin
    case (exp_344)
      0:exp_347_reg <= exp_334;
      1:exp_347_reg <= exp_345;
      default:exp_347_reg <= exp_346;
    endcase
  end
  assign exp_347 = exp_347_reg;
  assign exp_344 = exp_278 | exp_280;
  assign exp_278 = exp_268 == exp_277;
  assign exp_268 = exp_96[6:0];
  assign exp_277 = 111;
  assign exp_280 = exp_268 == exp_279;
  assign exp_279 = 103;
  assign exp_346 = 0;

  reg [2:0] exp_334_reg;
  always@(*) begin
    case (exp_276)
      0:exp_334_reg <= exp_321;
      1:exp_334_reg <= exp_332;
      default:exp_334_reg <= exp_333;
    endcase
  end
  assign exp_334 = exp_334_reg;
  assign exp_276 = exp_268 == exp_275;
  assign exp_275 = 23;
  assign exp_333 = 0;

  reg [2:0] exp_321_reg;
  always@(*) begin
    case (exp_274)
      0:exp_321_reg <= exp_270;
      1:exp_321_reg <= exp_319;
      default:exp_321_reg <= exp_320;
    endcase
  end
  assign exp_321 = exp_321_reg;
  assign exp_274 = exp_268 == exp_273;
  assign exp_273 = 55;
  assign exp_320 = 0;
  assign exp_270 = exp_96[14:12];
  assign exp_319 = 0;
  assign exp_332 = 0;
  assign exp_345 = 0;
  assign exp_351 = exp_232 & exp_237;
  assign exp_412 = 0;

  reg [31:0] exp_392_reg;
  always@(*) begin
    case (exp_358)
      0:exp_392_reg <= exp_389;
      1:exp_392_reg <= exp_390;
      default:exp_392_reg <= exp_391;
    endcase
  end
  assign exp_392 = exp_392_reg;

      reg [0:0] exp_358_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_358_reg <= exp_350;
        end
      end
      assign exp_358 = exp_358_reg;
      assign exp_350 = exp_336 & exp_349;
  assign exp_336 = exp_323 & exp_335;
  assign exp_323 = exp_309 & exp_322;
  assign exp_309 = exp_307 & exp_308;
  assign exp_307 = exp_96[30:30];
  assign exp_308 = ~exp_272;
  assign exp_272 = exp_268 == exp_271;
  assign exp_271 = 19;
  assign exp_322 = ~exp_274;
  assign exp_335 = ~exp_276;
  assign exp_349 = ~exp_348;
  assign exp_348 = exp_278 | exp_280;
  assign exp_391 = 0;
  assign exp_389 = exp_354 + exp_355;

      reg [31:0] exp_354_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_354_reg <= exp_340;
        end
      end
      assign exp_354 = exp_354_reg;
    
  reg [31:0] exp_340_reg;
  always@(*) begin
    case (exp_337)
      0:exp_340_reg <= exp_329;
      1:exp_340_reg <= exp_338;
      default:exp_340_reg <= exp_339;
    endcase
  end
  assign exp_340 = exp_340_reg;
  assign exp_337 = exp_278 | exp_280;
  assign exp_339 = 0;

  reg [31:0] exp_329_reg;
  always@(*) begin
    case (exp_276)
      0:exp_329_reg <= exp_315;
      1:exp_329_reg <= exp_327;
      default:exp_329_reg <= exp_328;
    endcase
  end
  assign exp_329 = exp_329_reg;
  assign exp_328 = 0;

  reg [31:0] exp_315_reg;
  always@(*) begin
    case (exp_274)
      0:exp_315_reg <= exp_290;
      1:exp_315_reg <= exp_313;
      default:exp_315_reg <= exp_314;
    endcase
  end
  assign exp_315 = exp_315_reg;
  assign exp_314 = 0;
  assign exp_313 = exp_311 << exp_312;
  assign exp_311 = exp_310;
  assign exp_310 = exp_96[31:12];
  assign exp_312 = 12;
  assign exp_327 = exp_325 << exp_326;
  assign exp_325 = exp_324;
  assign exp_324 = exp_96[31:12];
  assign exp_326 = 12;
  assign exp_338 = 4;

      reg [31:0] exp_355_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_355_reg <= exp_343;
        end
      end
      assign exp_355 = exp_355_reg;
    
  reg [31:0] exp_343_reg;
  always@(*) begin
    case (exp_341)
      0:exp_343_reg <= exp_331;
      1:exp_343_reg <= exp_244;
      default:exp_343_reg <= exp_342;
    endcase
  end
  assign exp_343 = exp_343_reg;
  assign exp_341 = exp_278 | exp_280;
  assign exp_342 = 0;

  reg [31:0] exp_331_reg;
  always@(*) begin
    case (exp_276)
      0:exp_331_reg <= exp_318;
      1:exp_331_reg <= exp_244;
      default:exp_331_reg <= exp_330;
    endcase
  end
  assign exp_331 = exp_331_reg;
  assign exp_330 = 0;

  reg [31:0] exp_318_reg;
  always@(*) begin
    case (exp_274)
      0:exp_318_reg <= exp_302;
      1:exp_318_reg <= exp_316;
      default:exp_318_reg <= exp_317;
    endcase
  end
  assign exp_318 = exp_318_reg;
  assign exp_317 = 0;

  reg [31:0] exp_302_reg;
  always@(*) begin
    case (exp_272)
      0:exp_302_reg <= exp_296;
      1:exp_302_reg <= exp_300;
      default:exp_302_reg <= exp_301;
    endcase
  end
  assign exp_302 = exp_302_reg;
  assign exp_301 = 0;

  reg [31:0] exp_296_reg;
  always@(*) begin
    case (exp_292)
      0:exp_296_reg <= exp_284;
      1:exp_296_reg <= exp_294;
      default:exp_296_reg <= exp_295;
    endcase
  end
  assign exp_296 = exp_296_reg;
  assign exp_292 = exp_267 == exp_291;
  assign exp_267 = exp_96[24:20];
  assign exp_291 = 0;
  assign exp_295 = 0;

  reg [31:0] exp_284_reg;
  always@(*) begin
    case (exp_264)
      0:exp_284_reg <= exp_260;
      1:exp_284_reg <= exp_265;
      default:exp_284_reg <= exp_283;
    endcase
  end
  assign exp_284 = exp_284_reg;
  assign exp_264 = exp_840;
  assign exp_840 = exp_839 & exp_232;
  assign exp_839 = exp_838 & exp_240;
  assign exp_838 = exp_837 & exp_827;
  assign exp_837 = exp_246 == exp_828;
  assign exp_246 = exp_96[24:20];
  assign exp_283 = 0;

  //Create RAM
  reg [31:0] exp_260_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_258) begin
      exp_260_ram[exp_254] <= exp_256;
    end
  end
  assign exp_260 = exp_260_ram[exp_255];
  assign exp_259 = exp_262;
  assign exp_262 = 1;
  assign exp_255 = exp_246;
  assign exp_258 = exp_832;
  assign exp_832 = exp_831 & exp_232;
  assign exp_831 = exp_827 & exp_240;
  assign exp_254 = exp_828;
  assign exp_256 = exp_826;
  assign exp_265 = exp_826;
  assign exp_294 = $signed(exp_293);
  assign exp_293 = 0;
  assign exp_300 = exp_297 + exp_299;
  assign exp_297 = 0;
  assign exp_299 = $signed(exp_298);
  assign exp_298 = exp_96[31:20];
  assign exp_316 = 0;

      reg [31:0] exp_244_reg = 0;
      always@(posedge clk) begin
        if (exp_243) begin
          exp_244_reg <= exp_242;
        end
      end
      assign exp_244 = exp_244_reg;
      assign exp_243 = exp_234 & exp_232;
  assign exp_390 = exp_354 - exp_355;
  assign exp_394 = exp_354 << exp_393;
  assign exp_393 = $signed(exp_388);
  assign exp_388 = exp_387 + exp_386;
  assign exp_387 = 0;
  assign exp_386 = exp_357;

      reg [4:0] exp_357_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_357_reg <= exp_306;
        end
      end
      assign exp_357 = exp_357_reg;
    
  reg [4:0] exp_306_reg;
  always@(*) begin
    case (exp_272)
      0:exp_306_reg <= exp_304;
      1:exp_306_reg <= exp_269;
      default:exp_306_reg <= exp_305;
    endcase
  end
  assign exp_306 = exp_306_reg;
  assign exp_305 = 0;
  assign exp_304 = exp_302[4:0];
  assign exp_269 = exp_96[24:20];
  assign exp_410 = $signed(exp_396);
  assign exp_396 = exp_395;
  assign exp_395 = $signed(exp_354) < $signed(exp_355);
  assign exp_411 = $signed(exp_402);
  assign exp_402 = exp_401;
  assign exp_401 = exp_398 < exp_400;
  assign exp_398 = exp_397 + exp_354;
  assign exp_397 = 0;
  assign exp_400 = exp_399 + exp_355;
  assign exp_399 = 0;
  assign exp_403 = exp_354 ^ exp_355;
  assign exp_407 = exp_406[31:0];
  assign exp_406 = $signed(exp_404) >>> $signed(exp_405);
  assign exp_404 = {exp_385, exp_354};
  reg [0:0] exp_385_reg;
  always@(*) begin
    case (exp_359)
      0:exp_385_reg <= exp_383;
      1:exp_385_reg <= exp_382;
      default:exp_385_reg <= exp_384;
    endcase
  end
  assign exp_385 = exp_385_reg;

      reg [0:0] exp_359_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_359_reg <= exp_303;
        end
      end
      assign exp_359 = exp_359_reg;
      assign exp_303 = exp_96[30:30];
  assign exp_384 = 0;
  assign exp_383 = 0;
  assign exp_382 = exp_354[31:31];
  assign exp_405 = $signed(exp_388);
  assign exp_408 = exp_354 | exp_355;
  assign exp_409 = exp_354 & exp_355;

  reg [31:0] exp_460_reg;
  always@(*) begin
    case (exp_363)
      0:exp_460_reg <= exp_450;
      1:exp_460_reg <= exp_453;
      2:exp_460_reg <= exp_226;
      3:exp_460_reg <= exp_454;
      4:exp_460_reg <= exp_455;
      5:exp_460_reg <= exp_456;
      6:exp_460_reg <= exp_457;
      7:exp_460_reg <= exp_458;
      default:exp_460_reg <= exp_459;
    endcase
  end
  assign exp_460 = exp_460_reg;
  assign exp_459 = 0;
  assign exp_450 = $signed(exp_449);
  assign exp_449 = exp_448 + exp_443;
  assign exp_448 = 0;

  reg [7:0] exp_443_reg;
  always@(*) begin
    case (exp_434)
      0:exp_443_reg <= exp_438;
      1:exp_443_reg <= exp_439;
      2:exp_443_reg <= exp_440;
      3:exp_443_reg <= exp_441;
      default:exp_443_reg <= exp_442;
    endcase
  end
  assign exp_443 = exp_443_reg;
  assign exp_434 = exp_433 + exp_432;
  assign exp_433 = 0;
  assign exp_432 = exp_431[1:0];
  assign exp_442 = 0;
  assign exp_438 = exp_226[7:0];
  assign exp_226 = exp_216;

  reg [31:0] exp_216_reg;
  always@(*) begin
    case (exp_213)
      0:exp_216_reg <= exp_194;
      1:exp_216_reg <= exp_204;
      default:exp_216_reg <= exp_215;
    endcase
  end
  assign exp_216 = exp_216_reg;
  assign exp_215 = 0;

  reg [31:0] exp_194_reg;
  always@(*) begin
    case (exp_191)
      0:exp_194_reg <= exp_153;
      1:exp_194_reg <= exp_182;
      default:exp_194_reg <= exp_193;
    endcase
  end
  assign exp_194 = exp_194_reg;
  assign exp_193 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 0;
    exp_54_ram[32] = 252;
    exp_54_ram[33] = 10;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 253;
    exp_54_ram[36] = 2;
    exp_54_ram[37] = 3;
    exp_54_ram[38] = 252;
    exp_54_ram[39] = 252;
    exp_54_ram[40] = 253;
    exp_54_ram[41] = 254;
    exp_54_ram[42] = 253;
    exp_54_ram[43] = 254;
    exp_54_ram[44] = 0;
    exp_54_ram[45] = 253;
    exp_54_ram[46] = 0;
    exp_54_ram[47] = 2;
    exp_54_ram[48] = 3;
    exp_54_ram[49] = 0;
    exp_54_ram[50] = 254;
    exp_54_ram[51] = 0;
    exp_54_ram[52] = 2;
    exp_54_ram[53] = 128;
    exp_54_ram[54] = 254;
    exp_54_ram[55] = 128;
    exp_54_ram[56] = 0;
    exp_54_ram[57] = 254;
    exp_54_ram[58] = 254;
    exp_54_ram[59] = 0;
    exp_54_ram[60] = 0;
    exp_54_ram[61] = 254;
    exp_54_ram[62] = 0;
    exp_54_ram[63] = 0;
    exp_54_ram[64] = 0;
    exp_54_ram[65] = 0;
    exp_54_ram[66] = 0;
    exp_54_ram[67] = 0;
    exp_54_ram[68] = 0;
    exp_54_ram[69] = 0;
    exp_54_ram[70] = 0;
    exp_54_ram[71] = 0;
    exp_54_ram[72] = 1;
    exp_54_ram[73] = 2;
    exp_54_ram[74] = 0;
    exp_54_ram[75] = 252;
    exp_54_ram[76] = 2;
    exp_54_ram[77] = 2;
    exp_54_ram[78] = 3;
    exp_54_ram[79] = 3;
    exp_54_ram[80] = 3;
    exp_54_ram[81] = 3;
    exp_54_ram[82] = 3;
    exp_54_ram[83] = 3;
    exp_54_ram[84] = 1;
    exp_54_ram[85] = 1;
    exp_54_ram[86] = 4;
    exp_54_ram[87] = 246;
    exp_54_ram[88] = 252;
    exp_54_ram[89] = 252;
    exp_54_ram[90] = 0;
    exp_54_ram[91] = 245;
    exp_54_ram[92] = 0;
    exp_54_ram[93] = 0;
    exp_54_ram[94] = 252;
    exp_54_ram[95] = 252;
    exp_54_ram[96] = 64;
    exp_54_ram[97] = 0;
    exp_54_ram[98] = 1;
    exp_54_ram[99] = 64;
    exp_54_ram[100] = 65;
    exp_54_ram[101] = 0;
    exp_54_ram[102] = 42;
    exp_54_ram[103] = 0;
    exp_54_ram[104] = 0;
    exp_54_ram[105] = 0;
    exp_54_ram[106] = 0;
    exp_54_ram[107] = 252;
    exp_54_ram[108] = 0;
    exp_54_ram[109] = 0;
    exp_54_ram[110] = 0;
    exp_54_ram[111] = 0;
    exp_54_ram[112] = 250;
    exp_54_ram[113] = 42;
    exp_54_ram[114] = 0;
    exp_54_ram[115] = 0;
    exp_54_ram[116] = 252;
    exp_54_ram[117] = 252;
    exp_54_ram[118] = 1;
    exp_54_ram[119] = 0;
    exp_54_ram[120] = 0;
    exp_54_ram[121] = 1;
    exp_54_ram[122] = 0;
    exp_54_ram[123] = 0;
    exp_54_ram[124] = 252;
    exp_54_ram[125] = 252;
    exp_54_ram[126] = 43;
    exp_54_ram[127] = 0;
    exp_54_ram[128] = 0;
    exp_54_ram[129] = 232;
    exp_54_ram[130] = 0;
    exp_54_ram[131] = 235;
    exp_54_ram[132] = 0;
    exp_54_ram[133] = 0;
    exp_54_ram[134] = 252;
    exp_54_ram[135] = 252;
    exp_54_ram[136] = 64;
    exp_54_ram[137] = 0;
    exp_54_ram[138] = 1;
    exp_54_ram[139] = 64;
    exp_54_ram[140] = 65;
    exp_54_ram[141] = 0;
    exp_54_ram[142] = 42;
    exp_54_ram[143] = 0;
    exp_54_ram[144] = 0;
    exp_54_ram[145] = 0;
    exp_54_ram[146] = 0;
    exp_54_ram[147] = 252;
    exp_54_ram[148] = 0;
    exp_54_ram[149] = 0;
    exp_54_ram[150] = 0;
    exp_54_ram[151] = 0;
    exp_54_ram[152] = 250;
    exp_54_ram[153] = 42;
    exp_54_ram[154] = 0;
    exp_54_ram[155] = 0;
    exp_54_ram[156] = 252;
    exp_54_ram[157] = 252;
    exp_54_ram[158] = 1;
    exp_54_ram[159] = 0;
    exp_54_ram[160] = 0;
    exp_54_ram[161] = 1;
    exp_54_ram[162] = 0;
    exp_54_ram[163] = 0;
    exp_54_ram[164] = 252;
    exp_54_ram[165] = 252;
    exp_54_ram[166] = 43;
    exp_54_ram[167] = 0;
    exp_54_ram[168] = 0;
    exp_54_ram[169] = 222;
    exp_54_ram[170] = 236;
    exp_54_ram[171] = 2;
    exp_54_ram[172] = 128;
    exp_54_ram[173] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_230;
  assign exp_230 = exp_511;

  reg [3:0] exp_511_reg;
  always@(*) begin
    case (exp_363)
      0:exp_511_reg <= exp_498;
      1:exp_511_reg <= exp_503;
      2:exp_511_reg <= exp_504;
      3:exp_511_reg <= exp_505;
      4:exp_511_reg <= exp_506;
      5:exp_511_reg <= exp_507;
      6:exp_511_reg <= exp_508;
      7:exp_511_reg <= exp_509;
      default:exp_511_reg <= exp_510;
    endcase
  end
  assign exp_511 = exp_511_reg;
  assign exp_510 = 0;
  assign exp_498 = exp_494 << exp_497;
  assign exp_494 = 1;
  assign exp_497 = exp_496 + exp_495;
  assign exp_496 = 0;
  assign exp_495 = exp_431[1:0];
  assign exp_503 = exp_499 << exp_502;
  assign exp_499 = 3;
  assign exp_502 = exp_501 + exp_500;
  assign exp_501 = 0;
  assign exp_500 = exp_431[1:1];
  assign exp_504 = 15;
  assign exp_505 = 0;
  assign exp_506 = 0;
  assign exp_507 = 0;
  assign exp_508 = 0;
  assign exp_509 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_225;
  assign exp_225 = exp_493;

  reg [31:0] exp_493_reg;
  always@(*) begin
    case (exp_363)
      0:exp_493_reg <= exp_480;
      1:exp_493_reg <= exp_484;
      2:exp_493_reg <= exp_486;
      3:exp_493_reg <= exp_487;
      4:exp_493_reg <= exp_488;
      5:exp_493_reg <= exp_489;
      6:exp_493_reg <= exp_490;
      7:exp_493_reg <= exp_491;
      default:exp_493_reg <= exp_492;
    endcase
  end
  assign exp_493 = exp_493_reg;
  assign exp_492 = 0;

  reg [31:0] exp_480_reg;
  always@(*) begin
    case (exp_434)
      0:exp_480_reg <= exp_466;
      1:exp_480_reg <= exp_474;
      2:exp_480_reg <= exp_476;
      3:exp_480_reg <= exp_478;
      default:exp_480_reg <= exp_479;
    endcase
  end
  assign exp_480 = exp_480_reg;
  assign exp_479 = 0;
  assign exp_466 = exp_465;
  assign exp_465 = exp_464 + exp_463;
  assign exp_464 = 0;
  assign exp_463 = exp_353[7:0];

      reg [31:0] exp_353_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_353_reg <= exp_296;
        end
      end
      assign exp_353 = exp_353_reg;
      assign exp_474 = exp_466 << exp_473;
  assign exp_473 = 8;
  assign exp_476 = exp_466 << exp_475;
  assign exp_475 = 16;
  assign exp_478 = exp_466 << exp_477;
  assign exp_477 = 24;

  reg [31:0] exp_484_reg;
  always@(*) begin
    case (exp_437)
      0:exp_484_reg <= exp_470;
      1:exp_484_reg <= exp_482;
      default:exp_484_reg <= exp_483;
    endcase
  end
  assign exp_484 = exp_484_reg;
  assign exp_437 = exp_436 + exp_435;
  assign exp_436 = 0;
  assign exp_435 = exp_431[1:1];
  assign exp_483 = 0;
  assign exp_470 = exp_469;
  assign exp_469 = exp_468 + exp_467;
  assign exp_468 = 0;
  assign exp_467 = exp_353[15:0];
  assign exp_482 = exp_470 << exp_481;
  assign exp_481 = 16;
  assign exp_486 = exp_485 + exp_472;
  assign exp_485 = 0;
  assign exp_472 = exp_471 + exp_353;
  assign exp_471 = 0;
  assign exp_487 = 0;
  assign exp_488 = 0;
  assign exp_489 = 0;
  assign exp_490 = 0;
  assign exp_491 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 0;
    exp_47_ram[32] = 1;
    exp_47_ram[33] = 128;
    exp_47_ram[34] = 0;
    exp_47_ram[35] = 1;
    exp_47_ram[36] = 129;
    exp_47_ram[37] = 1;
    exp_47_ram[38] = 164;
    exp_47_ram[39] = 180;
    exp_47_ram[40] = 132;
    exp_47_ram[41] = 244;
    exp_47_ram[42] = 196;
    exp_47_ram[43] = 196;
    exp_47_ram[44] = 231;
    exp_47_ram[45] = 196;
    exp_47_ram[46] = 7;
    exp_47_ram[47] = 193;
    exp_47_ram[48] = 1;
    exp_47_ram[49] = 0;
    exp_47_ram[50] = 1;
    exp_47_ram[51] = 129;
    exp_47_ram[52] = 1;
    exp_47_ram[53] = 0;
    exp_47_ram[54] = 212;
    exp_47_ram[55] = 0;
    exp_47_ram[56] = 70;
    exp_47_ram[57] = 212;
    exp_47_ram[58] = 196;
    exp_47_ram[59] = 6;
    exp_47_ram[60] = 70;
    exp_47_ram[61] = 132;
    exp_47_ram[62] = 72;
    exp_47_ram[63] = 8;
    exp_47_ram[64] = 8;
    exp_47_ram[65] = 0;
    exp_47_ram[66] = 230;
    exp_47_ram[67] = 246;
    exp_47_ram[68] = 5;
    exp_47_ram[69] = 5;
    exp_47_ram[70] = 7;
    exp_47_ram[71] = 7;
    exp_47_ram[72] = 193;
    exp_47_ram[73] = 1;
    exp_47_ram[74] = 0;
    exp_47_ram[75] = 1;
    exp_47_ram[76] = 17;
    exp_47_ram[77] = 129;
    exp_47_ram[78] = 33;
    exp_47_ram[79] = 49;
    exp_47_ram[80] = 65;
    exp_47_ram[81] = 81;
    exp_47_ram[82] = 97;
    exp_47_ram[83] = 113;
    exp_47_ram[84] = 129;
    exp_47_ram[85] = 145;
    exp_47_ram[86] = 1;
    exp_47_ram[87] = 223;
    exp_47_ram[88] = 164;
    exp_47_ram[89] = 180;
    exp_47_ram[90] = 0;
    exp_47_ram[91] = 223;
    exp_47_ram[92] = 5;
    exp_47_ram[93] = 5;
    exp_47_ram[94] = 132;
    exp_47_ram[95] = 196;
    exp_47_ram[96] = 166;
    exp_47_ram[97] = 7;
    exp_47_ram[98] = 6;
    exp_47_ram[99] = 182;
    exp_47_ram[100] = 7;
    exp_47_ram[101] = 6;
    exp_47_ram[102] = 192;
    exp_47_ram[103] = 6;
    exp_47_ram[104] = 0;
    exp_47_ram[105] = 7;
    exp_47_ram[106] = 11;
    exp_47_ram[107] = 198;
    exp_47_ram[108] = 7;
    exp_47_ram[109] = 11;
    exp_47_ram[110] = 214;
    exp_47_ram[111] = 11;
    exp_47_ram[112] = 231;
    exp_47_ram[113] = 192;
    exp_47_ram[114] = 7;
    exp_47_ram[115] = 0;
    exp_47_ram[116] = 132;
    exp_47_ram[117] = 196;
    exp_47_ram[118] = 70;
    exp_47_ram[119] = 7;
    exp_47_ram[120] = 197;
    exp_47_ram[121] = 86;
    exp_47_ram[122] = 245;
    exp_47_ram[123] = 6;
    exp_47_ram[124] = 228;
    exp_47_ram[125] = 244;
    exp_47_ram[126] = 0;
    exp_47_ram[127] = 7;
    exp_47_ram[128] = 16;
    exp_47_ram[129] = 159;
    exp_47_ram[130] = 0;
    exp_47_ram[131] = 223;
    exp_47_ram[132] = 5;
    exp_47_ram[133] = 5;
    exp_47_ram[134] = 132;
    exp_47_ram[135] = 196;
    exp_47_ram[136] = 166;
    exp_47_ram[137] = 7;
    exp_47_ram[138] = 6;
    exp_47_ram[139] = 182;
    exp_47_ram[140] = 7;
    exp_47_ram[141] = 6;
    exp_47_ram[142] = 192;
    exp_47_ram[143] = 6;
    exp_47_ram[144] = 0;
    exp_47_ram[145] = 7;
    exp_47_ram[146] = 12;
    exp_47_ram[147] = 198;
    exp_47_ram[148] = 7;
    exp_47_ram[149] = 12;
    exp_47_ram[150] = 214;
    exp_47_ram[151] = 12;
    exp_47_ram[152] = 231;
    exp_47_ram[153] = 192;
    exp_47_ram[154] = 7;
    exp_47_ram[155] = 0;
    exp_47_ram[156] = 132;
    exp_47_ram[157] = 196;
    exp_47_ram[158] = 38;
    exp_47_ram[159] = 7;
    exp_47_ram[160] = 197;
    exp_47_ram[161] = 54;
    exp_47_ram[162] = 245;
    exp_47_ram[163] = 6;
    exp_47_ram[164] = 228;
    exp_47_ram[165] = 244;
    exp_47_ram[166] = 0;
    exp_47_ram[167] = 7;
    exp_47_ram[168] = 0;
    exp_47_ram[169] = 159;
    exp_47_ram[170] = 31;
    exp_47_ram[171] = 250;
    exp_47_ram[172] = 0;
    exp_47_ram[173] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 33;
    exp_40_ram[32] = 1;
    exp_40_ram[33] = 0;
    exp_40_ram[34] = 0;
    exp_40_ram[35] = 1;
    exp_40_ram[36] = 38;
    exp_40_ram[37] = 4;
    exp_40_ram[38] = 46;
    exp_40_ram[39] = 44;
    exp_40_ram[40] = 39;
    exp_40_ram[41] = 38;
    exp_40_ram[42] = 39;
    exp_40_ram[43] = 39;
    exp_40_ram[44] = 160;
    exp_40_ram[45] = 39;
    exp_40_ram[46] = 133;
    exp_40_ram[47] = 36;
    exp_40_ram[48] = 1;
    exp_40_ram[49] = 128;
    exp_40_ram[50] = 1;
    exp_40_ram[51] = 46;
    exp_40_ram[52] = 4;
    exp_40_ram[53] = 6;
    exp_40_ram[54] = 38;
    exp_40_ram[55] = 6;
    exp_40_ram[56] = 134;
    exp_40_ram[57] = 36;
    exp_40_ram[58] = 38;
    exp_40_ram[59] = 166;
    exp_40_ram[60] = 166;
    exp_40_ram[61] = 40;
    exp_40_ram[62] = 40;
    exp_40_ram[63] = 40;
    exp_40_ram[64] = 23;
    exp_40_ram[65] = 7;
    exp_40_ram[66] = 101;
    exp_40_ram[67] = 229;
    exp_40_ram[68] = 7;
    exp_40_ram[69] = 135;
    exp_40_ram[70] = 5;
    exp_40_ram[71] = 133;
    exp_40_ram[72] = 36;
    exp_40_ram[73] = 1;
    exp_40_ram[74] = 128;
    exp_40_ram[75] = 1;
    exp_40_ram[76] = 46;
    exp_40_ram[77] = 44;
    exp_40_ram[78] = 42;
    exp_40_ram[79] = 40;
    exp_40_ram[80] = 38;
    exp_40_ram[81] = 36;
    exp_40_ram[82] = 34;
    exp_40_ram[83] = 32;
    exp_40_ram[84] = 46;
    exp_40_ram[85] = 44;
    exp_40_ram[86] = 4;
    exp_40_ram[87] = 240;
    exp_40_ram[88] = 36;
    exp_40_ram[89] = 38;
    exp_40_ram[90] = 0;
    exp_40_ram[91] = 240;
    exp_40_ram[92] = 6;
    exp_40_ram[93] = 134;
    exp_40_ram[94] = 37;
    exp_40_ram[95] = 37;
    exp_40_ram[96] = 7;
    exp_40_ram[97] = 8;
    exp_40_ram[98] = 56;
    exp_40_ram[99] = 135;
    exp_40_ram[100] = 134;
    exp_40_ram[101] = 135;
    exp_40_ram[102] = 38;
    exp_40_ram[103] = 139;
    exp_40_ram[104] = 11;
    exp_40_ram[105] = 134;
    exp_40_ram[106] = 134;
    exp_40_ram[107] = 224;
    exp_40_ram[108] = 134;
    exp_40_ram[109] = 134;
    exp_40_ram[110] = 22;
    exp_40_ram[111] = 7;
    exp_40_ram[112] = 230;
    exp_40_ram[113] = 39;
    exp_40_ram[114] = 138;
    exp_40_ram[115] = 10;
    exp_40_ram[116] = 38;
    exp_40_ram[117] = 38;
    exp_40_ram[118] = 7;
    exp_40_ram[119] = 5;
    exp_40_ram[120] = 181;
    exp_40_ram[121] = 135;
    exp_40_ram[122] = 134;
    exp_40_ram[123] = 135;
    exp_40_ram[124] = 36;
    exp_40_ram[125] = 38;
    exp_40_ram[126] = 39;
    exp_40_ram[127] = 133;
    exp_40_ram[128] = 5;
    exp_40_ram[129] = 240;
    exp_40_ram[130] = 0;
    exp_40_ram[131] = 240;
    exp_40_ram[132] = 6;
    exp_40_ram[133] = 134;
    exp_40_ram[134] = 37;
    exp_40_ram[135] = 37;
    exp_40_ram[136] = 7;
    exp_40_ram[137] = 8;
    exp_40_ram[138] = 56;
    exp_40_ram[139] = 135;
    exp_40_ram[140] = 134;
    exp_40_ram[141] = 135;
    exp_40_ram[142] = 38;
    exp_40_ram[143] = 140;
    exp_40_ram[144] = 12;
    exp_40_ram[145] = 134;
    exp_40_ram[146] = 134;
    exp_40_ram[147] = 224;
    exp_40_ram[148] = 134;
    exp_40_ram[149] = 134;
    exp_40_ram[150] = 22;
    exp_40_ram[151] = 7;
    exp_40_ram[152] = 230;
    exp_40_ram[153] = 39;
    exp_40_ram[154] = 137;
    exp_40_ram[155] = 9;
    exp_40_ram[156] = 38;
    exp_40_ram[157] = 38;
    exp_40_ram[158] = 7;
    exp_40_ram[159] = 5;
    exp_40_ram[160] = 181;
    exp_40_ram[161] = 135;
    exp_40_ram[162] = 134;
    exp_40_ram[163] = 135;
    exp_40_ram[164] = 36;
    exp_40_ram[165] = 38;
    exp_40_ram[166] = 39;
    exp_40_ram[167] = 133;
    exp_40_ram[168] = 5;
    exp_40_ram[169] = 240;
    exp_40_ram[170] = 240;
    exp_40_ram[171] = 240;
    exp_40_ram[172] = 0;
    exp_40_ram[173] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 55;
    exp_33_ram[32] = 19;
    exp_33_ram[33] = 239;
    exp_33_ram[34] = 111;
    exp_33_ram[35] = 19;
    exp_33_ram[36] = 35;
    exp_33_ram[37] = 19;
    exp_33_ram[38] = 35;
    exp_33_ram[39] = 35;
    exp_33_ram[40] = 131;
    exp_33_ram[41] = 35;
    exp_33_ram[42] = 3;
    exp_33_ram[43] = 131;
    exp_33_ram[44] = 35;
    exp_33_ram[45] = 131;
    exp_33_ram[46] = 19;
    exp_33_ram[47] = 3;
    exp_33_ram[48] = 19;
    exp_33_ram[49] = 103;
    exp_33_ram[50] = 19;
    exp_33_ram[51] = 35;
    exp_33_ram[52] = 19;
    exp_33_ram[53] = 183;
    exp_33_ram[54] = 35;
    exp_33_ram[55] = 183;
    exp_33_ram[56] = 147;
    exp_33_ram[57] = 35;
    exp_33_ram[58] = 131;
    exp_33_ram[59] = 3;
    exp_33_ram[60] = 131;
    exp_33_ram[61] = 3;
    exp_33_ram[62] = 131;
    exp_33_ram[63] = 3;
    exp_33_ram[64] = 147;
    exp_33_ram[65] = 19;
    exp_33_ram[66] = 51;
    exp_33_ram[67] = 179;
    exp_33_ram[68] = 19;
    exp_33_ram[69] = 147;
    exp_33_ram[70] = 19;
    exp_33_ram[71] = 147;
    exp_33_ram[72] = 3;
    exp_33_ram[73] = 19;
    exp_33_ram[74] = 103;
    exp_33_ram[75] = 19;
    exp_33_ram[76] = 35;
    exp_33_ram[77] = 35;
    exp_33_ram[78] = 35;
    exp_33_ram[79] = 35;
    exp_33_ram[80] = 35;
    exp_33_ram[81] = 35;
    exp_33_ram[82] = 35;
    exp_33_ram[83] = 35;
    exp_33_ram[84] = 35;
    exp_33_ram[85] = 35;
    exp_33_ram[86] = 19;
    exp_33_ram[87] = 239;
    exp_33_ram[88] = 35;
    exp_33_ram[89] = 35;
    exp_33_ram[90] = 19;
    exp_33_ram[91] = 239;
    exp_33_ram[92] = 19;
    exp_33_ram[93] = 147;
    exp_33_ram[94] = 3;
    exp_33_ram[95] = 131;
    exp_33_ram[96] = 51;
    exp_33_ram[97] = 19;
    exp_33_ram[98] = 51;
    exp_33_ram[99] = 179;
    exp_33_ram[100] = 179;
    exp_33_ram[101] = 147;
    exp_33_ram[102] = 131;
    exp_33_ram[103] = 19;
    exp_33_ram[104] = 147;
    exp_33_ram[105] = 19;
    exp_33_ram[106] = 147;
    exp_33_ram[107] = 227;
    exp_33_ram[108] = 19;
    exp_33_ram[109] = 147;
    exp_33_ram[110] = 99;
    exp_33_ram[111] = 147;
    exp_33_ram[112] = 227;
    exp_33_ram[113] = 131;
    exp_33_ram[114] = 19;
    exp_33_ram[115] = 147;
    exp_33_ram[116] = 3;
    exp_33_ram[117] = 131;
    exp_33_ram[118] = 51;
    exp_33_ram[119] = 147;
    exp_33_ram[120] = 179;
    exp_33_ram[121] = 179;
    exp_33_ram[122] = 179;
    exp_33_ram[123] = 147;
    exp_33_ram[124] = 35;
    exp_33_ram[125] = 35;
    exp_33_ram[126] = 131;
    exp_33_ram[127] = 147;
    exp_33_ram[128] = 19;
    exp_33_ram[129] = 239;
    exp_33_ram[130] = 19;
    exp_33_ram[131] = 239;
    exp_33_ram[132] = 19;
    exp_33_ram[133] = 147;
    exp_33_ram[134] = 3;
    exp_33_ram[135] = 131;
    exp_33_ram[136] = 51;
    exp_33_ram[137] = 19;
    exp_33_ram[138] = 51;
    exp_33_ram[139] = 179;
    exp_33_ram[140] = 179;
    exp_33_ram[141] = 147;
    exp_33_ram[142] = 131;
    exp_33_ram[143] = 19;
    exp_33_ram[144] = 147;
    exp_33_ram[145] = 19;
    exp_33_ram[146] = 147;
    exp_33_ram[147] = 227;
    exp_33_ram[148] = 19;
    exp_33_ram[149] = 147;
    exp_33_ram[150] = 99;
    exp_33_ram[151] = 147;
    exp_33_ram[152] = 227;
    exp_33_ram[153] = 131;
    exp_33_ram[154] = 19;
    exp_33_ram[155] = 147;
    exp_33_ram[156] = 3;
    exp_33_ram[157] = 131;
    exp_33_ram[158] = 51;
    exp_33_ram[159] = 147;
    exp_33_ram[160] = 179;
    exp_33_ram[161] = 179;
    exp_33_ram[162] = 179;
    exp_33_ram[163] = 147;
    exp_33_ram[164] = 35;
    exp_33_ram[165] = 35;
    exp_33_ram[166] = 131;
    exp_33_ram[167] = 147;
    exp_33_ram[168] = 19;
    exp_33_ram[169] = 239;
    exp_33_ram[170] = 111;
    exp_33_ram[171] = 128;
    exp_33_ram[172] = 12;
    exp_33_ram[173] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_179;

  reg [31:0] exp_179_reg;
  always@(*) begin
    case (exp_177)
      0:exp_179_reg <= exp_157;
      1:exp_179_reg <= exp_167;
      default:exp_179_reg <= exp_178;
    endcase
  end
  assign exp_179 = exp_179_reg;
  assign exp_177 = exp_139[2:2];
  assign exp_139 = exp_1;
  assign exp_178 = 0;

      reg [31:0] exp_157_reg = 0;
      always@(posedge clk) begin
        if (exp_156) begin
          exp_157_reg <= exp_164;
        end
      end
      assign exp_157 = exp_157_reg;
    
  reg [31:0] exp_164_reg;
  always@(*) begin
    case (exp_159)
      0:exp_164_reg <= exp_161;
      1:exp_164_reg <= exp_162;
      default:exp_164_reg <= exp_163;
    endcase
  end
  assign exp_164 = exp_164_reg;
  assign exp_159 = exp_157 == exp_158;
  assign exp_158 = 4294967295;
  assign exp_163 = 0;
  assign exp_161 = exp_157 + exp_160;
  assign exp_160 = 1;
  assign exp_162 = 0;
  assign exp_156 = 1;

      reg [31:0] exp_167_reg = 0;
      always@(posedge clk) begin
        if (exp_166) begin
          exp_167_reg <= exp_174;
        end
      end
      assign exp_167 = exp_167_reg;
    
  reg [31:0] exp_174_reg;
  always@(*) begin
    case (exp_169)
      0:exp_174_reg <= exp_171;
      1:exp_174_reg <= exp_172;
      default:exp_174_reg <= exp_173;
    endcase
  end
  assign exp_174 = exp_174_reg;
  assign exp_169 = exp_167 == exp_168;
  assign exp_168 = 4294967295;
  assign exp_173 = 0;
  assign exp_171 = exp_167 + exp_170;
  assign exp_170 = 1;
  assign exp_172 = 0;
  assign exp_166 = exp_159 & exp_165;
  assign exp_165 = 1;
  assign exp_182 = exp_201;
  assign exp_201 = 0;
  assign exp_204 = exp_219;
  assign exp_219 = stdin_in;
  assign exp_439 = exp_226[15:8];
  assign exp_440 = exp_226[23:16];
  assign exp_441 = exp_226[31:24];
  assign exp_453 = $signed(exp_452);
  assign exp_452 = exp_451 + exp_447;
  assign exp_451 = 0;

  reg [15:0] exp_447_reg;
  always@(*) begin
    case (exp_437)
      0:exp_447_reg <= exp_444;
      1:exp_447_reg <= exp_445;
      default:exp_447_reg <= exp_446;
    endcase
  end
  assign exp_447 = exp_447_reg;
  assign exp_446 = 0;
  assign exp_444 = exp_226[15:0];
  assign exp_445 = exp_226[31:16];
  assign exp_454 = 0;
  assign exp_455 = exp_443;
  assign exp_456 = exp_447;
  assign exp_457 = 0;
  assign exp_458 = 0;

  reg [31:0] exp_817_reg;
  always@(*) begin
    case (exp_607)
      0:exp_817_reg <= exp_813;
      1:exp_817_reg <= exp_815;
      default:exp_817_reg <= exp_816;
    endcase
  end
  assign exp_817 = exp_817_reg;
  assign exp_816 = 0;

  reg [31:0] exp_813_reg;
  always@(*) begin
    case (exp_584)
      0:exp_813_reg <= exp_808;
      1:exp_813_reg <= exp_809;
      default:exp_813_reg <= exp_812;
    endcase
  end
  assign exp_813 = exp_813_reg;
  assign exp_584 = exp_583 & exp_581;
  assign exp_583 = exp_576 == exp_582;
  assign exp_582 = 0;
  assign exp_812 = 0;
  assign exp_808 = exp_807[63:32];

  reg [63:0] exp_807_reg;
  always@(*) begin
    case (exp_804)
      0:exp_807_reg <= exp_803;
      1:exp_807_reg <= exp_805;
      default:exp_807_reg <= exp_806;
    endcase
  end
  assign exp_807 = exp_807_reg;

      reg [0:0] exp_804_reg = 0;
      always@(posedge clk) begin
        if (exp_789) begin
          exp_804_reg <= exp_787;
        end
      end
      assign exp_804 = exp_804_reg;
    
      reg [0:0] exp_787_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_787_reg <= exp_764;
        end
      end
      assign exp_787 = exp_787_reg;
    
      reg [0:0] exp_764_reg = 0;
      always@(posedge clk) begin
        if (exp_746) begin
          exp_764_reg <= exp_761;
        end
      end
      assign exp_764 = exp_764_reg;
      assign exp_761 = exp_759 ^ exp_760;
  assign exp_759 = exp_741 & exp_724;
  assign exp_741 = exp_740 + exp_739;
  assign exp_740 = 0;
  assign exp_739 = exp_737[31:31];

      reg [31:0] exp_737_reg = 0;
      always@(posedge clk) begin
        if (exp_736) begin
          exp_737_reg <= exp_354;
        end
      end
      assign exp_737 = exp_737_reg;
      assign exp_736 = exp_726 == exp_735;
  assign exp_735 = 0;
  assign exp_724 = exp_723 | exp_590;
  assign exp_723 = exp_584 | exp_587;
  assign exp_587 = exp_586 & exp_581;
  assign exp_586 = exp_576 == exp_585;
  assign exp_585 = 1;
  assign exp_590 = exp_589 & exp_581;
  assign exp_589 = exp_576 == exp_588;
  assign exp_588 = 2;
  assign exp_760 = exp_744 & exp_725;
  assign exp_744 = exp_743 + exp_742;
  assign exp_743 = 0;
  assign exp_742 = exp_738[31:31];

      reg [31:0] exp_738_reg = 0;
      always@(posedge clk) begin
        if (exp_736) begin
          exp_738_reg <= exp_355;
        end
      end
      assign exp_738 = exp_738_reg;
      assign exp_725 = exp_584 | exp_587;
  assign exp_746 = exp_726 == exp_745;
  assign exp_745 = 1;
  assign exp_766 = exp_726 == exp_765;
  assign exp_765 = 2;
  assign exp_789 = exp_726 == exp_788;
  assign exp_788 = 3;
  assign exp_806 = 0;

      reg [63:0] exp_803_reg = 0;
      always@(posedge clk) begin
        if (exp_789) begin
          exp_803_reg <= exp_802;
        end
      end
      assign exp_803 = exp_803_reg;
      assign exp_802 = exp_798 + exp_801;
  assign exp_798 = exp_794 + exp_797;
  assign exp_794 = exp_790 + exp_793;
  assign exp_790 = exp_783;

      reg [31:0] exp_783_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_783_reg <= exp_770;
        end
      end
      assign exp_783 = exp_783_reg;
      assign exp_770 = exp_768 * exp_769;
  assign exp_768 = exp_767;
  assign exp_767 = exp_762[15:0];

      reg [31:0] exp_762_reg = 0;
      always@(posedge clk) begin
        if (exp_746) begin
          exp_762_reg <= exp_752;
        end
      end
      assign exp_762 = exp_762_reg;
      assign exp_752 = exp_751 + exp_750;
  assign exp_751 = 0;

  reg [31:0] exp_750_reg;
  always@(*) begin
    case (exp_747)
      0:exp_750_reg <= exp_737;
      1:exp_750_reg <= exp_748;
      default:exp_750_reg <= exp_749;
    endcase
  end
  assign exp_750 = exp_750_reg;
  assign exp_747 = exp_741 & exp_724;
  assign exp_749 = 0;
  assign exp_748 = -exp_737;
  assign exp_769 = exp_763[15:0];

      reg [31:0] exp_763_reg = 0;
      always@(posedge clk) begin
        if (exp_746) begin
          exp_763_reg <= exp_758;
        end
      end
      assign exp_763 = exp_763_reg;
      assign exp_758 = exp_757 + exp_756;
  assign exp_757 = 0;

  reg [31:0] exp_756_reg;
  always@(*) begin
    case (exp_753)
      0:exp_756_reg <= exp_738;
      1:exp_756_reg <= exp_754;
      default:exp_756_reg <= exp_755;
    endcase
  end
  assign exp_756 = exp_756_reg;
  assign exp_753 = exp_744 & exp_725;
  assign exp_755 = 0;
  assign exp_754 = -exp_738;
  assign exp_793 = exp_791 << exp_792;
  assign exp_791 = exp_784;

      reg [31:0] exp_784_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_784_reg <= exp_774;
        end
      end
      assign exp_784 = exp_784_reg;
      assign exp_774 = exp_772 * exp_773;
  assign exp_772 = exp_771;
  assign exp_771 = exp_762[15:0];
  assign exp_773 = exp_763[31:16];
  assign exp_792 = 16;
  assign exp_797 = exp_795 << exp_796;
  assign exp_795 = exp_785;

      reg [31:0] exp_785_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_785_reg <= exp_778;
        end
      end
      assign exp_785 = exp_785_reg;
      assign exp_778 = exp_776 * exp_777;
  assign exp_776 = exp_775;
  assign exp_775 = exp_762[31:16];
  assign exp_777 = exp_763[15:0];
  assign exp_796 = 16;
  assign exp_801 = exp_799 << exp_800;
  assign exp_799 = exp_786;

      reg [31:0] exp_786_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_786_reg <= exp_782;
        end
      end
      assign exp_786 = exp_786_reg;
      assign exp_782 = exp_780 * exp_781;
  assign exp_780 = exp_779;
  assign exp_779 = exp_762[31:16];
  assign exp_781 = exp_763[31:16];
  assign exp_800 = 32;
  assign exp_805 = -exp_803;
  assign exp_809 = exp_807[31:0];

  reg [31:0] exp_815_reg;
  always@(*) begin
    case (exp_608)
      0:exp_815_reg <= exp_718;
      1:exp_815_reg <= exp_719;
      default:exp_815_reg <= exp_814;
    endcase
  end
  assign exp_815 = exp_815_reg;
  assign exp_608 = exp_576[1:1];
  assign exp_814 = 0;

      reg [31:0] exp_718_reg = 0;
      always@(posedge clk) begin
        if (exp_627) begin
          exp_718_reg <= exp_712;
        end
      end
      assign exp_718 = exp_718_reg;
    
  reg [31:0] exp_712_reg;
  always@(*) begin
    case (exp_708)
      0:exp_712_reg <= exp_699;
      1:exp_712_reg <= exp_710;
      default:exp_712_reg <= exp_711;
    endcase
  end
  assign exp_712 = exp_712_reg;
  assign exp_708 = exp_707 & exp_610;
  assign exp_707 = exp_656 == exp_706;

      reg [31:0] exp_656_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_656_reg <= exp_653;
        end
      end
      assign exp_656 = exp_656_reg;
      assign exp_653 = exp_652 + exp_651;
  assign exp_652 = 0;

  reg [31:0] exp_651_reg;
  always@(*) begin
    case (exp_648)
      0:exp_651_reg <= exp_633;
      1:exp_651_reg <= exp_649;
      default:exp_651_reg <= exp_650;
    endcase
  end
  assign exp_651 = exp_651_reg;
  assign exp_648 = exp_639 & exp_610;
  assign exp_639 = exp_638 + exp_637;
  assign exp_638 = 0;
  assign exp_637 = exp_633[31:31];

      reg [31:0] exp_633_reg = 0;
      always@(posedge clk) begin
        if (exp_631) begin
          exp_633_reg <= exp_355;
        end
      end
      assign exp_633 = exp_633_reg;
      assign exp_631 = exp_613 == exp_630;
  assign exp_630 = 0;
  assign exp_610 = ~exp_609;
  assign exp_609 = exp_576[0:0];
  assign exp_650 = 0;
  assign exp_649 = -exp_633;
  assign exp_641 = exp_613 == exp_640;
  assign exp_640 = 1;
  assign exp_706 = 0;
  assign exp_711 = 0;
  assign exp_699 = exp_698 + exp_697;
  assign exp_698 = 0;

  reg [31:0] exp_697_reg;
  always@(*) begin
    case (exp_694)
      0:exp_697_reg <= exp_692;
      1:exp_697_reg <= exp_695;
      default:exp_697_reg <= exp_696;
    endcase
  end
  assign exp_697 = exp_697_reg;
  assign exp_694 = exp_658 & exp_610;

      reg [0:0] exp_658_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_658_reg <= exp_654;
        end
      end
      assign exp_658 = exp_658_reg;
      assign exp_654 = exp_636 ^ exp_639;
  assign exp_636 = exp_635 + exp_634;
  assign exp_635 = 0;
  assign exp_634 = exp_632[31:31];

      reg [31:0] exp_632_reg = 0;
      always@(posedge clk) begin
        if (exp_631) begin
          exp_632_reg <= exp_354;
        end
      end
      assign exp_632 = exp_632_reg;
      assign exp_696 = 0;

      reg [31:0] exp_692_reg = 0;
      always@(posedge clk) begin
        if (exp_625) begin
          exp_692_reg <= exp_662;
        end
      end
      assign exp_692 = exp_692_reg;
    
      reg [31:0] exp_662_reg = 0;
      always@(posedge clk) begin
        if (exp_661) begin
          exp_662_reg <= exp_689;
        end
      end
      assign exp_662 = exp_662_reg;
    
  reg [31:0] exp_689_reg;
  always@(*) begin
    case (exp_623)
      0:exp_689_reg <= exp_681;
      1:exp_689_reg <= exp_687;
      default:exp_689_reg <= exp_688;
    endcase
  end
  assign exp_689 = exp_689_reg;
  assign exp_623 = exp_613 == exp_622;
  assign exp_622 = 2;
  assign exp_688 = 0;

  reg [31:0] exp_681_reg;
  always@(*) begin
    case (exp_671)
      0:exp_681_reg <= exp_675;
      1:exp_681_reg <= exp_679;
      default:exp_681_reg <= exp_680;
    endcase
  end
  assign exp_681 = exp_681_reg;
  assign exp_671 = ~exp_670;
  assign exp_670 = exp_669[32:32];
  assign exp_669 = exp_668 - exp_656;
  assign exp_668 = exp_667;
  assign exp_667 = {exp_665, exp_666};  assign exp_665 = exp_660[31:0];

      reg [31:0] exp_660_reg = 0;
      always@(posedge clk) begin
        if (exp_659) begin
          exp_660_reg <= exp_686;
        end
      end
      assign exp_660 = exp_660_reg;
    
  reg [32:0] exp_686_reg;
  always@(*) begin
    case (exp_623)
      0:exp_686_reg <= exp_673;
      1:exp_686_reg <= exp_684;
      default:exp_686_reg <= exp_685;
    endcase
  end
  assign exp_686 = exp_686_reg;
  assign exp_685 = 0;

  reg [32:0] exp_673_reg;
  always@(*) begin
    case (exp_671)
      0:exp_673_reg <= exp_667;
      1:exp_673_reg <= exp_669;
      default:exp_673_reg <= exp_672;
    endcase
  end
  assign exp_673 = exp_673_reg;
  assign exp_672 = 0;
  assign exp_684 = 0;
  assign exp_659 = 1;
  assign exp_666 = exp_664[31:31];

      reg [31:0] exp_664_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_664_reg <= exp_691;
        end
      end
      assign exp_664 = exp_664_reg;
    
  reg [31:0] exp_691_reg;
  always@(*) begin
    case (exp_623)
      0:exp_691_reg <= exp_683;
      1:exp_691_reg <= exp_655;
      default:exp_691_reg <= exp_690;
    endcase
  end
  assign exp_691 = exp_691_reg;
  assign exp_690 = 0;
  assign exp_683 = exp_664 << exp_682;
  assign exp_682 = 1;

      reg [31:0] exp_655_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_655_reg <= exp_647;
        end
      end
      assign exp_655 = exp_655_reg;
      assign exp_647 = exp_646 + exp_645;
  assign exp_646 = 0;

  reg [31:0] exp_645_reg;
  always@(*) begin
    case (exp_642)
      0:exp_645_reg <= exp_632;
      1:exp_645_reg <= exp_643;
      default:exp_645_reg <= exp_644;
    endcase
  end
  assign exp_645 = exp_645_reg;
  assign exp_642 = exp_636 & exp_610;
  assign exp_644 = 0;
  assign exp_643 = -exp_632;
  assign exp_663 = 1;
  assign exp_680 = 0;
  assign exp_675 = exp_662 << exp_674;
  assign exp_674 = 1;
  assign exp_679 = exp_677 | exp_678;
  assign exp_677 = exp_662 << exp_676;
  assign exp_676 = 1;
  assign exp_678 = 1;
  assign exp_687 = 0;
  assign exp_661 = 1;
  assign exp_625 = exp_613 == exp_624;
  assign exp_624 = 35;
  assign exp_695 = -exp_692;
  assign exp_710 = $signed(exp_709);
  assign exp_709 = -1;
  assign exp_627 = exp_613 == exp_626;
  assign exp_626 = 36;

      reg [31:0] exp_719_reg = 0;
      always@(posedge clk) begin
        if (exp_627) begin
          exp_719_reg <= exp_717;
        end
      end
      assign exp_719 = exp_719_reg;
    
  reg [31:0] exp_717_reg;
  always@(*) begin
    case (exp_715)
      0:exp_717_reg <= exp_705;
      1:exp_717_reg <= exp_632;
      default:exp_717_reg <= exp_716;
    endcase
  end
  assign exp_717 = exp_717_reg;
  assign exp_715 = exp_714 & exp_610;
  assign exp_714 = exp_656 == exp_713;
  assign exp_713 = 0;
  assign exp_716 = 0;
  assign exp_705 = exp_704 + exp_703;
  assign exp_704 = 0;

  reg [31:0] exp_703_reg;
  always@(*) begin
    case (exp_700)
      0:exp_703_reg <= exp_693;
      1:exp_703_reg <= exp_701;
      default:exp_703_reg <= exp_702;
    endcase
  end
  assign exp_703 = exp_703_reg;
  assign exp_700 = exp_657 & exp_610;

      reg [0:0] exp_657_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_657_reg <= exp_636;
        end
      end
      assign exp_657 = exp_657_reg;
      assign exp_702 = 0;

      reg [31:0] exp_693_reg = 0;
      always@(posedge clk) begin
        if (exp_625) begin
          exp_693_reg <= exp_660;
        end
      end
      assign exp_693 = exp_693_reg;
      assign exp_701 = -exp_693;
  assign exp_288 = $signed(exp_287);
  assign exp_287 = 0;
  assign exp_517 = exp_352 != exp_353;
  assign exp_530 = 0;
  assign exp_531 = 0;
  assign exp_518 = $signed(exp_352) < $signed(exp_353);
  assign exp_519 = $signed(exp_352) >= $signed(exp_353);
  assign exp_524 = exp_521 < exp_523;
  assign exp_521 = exp_520 + exp_352;
  assign exp_520 = 0;
  assign exp_523 = exp_522 + exp_353;
  assign exp_522 = 0;
  assign exp_529 = exp_526 >= exp_528;
  assign exp_526 = exp_525 + exp_352;
  assign exp_525 = 0;
  assign exp_528 = exp_527 + exp_353;
  assign exp_527 = 0;
  assign exp_844 = 0;
  assign exp_843 = exp_242 + exp_842;
  assign exp_842 = 4;

  reg [32:0] exp_574_reg;
  always@(*) begin
    case (exp_375)
      0:exp_574_reg <= exp_564;
      1:exp_574_reg <= exp_572;
      default:exp_574_reg <= exp_573;
    endcase
  end
  assign exp_574 = exp_574_reg;
  assign exp_573 = 0;
  assign exp_564 = exp_563 + exp_361;

  reg [31:0] exp_563_reg;
  always@(*) begin
    case (exp_373)
      0:exp_563_reg <= exp_549;
      1:exp_563_reg <= exp_561;
      default:exp_563_reg <= exp_562;
    endcase
  end
  assign exp_563 = exp_563_reg;
  assign exp_562 = 0;
  assign exp_549 = $signed(exp_548);
  assign exp_548 = exp_547 + exp_546;
  assign exp_547 = 0;
  assign exp_546 = {exp_545, exp_542};  assign exp_545 = {exp_544, exp_541};  assign exp_544 = {exp_543, exp_540};  assign exp_543 = {exp_538, exp_539};  assign exp_538 = exp_360[31:31];
  assign exp_539 = exp_360[7:7];
  assign exp_540 = exp_360[30:25];
  assign exp_541 = exp_360[11:8];
  assign exp_542 = 0;
  assign exp_561 = $signed(exp_560);
  assign exp_560 = exp_559 + exp_558;
  assign exp_559 = 0;
  assign exp_558 = {exp_557, exp_554};  assign exp_557 = {exp_556, exp_553};  assign exp_556 = {exp_555, exp_552};  assign exp_555 = {exp_550, exp_551};  assign exp_550 = exp_360[31:31];
  assign exp_551 = exp_360[19:12];
  assign exp_552 = exp_360[20:20];
  assign exp_553 = exp_360[30:21];
  assign exp_554 = 0;

      reg [31:0] exp_361_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_361_reg <= exp_244;
        end
      end
      assign exp_361 = exp_361_reg;
      assign exp_572 = exp_571 & exp_570;
  assign exp_571 = $signed(exp_569);
  assign exp_569 = exp_352 + exp_568;
  assign exp_568 = $signed(exp_567);
  assign exp_567 = exp_566 + exp_565;
  assign exp_566 = 0;
  assign exp_565 = exp_360[31:20];
  assign exp_570 = 4294967294;
  assign exp_241 = exp_234 & exp_232;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_243;
  assign exp_376 = 3;
  assign exp_222 = ~exp_207;
  assign exp_207 = exp_6;
  assign exp_200 = exp_184 & exp_185;
  assign exp_184 = exp_192;
  assign exp_192 = exp_5 & exp_191;
  assign exp_185 = exp_6;
  assign exp_181 = exp_2;
  assign stdin_ready_out = exp_223;
  assign stdout_valid_out = exp_200;
  assign stdout_out = exp_181;

endmodule