
module soc(clk, stdin_rx, stdout_tx, leds_out);
  input [0:0] stdin_rx;
  input [0:0] clk;
  output [0:0] stdout_tx;
  output [31:0] leds_out;
  wire [0:0] exp_280;
  wire [0:0] exp_277;
  wire [0:0] exp_201;
  wire [0:0] exp_204;
  wire [0:0] exp_199;
  wire [0:0] exp_262;
  wire [0:0] exp_247;
  wire [0:0] exp_261;
  wire [0:0] exp_258;
  wire [0:0] exp_257;
  wire [0:0] exp_221;
  wire [0:0] exp_245;
  wire [0:0] exp_241;
  wire [0:0] exp_206;
  wire [0:0] exp_219;
  wire [0:0] exp_216;
  wire [0:0] exp_198;
  wire [0:0] exp_184;
  wire [0:0] exp_192;
  wire [0:0] exp_5;
  wire [0:0] exp_396;
  wire [0:0] exp_743;
  wire [0:0] exp_680;
  wire [0:0] exp_545;
  wire [6:0] exp_530;
  wire [31:0] exp_528;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [12:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_410;
  wire [32:0] exp_1013;
  wire [0:0] exp_1009;
  wire [0:0] exp_705;
  wire [0:0] exp_683;
  wire [0:0] exp_541;
  wire [6:0] exp_540;
  wire [0:0] exp_543;
  wire [6:0] exp_542;
  wire [0:0] exp_704;
  wire [0:0] exp_549;
  wire [6:0] exp_548;
  wire [0:0] exp_703;
  wire [0:0] exp_702;
  wire [0:0] exp_701;
  wire [2:0] exp_531;
  wire [0:0] exp_700;
  wire [0:0] exp_684;
  wire [31:0] exp_520;
  wire [31:0] exp_458;
  wire [0:0] exp_454;
  wire [4:0] exp_434;
  wire [0:0] exp_453;
  wire [0:0] exp_457;
  wire [31:0] exp_450;
  wire [0:0] exp_431;
  wire [0:0] exp_1004;
  wire [0:0] exp_1003;
  wire [0:0] exp_1002;
  wire [0:0] exp_1001;
  wire [4:0] exp_413;
  wire [4:0] exp_996;
  wire [0:0] exp_995;
  wire [0:0] exp_587;
  wire [0:0] exp_586;
  wire [0:0] exp_585;
  wire [0:0] exp_584;
  wire [0:0] exp_583;
  wire [0:0] exp_582;
  wire [0:0] exp_533;
  wire [4:0] exp_532;
  wire [0:0] exp_535;
  wire [5:0] exp_534;
  wire [0:0] exp_537;
  wire [5:0] exp_536;
  wire [0:0] exp_539;
  wire [4:0] exp_538;
  wire [0:0] exp_990;
  wire [0:0] exp_989;
  wire [0:0] exp_775;
  wire [0:0] exp_749;
  wire [0:0] exp_747;
  wire [6:0] exp_745;
  wire [5:0] exp_746;
  wire [0:0] exp_748;
  wire [0:0] exp_774;
  wire [2:0] exp_744;
  wire [0:0] exp_988;
  wire [0:0] exp_986;
  wire [0:0] exp_979;
  wire [2:0] exp_894;
  wire [2:0] exp_901;
  wire [0:0] exp_896;
  wire [2:0] exp_895;
  wire [0:0] exp_900;
  wire [2:0] exp_898;
  wire [0:0] exp_897;
  wire [0:0] exp_899;
  wire [0:0] exp_890;
  wire [0:0] exp_889;
  wire [0:0] exp_888;
  wire [2:0] exp_978;
  wire [0:0] exp_987;
  wire [0:0] exp_797;
  wire [5:0] exp_781;
  wire [5:0] exp_788;
  wire [0:0] exp_783;
  wire [5:0] exp_782;
  wire [0:0] exp_787;
  wire [5:0] exp_785;
  wire [0:0] exp_784;
  wire [0:0] exp_786;
  wire [5:0] exp_796;
  wire [0:0] exp_408;
  wire [0:0] exp_407;
  wire [0:0] exp_405;
  wire [0:0] exp_404;
  wire [0:0] exp_402;
  wire [0:0] exp_403;
  wire [0:0] exp_401;
  wire [0:0] exp_1014;
  wire [0:0] exp_400;
  wire [0:0] exp_399;
  wire [0:0] exp_1018;
  wire [0:0] exp_1017;
  wire [0:0] exp_1016;
  wire [0:0] exp_1015;
  wire [0:0] exp_395;
  wire [0:0] exp_321;
  wire [0:0] exp_316;
  wire [0:0] exp_313;
  wire [31:0] exp_1;
  wire [31:0] exp_392;
  wire [31:0] exp_599;
  wire [31:0] exp_598;
  wire [31:0] exp_597;
  wire [31:0] exp_596;
  wire [11:0] exp_595;
  wire [11:0] exp_594;
  wire [11:0] exp_593;
  wire [0:0] exp_547;
  wire [5:0] exp_546;
  wire [0:0] exp_592;
  wire [11:0] exp_588;
  wire [11:0] exp_591;
  wire [6:0] exp_589;
  wire [4:0] exp_590;
  wire [31:0] exp_312;
  wire [0:0] exp_315;
  wire [31:0] exp_314;
  wire [0:0] exp_320;
  wire [0:0] exp_298;
  wire [0:0] exp_293;
  wire [0:0] exp_290;
  wire [31:0] exp_289;
  wire [0:0] exp_292;
  wire [31:0] exp_291;
  wire [0:0] exp_297;
  wire [0:0] exp_196;
  wire [0:0] exp_191;
  wire [0:0] exp_188;
  wire [31:0] exp_187;
  wire [0:0] exp_190;
  wire [31:0] exp_189;
  wire [0:0] exp_195;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [31:0] exp_146;
  wire [0:0] exp_149;
  wire [31:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [14:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_397;
  wire [0:0] exp_682;
  wire [0:0] exp_681;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_176;
  wire [0:0] exp_183;
  wire [0:0] exp_285;
  wire [0:0] exp_303;
  wire [0:0] exp_308;
  wire [0:0] exp_378;
  wire [0:0] exp_383;
  wire [0:0] exp_380;
  wire [0:0] exp_379;
  wire [0:0] exp_352;
  wire [0:0] exp_376;
  wire [0:0] exp_372;
  wire [0:0] exp_336;
  wire [0:0] exp_350;
  wire [0:0] exp_347;
  wire [0:0] exp_332;
  wire [0:0] exp_334;
  wire [0:0] exp_330;
  wire [0:0] exp_384;
  wire [0:0] exp_323;
  wire [0:0] exp_309;
  wire [0:0] exp_317;
  wire [0:0] exp_322;
  wire [0:0] exp_310;
  wire [0:0] exp_333;
  wire [0:0] exp_329;
  wire [0:0] exp_327;
  wire [0:0] exp_325;
  wire [0:0] exp_304;
  wire [0:0] exp_324;
  wire [0:0] exp_326;
  wire [0:0] exp_328;
  wire [0:0] exp_331;
  wire [0:0] exp_346;
  wire [0:0] exp_349;
  wire [0:0] exp_348;
  wire [0:0] exp_345;
  wire [0:0] exp_339;
  wire [9:0] exp_337;
  wire [9:0] exp_344;
  wire [0:0] exp_343;
  wire [9:0] exp_341;
  wire [0:0] exp_340;
  wire [0:0] exp_342;
  wire [9:0] exp_338;
  wire [0:0] exp_335;
  wire [0:0] exp_375;
  wire [0:0] exp_374;
  wire [0:0] exp_373;
  wire [0:0] exp_361;
  wire [0:0] exp_355;
  wire [8:0] exp_353;
  wire [8:0] exp_360;
  wire [0:0] exp_359;
  wire [8:0] exp_357;
  wire [0:0] exp_356;
  wire [0:0] exp_358;
  wire [8:0] exp_354;
  wire [0:0] exp_371;
  wire [0:0] exp_365;
  wire [2:0] exp_363;
  wire [2:0] exp_370;
  wire [0:0] exp_369;
  wire [2:0] exp_367;
  wire [0:0] exp_366;
  wire [0:0] exp_368;
  wire [0:0] exp_362;
  wire [2:0] exp_364;
  wire [0:0] exp_351;
  wire [0:0] exp_382;
  wire [0:0] exp_381;
  wire [0:0] exp_377;
  wire [0:0] exp_992;
  wire [0:0] exp_991;
  wire [0:0] exp_406;
  wire [0:0] exp_449;
  wire [31:0] exp_421;
  wire [0:0] exp_420;
  wire [1:0] exp_429;
  wire [4:0] exp_416;
  wire [0:0] exp_419;
  wire [0:0] exp_998;
  wire [0:0] exp_997;
  wire [4:0] exp_415;
  wire [31:0] exp_417;
  wire [31:0] exp_994;
  wire [0:0] exp_993;
  wire [31:0] exp_630;
  wire [0:0] exp_629;
  wire [31:0] exp_581;
  wire [2:0] exp_524;
  wire [2:0] exp_515;
  wire [0:0] exp_512;
  wire [0:0] exp_446;
  wire [6:0] exp_436;
  wire [6:0] exp_445;
  wire [0:0] exp_448;
  wire [6:0] exp_447;
  wire [0:0] exp_514;
  wire [2:0] exp_502;
  wire [0:0] exp_444;
  wire [4:0] exp_443;
  wire [0:0] exp_501;
  wire [2:0] exp_489;
  wire [0:0] exp_442;
  wire [5:0] exp_441;
  wire [0:0] exp_488;
  wire [2:0] exp_438;
  wire [0:0] exp_487;
  wire [0:0] exp_500;
  wire [0:0] exp_513;
  wire [0:0] exp_519;
  wire [0:0] exp_580;
  wire [31:0] exp_560;
  wire [0:0] exp_526;
  wire [0:0] exp_518;
  wire [0:0] exp_504;
  wire [0:0] exp_491;
  wire [0:0] exp_477;
  wire [0:0] exp_475;
  wire [0:0] exp_476;
  wire [0:0] exp_440;
  wire [4:0] exp_439;
  wire [0:0] exp_490;
  wire [0:0] exp_503;
  wire [0:0] exp_517;
  wire [0:0] exp_516;
  wire [0:0] exp_559;
  wire [31:0] exp_557;
  wire [31:0] exp_522;
  wire [31:0] exp_508;
  wire [0:0] exp_505;
  wire [0:0] exp_507;
  wire [31:0] exp_497;
  wire [0:0] exp_496;
  wire [31:0] exp_483;
  wire [0:0] exp_482;
  wire [31:0] exp_481;
  wire [31:0] exp_479;
  wire [19:0] exp_478;
  wire [3:0] exp_480;
  wire [31:0] exp_495;
  wire [31:0] exp_493;
  wire [19:0] exp_492;
  wire [3:0] exp_494;
  wire [31:0] exp_506;
  wire [31:0] exp_523;
  wire [31:0] exp_511;
  wire [0:0] exp_509;
  wire [0:0] exp_510;
  wire [31:0] exp_499;
  wire [0:0] exp_498;
  wire [31:0] exp_486;
  wire [0:0] exp_485;
  wire [31:0] exp_470;
  wire [0:0] exp_469;
  wire [31:0] exp_464;
  wire [0:0] exp_460;
  wire [4:0] exp_435;
  wire [0:0] exp_459;
  wire [0:0] exp_463;
  wire [31:0] exp_452;
  wire [0:0] exp_432;
  wire [0:0] exp_1008;
  wire [0:0] exp_1007;
  wire [0:0] exp_1006;
  wire [0:0] exp_1005;
  wire [4:0] exp_414;
  wire [0:0] exp_451;
  wire [31:0] exp_428;
  wire [0:0] exp_427;
  wire [1:0] exp_430;
  wire [4:0] exp_423;
  wire [0:0] exp_426;
  wire [0:0] exp_1000;
  wire [0:0] exp_999;
  wire [4:0] exp_422;
  wire [31:0] exp_424;
  wire [31:0] exp_433;
  wire [31:0] exp_462;
  wire [0:0] exp_461;
  wire [31:0] exp_468;
  wire [31:0] exp_465;
  wire [31:0] exp_467;
  wire [11:0] exp_466;
  wire [31:0] exp_484;
  wire [31:0] exp_412;
  wire [0:0] exp_411;
  wire [31:0] exp_558;
  wire [31:0] exp_562;
  wire [31:0] exp_561;
  wire [5:0] exp_556;
  wire [5:0] exp_555;
  wire [5:0] exp_554;
  wire [4:0] exp_525;
  wire [4:0] exp_474;
  wire [0:0] exp_473;
  wire [4:0] exp_472;
  wire [4:0] exp_437;
  wire [31:0] exp_578;
  wire [1:0] exp_564;
  wire [0:0] exp_563;
  wire [31:0] exp_579;
  wire [1:0] exp_570;
  wire [0:0] exp_569;
  wire [31:0] exp_566;
  wire [31:0] exp_565;
  wire [31:0] exp_568;
  wire [31:0] exp_567;
  wire [31:0] exp_571;
  wire [31:0] exp_575;
  wire [32:0] exp_574;
  wire [32:0] exp_572;
  wire [0:0] exp_553;
  wire [0:0] exp_527;
  wire [0:0] exp_471;
  wire [0:0] exp_552;
  wire [0:0] exp_551;
  wire [0:0] exp_550;
  wire [32:0] exp_573;
  wire [31:0] exp_576;
  wire [31:0] exp_577;
  wire [31:0] exp_628;
  wire [0:0] exp_627;
  wire [31:0] exp_618;
  wire [7:0] exp_617;
  wire [7:0] exp_616;
  wire [7:0] exp_611;
  wire [1:0] exp_602;
  wire [1:0] exp_601;
  wire [1:0] exp_600;
  wire [0:0] exp_610;
  wire [7:0] exp_606;
  wire [31:0] exp_394;
  wire [31:0] exp_319;
  wire [0:0] exp_318;
  wire [31:0] exp_296;
  wire [0:0] exp_295;
  wire [31:0] exp_194;
  wire [0:0] exp_193;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [12:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_398;
  wire [3:0] exp_679;
  wire [0:0] exp_678;
  wire [3:0] exp_666;
  wire [3:0] exp_662;
  wire [1:0] exp_665;
  wire [1:0] exp_664;
  wire [1:0] exp_663;
  wire [3:0] exp_671;
  wire [3:0] exp_667;
  wire [0:0] exp_670;
  wire [0:0] exp_669;
  wire [0:0] exp_668;
  wire [3:0] exp_672;
  wire [3:0] exp_673;
  wire [3:0] exp_674;
  wire [3:0] exp_675;
  wire [3:0] exp_676;
  wire [3:0] exp_677;
  wire [12:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_393;
  wire [31:0] exp_661;
  wire [0:0] exp_660;
  wire [31:0] exp_648;
  wire [0:0] exp_647;
  wire [31:0] exp_634;
  wire [7:0] exp_633;
  wire [7:0] exp_632;
  wire [7:0] exp_631;
  wire [31:0] exp_521;
  wire [31:0] exp_642;
  wire [3:0] exp_641;
  wire [31:0] exp_644;
  wire [4:0] exp_643;
  wire [31:0] exp_646;
  wire [4:0] exp_645;
  wire [31:0] exp_652;
  wire [0:0] exp_605;
  wire [0:0] exp_604;
  wire [0:0] exp_603;
  wire [0:0] exp_651;
  wire [31:0] exp_638;
  wire [15:0] exp_637;
  wire [15:0] exp_636;
  wire [15:0] exp_635;
  wire [31:0] exp_650;
  wire [4:0] exp_649;
  wire [31:0] exp_654;
  wire [31:0] exp_653;
  wire [31:0] exp_640;
  wire [31:0] exp_639;
  wire [31:0] exp_655;
  wire [31:0] exp_656;
  wire [31:0] exp_657;
  wire [31:0] exp_658;
  wire [31:0] exp_659;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [12:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [12:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [12:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [12:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [12:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [12:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [12:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [12:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [12:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [12:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [12:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [12:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_179;
  wire [0:0] exp_177;
  wire [31:0] exp_139;
  wire [0:0] exp_178;
  wire [31:0] exp_157;
  wire [31:0] exp_164;
  wire [0:0] exp_159;
  wire [31:0] exp_158;
  wire [0:0] exp_163;
  wire [31:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [31:0] exp_167;
  wire [31:0] exp_174;
  wire [0:0] exp_169;
  wire [31:0] exp_168;
  wire [0:0] exp_173;
  wire [31:0] exp_171;
  wire [0:0] exp_170;
  wire [0:0] exp_172;
  wire [0:0] exp_166;
  wire [0:0] exp_165;
  wire [31:0] exp_182;
  wire [31:0] exp_281;
  wire [31:0] exp_284;
  wire [31:0] exp_302;
  wire [31:0] exp_307;
  wire [31:0] exp_391;
  wire [7:0] exp_388;
  wire [7:0] exp_390;
  wire [6:0] exp_389;
  wire [0:0] exp_387;
  wire [0:0] exp_386;
  wire [0:0] exp_385;
  wire [7:0] exp_607;
  wire [7:0] exp_608;
  wire [7:0] exp_609;
  wire [31:0] exp_621;
  wire [15:0] exp_620;
  wire [15:0] exp_619;
  wire [15:0] exp_615;
  wire [0:0] exp_614;
  wire [15:0] exp_612;
  wire [15:0] exp_613;
  wire [31:0] exp_622;
  wire [31:0] exp_623;
  wire [31:0] exp_624;
  wire [31:0] exp_625;
  wire [31:0] exp_626;
  wire [31:0] exp_985;
  wire [0:0] exp_984;
  wire [31:0] exp_981;
  wire [0:0] exp_752;
  wire [0:0] exp_751;
  wire [0:0] exp_750;
  wire [0:0] exp_980;
  wire [31:0] exp_976;
  wire [63:0] exp_975;
  wire [0:0] exp_972;
  wire [0:0] exp_955;
  wire [0:0] exp_932;
  wire [0:0] exp_929;
  wire [0:0] exp_927;
  wire [0:0] exp_909;
  wire [0:0] exp_908;
  wire [0:0] exp_907;
  wire [31:0] exp_905;
  wire [0:0] exp_904;
  wire [0:0] exp_903;
  wire [0:0] exp_892;
  wire [0:0] exp_891;
  wire [0:0] exp_755;
  wire [0:0] exp_754;
  wire [0:0] exp_753;
  wire [0:0] exp_758;
  wire [0:0] exp_757;
  wire [1:0] exp_756;
  wire [0:0] exp_928;
  wire [0:0] exp_912;
  wire [0:0] exp_911;
  wire [0:0] exp_910;
  wire [31:0] exp_906;
  wire [0:0] exp_893;
  wire [0:0] exp_914;
  wire [0:0] exp_913;
  wire [0:0] exp_934;
  wire [1:0] exp_933;
  wire [0:0] exp_957;
  wire [1:0] exp_956;
  wire [0:0] exp_974;
  wire [63:0] exp_971;
  wire [63:0] exp_970;
  wire [63:0] exp_966;
  wire [63:0] exp_962;
  wire [63:0] exp_958;
  wire [31:0] exp_951;
  wire [31:0] exp_938;
  wire [31:0] exp_936;
  wire [15:0] exp_935;
  wire [31:0] exp_930;
  wire [31:0] exp_920;
  wire [31:0] exp_919;
  wire [31:0] exp_918;
  wire [0:0] exp_915;
  wire [0:0] exp_917;
  wire [31:0] exp_916;
  wire [15:0] exp_937;
  wire [31:0] exp_931;
  wire [31:0] exp_926;
  wire [31:0] exp_925;
  wire [31:0] exp_924;
  wire [0:0] exp_921;
  wire [0:0] exp_923;
  wire [31:0] exp_922;
  wire [63:0] exp_961;
  wire [63:0] exp_959;
  wire [31:0] exp_952;
  wire [31:0] exp_942;
  wire [31:0] exp_940;
  wire [15:0] exp_939;
  wire [15:0] exp_941;
  wire [4:0] exp_960;
  wire [63:0] exp_965;
  wire [63:0] exp_963;
  wire [31:0] exp_953;
  wire [31:0] exp_946;
  wire [31:0] exp_944;
  wire [15:0] exp_943;
  wire [15:0] exp_945;
  wire [4:0] exp_964;
  wire [63:0] exp_969;
  wire [63:0] exp_967;
  wire [31:0] exp_954;
  wire [31:0] exp_950;
  wire [31:0] exp_948;
  wire [15:0] exp_947;
  wire [15:0] exp_949;
  wire [5:0] exp_968;
  wire [63:0] exp_973;
  wire [31:0] exp_977;
  wire [31:0] exp_983;
  wire [0:0] exp_776;
  wire [0:0] exp_982;
  wire [31:0] exp_886;
  wire [31:0] exp_880;
  wire [0:0] exp_876;
  wire [0:0] exp_875;
  wire [31:0] exp_824;
  wire [31:0] exp_821;
  wire [31:0] exp_820;
  wire [31:0] exp_819;
  wire [0:0] exp_816;
  wire [0:0] exp_807;
  wire [0:0] exp_806;
  wire [0:0] exp_805;
  wire [31:0] exp_801;
  wire [0:0] exp_799;
  wire [0:0] exp_798;
  wire [0:0] exp_778;
  wire [0:0] exp_777;
  wire [0:0] exp_818;
  wire [31:0] exp_817;
  wire [0:0] exp_809;
  wire [0:0] exp_808;
  wire [0:0] exp_874;
  wire [0:0] exp_879;
  wire [31:0] exp_867;
  wire [31:0] exp_866;
  wire [31:0] exp_865;
  wire [0:0] exp_862;
  wire [0:0] exp_826;
  wire [0:0] exp_822;
  wire [0:0] exp_804;
  wire [0:0] exp_803;
  wire [0:0] exp_802;
  wire [31:0] exp_800;
  wire [0:0] exp_864;
  wire [31:0] exp_860;
  wire [31:0] exp_830;
  wire [31:0] exp_857;
  wire [0:0] exp_791;
  wire [1:0] exp_790;
  wire [0:0] exp_856;
  wire [31:0] exp_849;
  wire [0:0] exp_839;
  wire [0:0] exp_838;
  wire [32:0] exp_837;
  wire [32:0] exp_836;
  wire [32:0] exp_835;
  wire [31:0] exp_833;
  wire [31:0] exp_828;
  wire [32:0] exp_854;
  wire [0:0] exp_853;
  wire [32:0] exp_841;
  wire [0:0] exp_840;
  wire [0:0] exp_852;
  wire [0:0] exp_827;
  wire [0:0] exp_834;
  wire [31:0] exp_832;
  wire [31:0] exp_859;
  wire [0:0] exp_858;
  wire [31:0] exp_851;
  wire [0:0] exp_850;
  wire [31:0] exp_823;
  wire [31:0] exp_815;
  wire [31:0] exp_814;
  wire [31:0] exp_813;
  wire [0:0] exp_810;
  wire [0:0] exp_812;
  wire [31:0] exp_811;
  wire [0:0] exp_831;
  wire [0:0] exp_848;
  wire [31:0] exp_843;
  wire [0:0] exp_842;
  wire [31:0] exp_847;
  wire [31:0] exp_845;
  wire [0:0] exp_844;
  wire [0:0] exp_846;
  wire [0:0] exp_855;
  wire [0:0] exp_829;
  wire [0:0] exp_793;
  wire [5:0] exp_792;
  wire [31:0] exp_863;
  wire [31:0] exp_878;
  wire [0:0] exp_877;
  wire [0:0] exp_795;
  wire [5:0] exp_794;
  wire [31:0] exp_887;
  wire [31:0] exp_885;
  wire [0:0] exp_883;
  wire [0:0] exp_882;
  wire [0:0] exp_881;
  wire [0:0] exp_884;
  wire [31:0] exp_873;
  wire [31:0] exp_872;
  wire [31:0] exp_871;
  wire [0:0] exp_868;
  wire [0:0] exp_825;
  wire [0:0] exp_870;
  wire [31:0] exp_861;
  wire [31:0] exp_869;
  wire [31:0] exp_456;
  wire [0:0] exp_455;
  wire [0:0] exp_685;
  wire [0:0] exp_698;
  wire [0:0] exp_699;
  wire [0:0] exp_686;
  wire [0:0] exp_687;
  wire [0:0] exp_692;
  wire [31:0] exp_689;
  wire [31:0] exp_688;
  wire [31:0] exp_691;
  wire [31:0] exp_690;
  wire [0:0] exp_697;
  wire [31:0] exp_694;
  wire [31:0] exp_693;
  wire [31:0] exp_696;
  wire [31:0] exp_695;
  wire [0:0] exp_1012;
  wire [31:0] exp_1011;
  wire [2:0] exp_1010;
  wire [32:0] exp_742;
  wire [0:0] exp_741;
  wire [31:0] exp_732;
  wire [31:0] exp_731;
  wire [0:0] exp_730;
  wire [31:0] exp_717;
  wire [12:0] exp_716;
  wire [12:0] exp_715;
  wire [12:0] exp_714;
  wire [11:0] exp_713;
  wire [7:0] exp_712;
  wire [1:0] exp_711;
  wire [0:0] exp_706;
  wire [0:0] exp_707;
  wire [5:0] exp_708;
  wire [3:0] exp_709;
  wire [0:0] exp_710;
  wire [31:0] exp_729;
  wire [20:0] exp_728;
  wire [20:0] exp_727;
  wire [20:0] exp_726;
  wire [19:0] exp_725;
  wire [9:0] exp_724;
  wire [8:0] exp_723;
  wire [0:0] exp_718;
  wire [7:0] exp_719;
  wire [0:0] exp_720;
  wire [9:0] exp_721;
  wire [0:0] exp_722;
  wire [31:0] exp_529;
  wire [32:0] exp_740;
  wire [32:0] exp_739;
  wire [31:0] exp_737;
  wire [31:0] exp_736;
  wire [11:0] exp_735;
  wire [11:0] exp_734;
  wire [11:0] exp_733;
  wire [32:0] exp_738;
  wire [0:0] exp_409;
  wire [0:0] exp_80;
  wire [12:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_544;
  wire [0:0] exp_185;
  wire [0:0] exp_218;
  wire [0:0] exp_217;
  wire [0:0] exp_215;
  wire [0:0] exp_209;
  wire [8:0] exp_207;
  wire [8:0] exp_214;
  wire [0:0] exp_213;
  wire [8:0] exp_211;
  wire [0:0] exp_210;
  wire [0:0] exp_212;
  wire [8:0] exp_208;
  wire [0:0] exp_205;
  wire [0:0] exp_244;
  wire [0:0] exp_243;
  wire [0:0] exp_242;
  wire [0:0] exp_230;
  wire [0:0] exp_224;
  wire [8:0] exp_222;
  wire [8:0] exp_229;
  wire [0:0] exp_228;
  wire [8:0] exp_226;
  wire [0:0] exp_225;
  wire [0:0] exp_227;
  wire [8:0] exp_223;
  wire [0:0] exp_240;
  wire [0:0] exp_234;
  wire [2:0] exp_232;
  wire [2:0] exp_239;
  wire [0:0] exp_238;
  wire [2:0] exp_236;
  wire [0:0] exp_235;
  wire [0:0] exp_237;
  wire [0:0] exp_231;
  wire [2:0] exp_233;
  wire [0:0] exp_220;
  wire [0:0] exp_260;
  wire [0:0] exp_259;
  wire [0:0] exp_256;
  wire [0:0] exp_250;
  wire [8:0] exp_248;
  wire [8:0] exp_255;
  wire [0:0] exp_254;
  wire [8:0] exp_252;
  wire [0:0] exp_251;
  wire [0:0] exp_253;
  wire [8:0] exp_249;
  wire [0:0] exp_246;
  wire [0:0] exp_203;
  wire [0:0] exp_202;
  wire [0:0] exp_200;
  wire [0:0] exp_279;
  wire [0:0] exp_276;
  wire [0:0] exp_275;
  wire [0:0] exp_273;
  wire [7:0] exp_264;
  wire [7:0] exp_272;
  wire [0:0] exp_270;
  wire [0:0] exp_271;
  wire [7:0] exp_269;
  wire [0:0] exp_265;
  wire [0:0] exp_268;
  wire [7:0] exp_267;
  wire [0:0] exp_266;
  wire [7:0] exp_197;
  wire [31:0] exp_181;
  wire [0:0] exp_263;
  wire [0:0] exp_274;
  wire [0:0] exp_278;
  wire [31:0] exp_301;
  wire [31:0] exp_283;
  wire [0:0] exp_300;
  wire [0:0] exp_286;
  wire [0:0] exp_294;
  wire [0:0] exp_287;


  reg [0:0] exp_280_reg;
  always@(*) begin
    case (exp_277)
      0:exp_280_reg <= exp_276;
      1:exp_280_reg <= exp_278;
      default:exp_280_reg <= exp_279;
    endcase
  end
  assign exp_280 = exp_280_reg;
  assign exp_277 = exp_201 | exp_247;

      reg [0:0] exp_201_reg = 1;
      always@(posedge clk) begin
        if (exp_200) begin
          exp_201_reg <= exp_204;
        end
      end
      assign exp_201 = exp_201_reg;
      assign exp_204 = exp_199 | exp_203;
  assign exp_199 = exp_262;
  assign exp_262 = exp_247 & exp_256;

      reg [0:0] exp_247_reg = 0;
      always@(posedge clk) begin
        if (exp_246) begin
          exp_247_reg <= exp_261;
        end
      end
      assign exp_247 = exp_247_reg;
      assign exp_261 = exp_258 | exp_260;
  assign exp_258 = exp_257 & exp_240;
  assign exp_257 = exp_221 & exp_230;

      reg [0:0] exp_221_reg = 0;
      always@(posedge clk) begin
        if (exp_220) begin
          exp_221_reg <= exp_245;
        end
      end
      assign exp_221 = exp_221_reg;
      assign exp_245 = exp_241 | exp_244;
  assign exp_241 = exp_206 & exp_215;

      reg [0:0] exp_206_reg = 0;
      always@(posedge clk) begin
        if (exp_205) begin
          exp_206_reg <= exp_219;
        end
      end
      assign exp_206 = exp_206_reg;
      assign exp_219 = exp_216 | exp_218;
  assign exp_216 = exp_201 & exp_198;
  assign exp_198 = exp_184 & exp_185;
  assign exp_184 = exp_192;
  assign exp_192 = exp_5 & exp_191;
  assign exp_5 = exp_396;
  assign exp_396 = exp_743;
  assign exp_743 = exp_680 & exp_408;
  assign exp_680 = exp_545 | exp_547;
  assign exp_545 = exp_530 == exp_544;
  assign exp_530 = exp_528[6:0];

      reg [31:0] exp_528_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_528_reg <= exp_96;
        end
      end
      assign exp_528 = exp_528_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_410;

      reg [31:0] exp_410_reg = 0;
      always@(posedge clk) begin
        if (exp_409) begin
          exp_410_reg <= exp_1013;
        end
      end
      assign exp_410 = exp_410_reg;
    
  reg [32:0] exp_1013_reg;
  always@(*) begin
    case (exp_1009)
      0:exp_1013_reg <= exp_1011;
      1:exp_1013_reg <= exp_742;
      default:exp_1013_reg <= exp_1012;
    endcase
  end
  assign exp_1013 = exp_1013_reg;
  assign exp_1009 = exp_705 & exp_408;
  assign exp_705 = exp_683 | exp_704;
  assign exp_683 = exp_541 | exp_543;
  assign exp_541 = exp_530 == exp_540;
  assign exp_540 = 111;
  assign exp_543 = exp_530 == exp_542;
  assign exp_542 = 103;

  reg [0:0] exp_704_reg;
  always@(*) begin
    case (exp_549)
      0:exp_704_reg <= exp_702;
      1:exp_704_reg <= exp_701;
      default:exp_704_reg <= exp_703;
    endcase
  end
  assign exp_704 = exp_704_reg;
  assign exp_549 = exp_530 == exp_548;
  assign exp_548 = 99;
  assign exp_703 = 0;
  assign exp_702 = 0;

  reg [0:0] exp_701_reg;
  always@(*) begin
    case (exp_531)
      0:exp_701_reg <= exp_684;
      1:exp_701_reg <= exp_685;
      2:exp_701_reg <= exp_698;
      3:exp_701_reg <= exp_699;
      4:exp_701_reg <= exp_686;
      5:exp_701_reg <= exp_687;
      6:exp_701_reg <= exp_692;
      7:exp_701_reg <= exp_697;
      default:exp_701_reg <= exp_700;
    endcase
  end
  assign exp_701 = exp_701_reg;
  assign exp_531 = exp_528[14:12];
  assign exp_700 = 0;
  assign exp_684 = exp_520 == exp_521;

      reg [31:0] exp_520_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_520_reg <= exp_458;
        end
      end
      assign exp_520 = exp_520_reg;
    
  reg [31:0] exp_458_reg;
  always@(*) begin
    case (exp_454)
      0:exp_458_reg <= exp_450;
      1:exp_458_reg <= exp_456;
      default:exp_458_reg <= exp_457;
    endcase
  end
  assign exp_458 = exp_458_reg;
  assign exp_454 = exp_434 == exp_453;
  assign exp_434 = exp_96[19:15];
  assign exp_453 = 0;
  assign exp_457 = 0;

  reg [31:0] exp_450_reg;
  always@(*) begin
    case (exp_431)
      0:exp_450_reg <= exp_421;
      1:exp_450_reg <= exp_433;
      default:exp_450_reg <= exp_449;
    endcase
  end
  assign exp_450 = exp_450_reg;
  assign exp_431 = exp_1004;
  assign exp_1004 = exp_1003 & exp_400;
  assign exp_1003 = exp_1002 & exp_408;
  assign exp_1002 = exp_1001 & exp_995;
  assign exp_1001 = exp_413 == exp_996;
  assign exp_413 = exp_96[19:15];
  assign exp_996 = exp_528[11:7];
  assign exp_995 = exp_587 | exp_990;
  assign exp_587 = exp_586 | exp_545;
  assign exp_586 = exp_585 | exp_539;
  assign exp_585 = exp_584 | exp_537;
  assign exp_584 = exp_583 | exp_543;
  assign exp_583 = exp_582 | exp_541;
  assign exp_582 = exp_533 | exp_535;
  assign exp_533 = exp_530 == exp_532;
  assign exp_532 = 19;
  assign exp_535 = exp_530 == exp_534;
  assign exp_534 = 51;
  assign exp_537 = exp_530 == exp_536;
  assign exp_536 = 55;
  assign exp_539 = exp_530 == exp_538;
  assign exp_538 = 23;
  assign exp_990 = exp_989 & exp_749;

  reg [0:0] exp_989_reg;
  always@(*) begin
    case (exp_775)
      0:exp_989_reg <= exp_986;
      1:exp_989_reg <= exp_987;
      default:exp_989_reg <= exp_988;
    endcase
  end
  assign exp_989 = exp_989_reg;
  assign exp_775 = exp_749 & exp_774;
  assign exp_749 = exp_747 & exp_748;
  assign exp_747 = exp_745 == exp_746;
  assign exp_745 = exp_528[6:0];
  assign exp_746 = 51;
  assign exp_748 = exp_528[25:25];
  assign exp_774 = exp_744[2:2];
  assign exp_744 = exp_528[14:12];
  assign exp_988 = 0;
  assign exp_986 = exp_979 & exp_749;
  assign exp_979 = exp_894 == exp_978;

      reg [2:0] exp_894_reg = 0;
      always@(posedge clk) begin
        if (exp_890) begin
          exp_894_reg <= exp_901;
        end
      end
      assign exp_894 = exp_894_reg;
    
  reg [2:0] exp_901_reg;
  always@(*) begin
    case (exp_896)
      0:exp_901_reg <= exp_898;
      1:exp_901_reg <= exp_899;
      default:exp_901_reg <= exp_900;
    endcase
  end
  assign exp_901 = exp_901_reg;
  assign exp_896 = exp_894 == exp_895;
  assign exp_895 = 4;
  assign exp_900 = 0;
  assign exp_898 = exp_894 + exp_897;
  assign exp_897 = 1;
  assign exp_899 = 0;
  assign exp_890 = exp_749 & exp_889;
  assign exp_889 = ~exp_888;
  assign exp_888 = exp_744[2:2];
  assign exp_978 = 4;
  assign exp_987 = exp_797 & exp_749;
  assign exp_797 = exp_781 == exp_796;

      reg [5:0] exp_781_reg = 0;
      always@(posedge clk) begin
        if (exp_775) begin
          exp_781_reg <= exp_788;
        end
      end
      assign exp_781 = exp_781_reg;
    
  reg [5:0] exp_788_reg;
  always@(*) begin
    case (exp_783)
      0:exp_788_reg <= exp_785;
      1:exp_788_reg <= exp_786;
      default:exp_788_reg <= exp_787;
    endcase
  end
  assign exp_788 = exp_788_reg;
  assign exp_783 = exp_781 == exp_782;
  assign exp_782 = 37;
  assign exp_787 = 0;
  assign exp_785 = exp_781 + exp_784;
  assign exp_784 = 1;
  assign exp_786 = 0;
  assign exp_796 = 37;

      reg [0:0] exp_408_reg = 0;
      always@(posedge clk) begin
        if (exp_400) begin
          exp_408_reg <= exp_407;
        end
      end
      assign exp_408 = exp_408_reg;
      assign exp_407 = exp_405 & exp_406;

      reg [0:0] exp_405_reg = 0;
      always@(posedge clk) begin
        if (exp_400) begin
          exp_405_reg <= exp_404;
        end
      end
      assign exp_405 = exp_405_reg;
      assign exp_404 = exp_402 & exp_403;
  assign exp_402 = 1;
  assign exp_403 = ~exp_401;
  assign exp_401 = exp_1014;
  assign exp_1014 = exp_408 & exp_705;
  assign exp_400 = ~exp_399;
  assign exp_399 = exp_1018;
  assign exp_1018 = exp_408 & exp_1017;
  assign exp_1017 = exp_1016 | exp_992;
  assign exp_1016 = exp_396 & exp_1015;
  assign exp_1015 = ~exp_395;
  assign exp_395 = exp_321;

  reg [0:0] exp_321_reg;
  always@(*) begin
    case (exp_316)
      0:exp_321_reg <= exp_298;
      1:exp_321_reg <= exp_308;
      default:exp_321_reg <= exp_320;
    endcase
  end
  assign exp_321 = exp_321_reg;
  assign exp_316 = exp_313 & exp_315;
  assign exp_313 = exp_1 >= exp_312;
  assign exp_1 = exp_392;
  assign exp_392 = exp_599;
  assign exp_599 = exp_598 + exp_597;
  assign exp_598 = 0;
  assign exp_597 = exp_520 + exp_596;
  assign exp_596 = $signed(exp_595);
  assign exp_595 = exp_594 + exp_593;
  assign exp_594 = 0;

  reg [11:0] exp_593_reg;
  always@(*) begin
    case (exp_547)
      0:exp_593_reg <= exp_588;
      1:exp_593_reg <= exp_591;
      default:exp_593_reg <= exp_592;
    endcase
  end
  assign exp_593 = exp_593_reg;
  assign exp_547 = exp_530 == exp_546;
  assign exp_546 = 35;
  assign exp_592 = 0;
  assign exp_588 = exp_528[31:20];
  assign exp_591 = {exp_589, exp_590};  assign exp_589 = exp_528[31:25];
  assign exp_590 = exp_528[11:7];
  assign exp_312 = 2147483664;
  assign exp_315 = exp_1 <= exp_314;
  assign exp_314 = 2147483664;
  assign exp_320 = 0;

  reg [0:0] exp_298_reg;
  always@(*) begin
    case (exp_293)
      0:exp_298_reg <= exp_196;
      1:exp_298_reg <= exp_285;
      default:exp_298_reg <= exp_297;
    endcase
  end
  assign exp_298 = exp_298_reg;
  assign exp_293 = exp_290 & exp_292;
  assign exp_290 = exp_1 >= exp_289;
  assign exp_289 = 2147483660;
  assign exp_292 = exp_1 <= exp_291;
  assign exp_291 = 2147483660;
  assign exp_297 = 0;

  reg [0:0] exp_196_reg;
  always@(*) begin
    case (exp_191)
      0:exp_196_reg <= exp_155;
      1:exp_196_reg <= exp_183;
      default:exp_196_reg <= exp_195;
    endcase
  end
  assign exp_196 = exp_196_reg;
  assign exp_191 = exp_188 & exp_190;
  assign exp_188 = exp_1 >= exp_187;
  assign exp_187 = 2147483656;
  assign exp_190 = exp_1 <= exp_189;
  assign exp_189 = 2147483656;
  assign exp_195 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 2147483648;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 2147483652;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 20476;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_397;
  assign exp_397 = exp_682;
  assign exp_682 = exp_681 + exp_547;
  assign exp_681 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_176;
  assign exp_176 = 1;
  assign exp_183 = exp_201;
  assign exp_285 = exp_303;
  assign exp_303 = 1;
  assign exp_308 = exp_378;

      reg [0:0] exp_378_reg = 0;
      always@(posedge clk) begin
        if (exp_377) begin
          exp_378_reg <= exp_383;
        end
      end
      assign exp_378 = exp_378_reg;
      assign exp_383 = exp_380 | exp_382;
  assign exp_380 = exp_379 & exp_371;
  assign exp_379 = exp_352 & exp_361;

      reg [0:0] exp_352_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_352_reg <= exp_376;
        end
      end
      assign exp_352 = exp_352_reg;
      assign exp_376 = exp_372 | exp_375;
  assign exp_372 = exp_336 & exp_345;

      reg [0:0] exp_336_reg = 0;
      always@(posedge clk) begin
        if (exp_335) begin
          exp_336_reg <= exp_350;
        end
      end
      assign exp_336 = exp_336_reg;
      assign exp_350 = exp_347 | exp_349;
  assign exp_347 = exp_332 & exp_346;

      reg [0:0] exp_332_reg = 1;
      always@(posedge clk) begin
        if (exp_331) begin
          exp_332_reg <= exp_334;
        end
      end
      assign exp_332 = exp_332_reg;
      assign exp_334 = exp_330 | exp_333;
  assign exp_330 = exp_384;
  assign exp_384 = exp_378 & exp_323;
  assign exp_323 = exp_309 & exp_322;
  assign exp_309 = exp_317;
  assign exp_317 = exp_5 & exp_316;
  assign exp_322 = ~exp_310;
  assign exp_310 = exp_6;
  assign exp_333 = exp_332 & exp_329;

      reg [0:0] exp_329_reg = 1;
      always@(posedge clk) begin
        if (exp_328) begin
          exp_329_reg <= exp_327;
        end
      end
      assign exp_329 = exp_329_reg;
    
      reg [0:0] exp_327_reg = 1;
      always@(posedge clk) begin
        if (exp_326) begin
          exp_327_reg <= exp_325;
        end
      end
      assign exp_327 = exp_327_reg;
    
      reg [0:0] exp_325_reg = 1;
      always@(posedge clk) begin
        if (exp_324) begin
          exp_325_reg <= exp_304;
        end
      end
      assign exp_325 = exp_325_reg;
      assign exp_304 = stdin_rx;
  assign exp_324 = 1;
  assign exp_326 = 1;
  assign exp_328 = 1;
  assign exp_331 = 1;
  assign exp_346 = ~exp_329;
  assign exp_349 = exp_336 & exp_348;
  assign exp_348 = ~exp_345;
  assign exp_345 = exp_339 & exp_336;
  assign exp_339 = exp_337 == exp_338;

      reg [9:0] exp_337_reg = 0;
      always@(posedge clk) begin
        if (exp_336) begin
          exp_337_reg <= exp_344;
        end
      end
      assign exp_337 = exp_337_reg;
    
  reg [9:0] exp_344_reg;
  always@(*) begin
    case (exp_339)
      0:exp_344_reg <= exp_341;
      1:exp_344_reg <= exp_342;
      default:exp_344_reg <= exp_343;
    endcase
  end
  assign exp_344 = exp_344_reg;
  assign exp_343 = 0;
  assign exp_341 = exp_337 + exp_340;
  assign exp_340 = 1;
  assign exp_342 = 0;
  assign exp_338 = 649;
  assign exp_335 = 1;
  assign exp_375 = exp_352 & exp_374;
  assign exp_374 = ~exp_373;
  assign exp_373 = exp_361 & exp_371;
  assign exp_361 = exp_355 & exp_352;
  assign exp_355 = exp_353 == exp_354;

      reg [8:0] exp_353_reg = 0;
      always@(posedge clk) begin
        if (exp_352) begin
          exp_353_reg <= exp_360;
        end
      end
      assign exp_353 = exp_353_reg;
    
  reg [8:0] exp_360_reg;
  always@(*) begin
    case (exp_355)
      0:exp_360_reg <= exp_357;
      1:exp_360_reg <= exp_358;
      default:exp_360_reg <= exp_359;
    endcase
  end
  assign exp_360 = exp_360_reg;
  assign exp_359 = 0;
  assign exp_357 = exp_353 + exp_356;
  assign exp_356 = 1;
  assign exp_358 = 0;
  assign exp_354 = 433;
  assign exp_371 = exp_365 & exp_362;
  assign exp_365 = exp_363 == exp_364;

      reg [2:0] exp_363_reg = 0;
      always@(posedge clk) begin
        if (exp_362) begin
          exp_363_reg <= exp_370;
        end
      end
      assign exp_363 = exp_363_reg;
    
  reg [2:0] exp_370_reg;
  always@(*) begin
    case (exp_365)
      0:exp_370_reg <= exp_367;
      1:exp_370_reg <= exp_368;
      default:exp_370_reg <= exp_369;
    endcase
  end
  assign exp_370 = exp_370_reg;
  assign exp_369 = 0;
  assign exp_367 = exp_363 + exp_366;
  assign exp_366 = 1;
  assign exp_368 = 0;
  assign exp_362 = exp_352 & exp_361;
  assign exp_364 = 7;
  assign exp_351 = 1;
  assign exp_382 = exp_378 & exp_381;
  assign exp_381 = ~exp_323;
  assign exp_377 = 1;
  assign exp_992 = exp_749 & exp_991;
  assign exp_991 = ~exp_989;
  assign exp_406 = ~exp_401;
  assign exp_449 = 0;

  //Create RAM
  reg [31:0] exp_421_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_419) begin
      exp_421_ram[exp_415] <= exp_417;
    end
  end
  assign exp_421 = exp_421_ram[exp_416];
  assign exp_420 = exp_429;
  assign exp_429 = 1;
  assign exp_416 = exp_413;
  assign exp_419 = exp_998;
  assign exp_998 = exp_997 & exp_400;
  assign exp_997 = exp_995 & exp_408;
  assign exp_415 = exp_996;
  assign exp_417 = exp_994;

  reg [31:0] exp_994_reg;
  always@(*) begin
    case (exp_990)
      0:exp_994_reg <= exp_630;
      1:exp_994_reg <= exp_985;
      default:exp_994_reg <= exp_993;
    endcase
  end
  assign exp_994 = exp_994_reg;
  assign exp_993 = 0;

  reg [31:0] exp_630_reg;
  always@(*) begin
    case (exp_545)
      0:exp_630_reg <= exp_581;
      1:exp_630_reg <= exp_628;
      default:exp_630_reg <= exp_629;
    endcase
  end
  assign exp_630 = exp_630_reg;
  assign exp_629 = 0;

  reg [31:0] exp_581_reg;
  always@(*) begin
    case (exp_524)
      0:exp_581_reg <= exp_560;
      1:exp_581_reg <= exp_562;
      2:exp_581_reg <= exp_578;
      3:exp_581_reg <= exp_579;
      4:exp_581_reg <= exp_571;
      5:exp_581_reg <= exp_575;
      6:exp_581_reg <= exp_576;
      7:exp_581_reg <= exp_577;
      default:exp_581_reg <= exp_580;
    endcase
  end
  assign exp_581 = exp_581_reg;

      reg [2:0] exp_524_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_524_reg <= exp_515;
        end
      end
      assign exp_524 = exp_524_reg;
    
  reg [2:0] exp_515_reg;
  always@(*) begin
    case (exp_512)
      0:exp_515_reg <= exp_502;
      1:exp_515_reg <= exp_513;
      default:exp_515_reg <= exp_514;
    endcase
  end
  assign exp_515 = exp_515_reg;
  assign exp_512 = exp_446 | exp_448;
  assign exp_446 = exp_436 == exp_445;
  assign exp_436 = exp_96[6:0];
  assign exp_445 = 111;
  assign exp_448 = exp_436 == exp_447;
  assign exp_447 = 103;
  assign exp_514 = 0;

  reg [2:0] exp_502_reg;
  always@(*) begin
    case (exp_444)
      0:exp_502_reg <= exp_489;
      1:exp_502_reg <= exp_500;
      default:exp_502_reg <= exp_501;
    endcase
  end
  assign exp_502 = exp_502_reg;
  assign exp_444 = exp_436 == exp_443;
  assign exp_443 = 23;
  assign exp_501 = 0;

  reg [2:0] exp_489_reg;
  always@(*) begin
    case (exp_442)
      0:exp_489_reg <= exp_438;
      1:exp_489_reg <= exp_487;
      default:exp_489_reg <= exp_488;
    endcase
  end
  assign exp_489 = exp_489_reg;
  assign exp_442 = exp_436 == exp_441;
  assign exp_441 = 55;
  assign exp_488 = 0;
  assign exp_438 = exp_96[14:12];
  assign exp_487 = 0;
  assign exp_500 = 0;
  assign exp_513 = 0;
  assign exp_519 = exp_400 & exp_405;
  assign exp_580 = 0;

  reg [31:0] exp_560_reg;
  always@(*) begin
    case (exp_526)
      0:exp_560_reg <= exp_557;
      1:exp_560_reg <= exp_558;
      default:exp_560_reg <= exp_559;
    endcase
  end
  assign exp_560 = exp_560_reg;

      reg [0:0] exp_526_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_526_reg <= exp_518;
        end
      end
      assign exp_526 = exp_526_reg;
      assign exp_518 = exp_504 & exp_517;
  assign exp_504 = exp_491 & exp_503;
  assign exp_491 = exp_477 & exp_490;
  assign exp_477 = exp_475 & exp_476;
  assign exp_475 = exp_96[30:30];
  assign exp_476 = ~exp_440;
  assign exp_440 = exp_436 == exp_439;
  assign exp_439 = 19;
  assign exp_490 = ~exp_442;
  assign exp_503 = ~exp_444;
  assign exp_517 = ~exp_516;
  assign exp_516 = exp_446 | exp_448;
  assign exp_559 = 0;
  assign exp_557 = exp_522 + exp_523;

      reg [31:0] exp_522_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_522_reg <= exp_508;
        end
      end
      assign exp_522 = exp_522_reg;
    
  reg [31:0] exp_508_reg;
  always@(*) begin
    case (exp_505)
      0:exp_508_reg <= exp_497;
      1:exp_508_reg <= exp_506;
      default:exp_508_reg <= exp_507;
    endcase
  end
  assign exp_508 = exp_508_reg;
  assign exp_505 = exp_446 | exp_448;
  assign exp_507 = 0;

  reg [31:0] exp_497_reg;
  always@(*) begin
    case (exp_444)
      0:exp_497_reg <= exp_483;
      1:exp_497_reg <= exp_495;
      default:exp_497_reg <= exp_496;
    endcase
  end
  assign exp_497 = exp_497_reg;
  assign exp_496 = 0;

  reg [31:0] exp_483_reg;
  always@(*) begin
    case (exp_442)
      0:exp_483_reg <= exp_458;
      1:exp_483_reg <= exp_481;
      default:exp_483_reg <= exp_482;
    endcase
  end
  assign exp_483 = exp_483_reg;
  assign exp_482 = 0;
  assign exp_481 = exp_479 << exp_480;
  assign exp_479 = exp_478;
  assign exp_478 = exp_96[31:12];
  assign exp_480 = 12;
  assign exp_495 = exp_493 << exp_494;
  assign exp_493 = exp_492;
  assign exp_492 = exp_96[31:12];
  assign exp_494 = 12;
  assign exp_506 = 4;

      reg [31:0] exp_523_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_523_reg <= exp_511;
        end
      end
      assign exp_523 = exp_523_reg;
    
  reg [31:0] exp_511_reg;
  always@(*) begin
    case (exp_509)
      0:exp_511_reg <= exp_499;
      1:exp_511_reg <= exp_412;
      default:exp_511_reg <= exp_510;
    endcase
  end
  assign exp_511 = exp_511_reg;
  assign exp_509 = exp_446 | exp_448;
  assign exp_510 = 0;

  reg [31:0] exp_499_reg;
  always@(*) begin
    case (exp_444)
      0:exp_499_reg <= exp_486;
      1:exp_499_reg <= exp_412;
      default:exp_499_reg <= exp_498;
    endcase
  end
  assign exp_499 = exp_499_reg;
  assign exp_498 = 0;

  reg [31:0] exp_486_reg;
  always@(*) begin
    case (exp_442)
      0:exp_486_reg <= exp_470;
      1:exp_486_reg <= exp_484;
      default:exp_486_reg <= exp_485;
    endcase
  end
  assign exp_486 = exp_486_reg;
  assign exp_485 = 0;

  reg [31:0] exp_470_reg;
  always@(*) begin
    case (exp_440)
      0:exp_470_reg <= exp_464;
      1:exp_470_reg <= exp_468;
      default:exp_470_reg <= exp_469;
    endcase
  end
  assign exp_470 = exp_470_reg;
  assign exp_469 = 0;

  reg [31:0] exp_464_reg;
  always@(*) begin
    case (exp_460)
      0:exp_464_reg <= exp_452;
      1:exp_464_reg <= exp_462;
      default:exp_464_reg <= exp_463;
    endcase
  end
  assign exp_464 = exp_464_reg;
  assign exp_460 = exp_435 == exp_459;
  assign exp_435 = exp_96[24:20];
  assign exp_459 = 0;
  assign exp_463 = 0;

  reg [31:0] exp_452_reg;
  always@(*) begin
    case (exp_432)
      0:exp_452_reg <= exp_428;
      1:exp_452_reg <= exp_433;
      default:exp_452_reg <= exp_451;
    endcase
  end
  assign exp_452 = exp_452_reg;
  assign exp_432 = exp_1008;
  assign exp_1008 = exp_1007 & exp_400;
  assign exp_1007 = exp_1006 & exp_408;
  assign exp_1006 = exp_1005 & exp_995;
  assign exp_1005 = exp_414 == exp_996;
  assign exp_414 = exp_96[24:20];
  assign exp_451 = 0;

  //Create RAM
  reg [31:0] exp_428_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_426) begin
      exp_428_ram[exp_422] <= exp_424;
    end
  end
  assign exp_428 = exp_428_ram[exp_423];
  assign exp_427 = exp_430;
  assign exp_430 = 1;
  assign exp_423 = exp_414;
  assign exp_426 = exp_1000;
  assign exp_1000 = exp_999 & exp_400;
  assign exp_999 = exp_995 & exp_408;
  assign exp_422 = exp_996;
  assign exp_424 = exp_994;
  assign exp_433 = exp_994;
  assign exp_462 = $signed(exp_461);
  assign exp_461 = 0;
  assign exp_468 = exp_465 + exp_467;
  assign exp_465 = 0;
  assign exp_467 = $signed(exp_466);
  assign exp_466 = exp_96[31:20];
  assign exp_484 = 0;

      reg [31:0] exp_412_reg = 0;
      always@(posedge clk) begin
        if (exp_411) begin
          exp_412_reg <= exp_410;
        end
      end
      assign exp_412 = exp_412_reg;
      assign exp_411 = exp_402 & exp_400;
  assign exp_558 = exp_522 - exp_523;
  assign exp_562 = exp_522 << exp_561;
  assign exp_561 = $signed(exp_556);
  assign exp_556 = exp_555 + exp_554;
  assign exp_555 = 0;
  assign exp_554 = exp_525;

      reg [4:0] exp_525_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_525_reg <= exp_474;
        end
      end
      assign exp_525 = exp_525_reg;
    
  reg [4:0] exp_474_reg;
  always@(*) begin
    case (exp_440)
      0:exp_474_reg <= exp_472;
      1:exp_474_reg <= exp_437;
      default:exp_474_reg <= exp_473;
    endcase
  end
  assign exp_474 = exp_474_reg;
  assign exp_473 = 0;
  assign exp_472 = exp_470[4:0];
  assign exp_437 = exp_96[24:20];
  assign exp_578 = $signed(exp_564);
  assign exp_564 = exp_563;
  assign exp_563 = $signed(exp_522) < $signed(exp_523);
  assign exp_579 = $signed(exp_570);
  assign exp_570 = exp_569;
  assign exp_569 = exp_566 < exp_568;
  assign exp_566 = exp_565 + exp_522;
  assign exp_565 = 0;
  assign exp_568 = exp_567 + exp_523;
  assign exp_567 = 0;
  assign exp_571 = exp_522 ^ exp_523;
  assign exp_575 = exp_574[31:0];
  assign exp_574 = $signed(exp_572) >>> $signed(exp_573);
  assign exp_572 = {exp_553, exp_522};
  reg [0:0] exp_553_reg;
  always@(*) begin
    case (exp_527)
      0:exp_553_reg <= exp_551;
      1:exp_553_reg <= exp_550;
      default:exp_553_reg <= exp_552;
    endcase
  end
  assign exp_553 = exp_553_reg;

      reg [0:0] exp_527_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_527_reg <= exp_471;
        end
      end
      assign exp_527 = exp_527_reg;
      assign exp_471 = exp_96[30:30];
  assign exp_552 = 0;
  assign exp_551 = 0;
  assign exp_550 = exp_522[31:31];
  assign exp_573 = $signed(exp_556);
  assign exp_576 = exp_522 | exp_523;
  assign exp_577 = exp_522 & exp_523;

  reg [31:0] exp_628_reg;
  always@(*) begin
    case (exp_531)
      0:exp_628_reg <= exp_618;
      1:exp_628_reg <= exp_621;
      2:exp_628_reg <= exp_394;
      3:exp_628_reg <= exp_622;
      4:exp_628_reg <= exp_623;
      5:exp_628_reg <= exp_624;
      6:exp_628_reg <= exp_625;
      7:exp_628_reg <= exp_626;
      default:exp_628_reg <= exp_627;
    endcase
  end
  assign exp_628 = exp_628_reg;
  assign exp_627 = 0;
  assign exp_618 = $signed(exp_617);
  assign exp_617 = exp_616 + exp_611;
  assign exp_616 = 0;

  reg [7:0] exp_611_reg;
  always@(*) begin
    case (exp_602)
      0:exp_611_reg <= exp_606;
      1:exp_611_reg <= exp_607;
      2:exp_611_reg <= exp_608;
      3:exp_611_reg <= exp_609;
      default:exp_611_reg <= exp_610;
    endcase
  end
  assign exp_611 = exp_611_reg;
  assign exp_602 = exp_601 + exp_600;
  assign exp_601 = 0;
  assign exp_600 = exp_599[1:0];
  assign exp_610 = 0;
  assign exp_606 = exp_394[7:0];
  assign exp_394 = exp_319;

  reg [31:0] exp_319_reg;
  always@(*) begin
    case (exp_316)
      0:exp_319_reg <= exp_296;
      1:exp_319_reg <= exp_307;
      default:exp_319_reg <= exp_318;
    endcase
  end
  assign exp_319 = exp_319_reg;
  assign exp_318 = 0;

  reg [31:0] exp_296_reg;
  always@(*) begin
    case (exp_293)
      0:exp_296_reg <= exp_194;
      1:exp_296_reg <= exp_284;
      default:exp_296_reg <= exp_295;
    endcase
  end
  assign exp_296 = exp_296_reg;
  assign exp_295 = 0;

  reg [31:0] exp_194_reg;
  always@(*) begin
    case (exp_191)
      0:exp_194_reg <= exp_153;
      1:exp_194_reg <= exp_182;
      default:exp_194_reg <= exp_193;
    endcase
  end
  assign exp_194 = exp_194_reg;
  assign exp_193 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 0;
    exp_54_ram[32] = 252;
    exp_54_ram[33] = 117;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 0;
    exp_54_ram[36] = 0;
    exp_54_ram[37] = 0;
    exp_54_ram[38] = 0;
    exp_54_ram[39] = 0;
    exp_54_ram[40] = 40;
    exp_54_ram[41] = 0;
    exp_54_ram[42] = 165;
    exp_54_ram[43] = 14;
    exp_54_ram[44] = 0;
    exp_54_ram[45] = 12;
    exp_54_ram[46] = 15;
    exp_54_ram[47] = 0;
    exp_54_ram[48] = 0;
    exp_54_ram[49] = 0;
    exp_54_ram[50] = 0;
    exp_54_ram[51] = 0;
    exp_54_ram[52] = 2;
    exp_54_ram[53] = 0;
    exp_54_ram[54] = 64;
    exp_54_ram[55] = 0;
    exp_54_ram[56] = 0;
    exp_54_ram[57] = 0;
    exp_54_ram[58] = 0;
    exp_54_ram[59] = 0;
    exp_54_ram[60] = 0;
    exp_54_ram[61] = 1;
    exp_54_ram[62] = 3;
    exp_54_ram[63] = 1;
    exp_54_ram[64] = 1;
    exp_54_ram[65] = 1;
    exp_54_ram[66] = 3;
    exp_54_ram[67] = 0;
    exp_54_ram[68] = 2;
    exp_54_ram[69] = 1;
    exp_54_ram[70] = 0;
    exp_54_ram[71] = 0;
    exp_54_ram[72] = 1;
    exp_54_ram[73] = 255;
    exp_54_ram[74] = 1;
    exp_54_ram[75] = 0;
    exp_54_ram[76] = 255;
    exp_54_ram[77] = 1;
    exp_54_ram[78] = 64;
    exp_54_ram[79] = 3;
    exp_54_ram[80] = 1;
    exp_54_ram[81] = 1;
    exp_54_ram[82] = 3;
    exp_54_ram[83] = 1;
    exp_54_ram[84] = 0;
    exp_54_ram[85] = 2;
    exp_54_ram[86] = 0;
    exp_54_ram[87] = 0;
    exp_54_ram[88] = 0;
    exp_54_ram[89] = 255;
    exp_54_ram[90] = 1;
    exp_54_ram[91] = 0;
    exp_54_ram[92] = 255;
    exp_54_ram[93] = 1;
    exp_54_ram[94] = 0;
    exp_54_ram[95] = 0;
    exp_54_ram[96] = 14;
    exp_54_ram[97] = 1;
    exp_54_ram[98] = 1;
    exp_54_ram[99] = 242;
    exp_54_ram[100] = 1;
    exp_54_ram[101] = 243;
    exp_54_ram[102] = 0;
    exp_54_ram[103] = 0;
    exp_54_ram[104] = 2;
    exp_54_ram[105] = 0;
    exp_54_ram[106] = 12;
    exp_54_ram[107] = 15;
    exp_54_ram[108] = 1;
    exp_54_ram[109] = 0;
    exp_54_ram[110] = 0;
    exp_54_ram[111] = 0;
    exp_54_ram[112] = 0;
    exp_54_ram[113] = 2;
    exp_54_ram[114] = 0;
    exp_54_ram[115] = 64;
    exp_54_ram[116] = 10;
    exp_54_ram[117] = 65;
    exp_54_ram[118] = 0;
    exp_54_ram[119] = 1;
    exp_54_ram[120] = 1;
    exp_54_ram[121] = 1;
    exp_54_ram[122] = 1;
    exp_54_ram[123] = 3;
    exp_54_ram[124] = 3;
    exp_54_ram[125] = 1;
    exp_54_ram[126] = 0;
    exp_54_ram[127] = 2;
    exp_54_ram[128] = 0;
    exp_54_ram[129] = 1;
    exp_54_ram[130] = 1;
    exp_54_ram[131] = 255;
    exp_54_ram[132] = 1;
    exp_54_ram[133] = 1;
    exp_54_ram[134] = 255;
    exp_54_ram[135] = 1;
    exp_54_ram[136] = 65;
    exp_54_ram[137] = 3;
    exp_54_ram[138] = 1;
    exp_54_ram[139] = 1;
    exp_54_ram[140] = 3;
    exp_54_ram[141] = 1;
    exp_54_ram[142] = 0;
    exp_54_ram[143] = 2;
    exp_54_ram[144] = 0;
    exp_54_ram[145] = 0;
    exp_54_ram[146] = 0;
    exp_54_ram[147] = 255;
    exp_54_ram[148] = 1;
    exp_54_ram[149] = 0;
    exp_54_ram[150] = 255;
    exp_54_ram[151] = 1;
    exp_54_ram[152] = 0;
    exp_54_ram[153] = 0;
    exp_54_ram[154] = 1;
    exp_54_ram[155] = 1;
    exp_54_ram[156] = 244;
    exp_54_ram[157] = 1;
    exp_54_ram[158] = 244;
    exp_54_ram[159] = 0;
    exp_54_ram[160] = 0;
    exp_54_ram[161] = 0;
    exp_54_ram[162] = 0;
    exp_54_ram[163] = 0;
    exp_54_ram[164] = 1;
    exp_54_ram[165] = 0;
    exp_54_ram[166] = 3;
    exp_54_ram[167] = 1;
    exp_54_ram[168] = 1;
    exp_54_ram[169] = 1;
    exp_54_ram[170] = 3;
    exp_54_ram[171] = 1;
    exp_54_ram[172] = 0;
    exp_54_ram[173] = 2;
    exp_54_ram[174] = 0;
    exp_54_ram[175] = 0;
    exp_54_ram[176] = 1;
    exp_54_ram[177] = 255;
    exp_54_ram[178] = 1;
    exp_54_ram[179] = 0;
    exp_54_ram[180] = 255;
    exp_54_ram[181] = 1;
    exp_54_ram[182] = 64;
    exp_54_ram[183] = 3;
    exp_54_ram[184] = 1;
    exp_54_ram[185] = 1;
    exp_54_ram[186] = 3;
    exp_54_ram[187] = 1;
    exp_54_ram[188] = 2;
    exp_54_ram[189] = 0;
    exp_54_ram[190] = 0;
    exp_54_ram[191] = 0;
    exp_54_ram[192] = 1;
    exp_54_ram[193] = 255;
    exp_54_ram[194] = 1;
    exp_54_ram[195] = 0;
    exp_54_ram[196] = 255;
    exp_54_ram[197] = 1;
    exp_54_ram[198] = 1;
    exp_54_ram[199] = 64;
    exp_54_ram[200] = 0;
    exp_54_ram[201] = 235;
    exp_54_ram[202] = 24;
    exp_54_ram[203] = 0;
    exp_54_ram[204] = 4;
    exp_54_ram[205] = 15;
    exp_54_ram[206] = 0;
    exp_54_ram[207] = 0;
    exp_54_ram[208] = 0;
    exp_54_ram[209] = 0;
    exp_54_ram[210] = 165;
    exp_54_ram[211] = 0;
    exp_54_ram[212] = 0;
    exp_54_ram[213] = 2;
    exp_54_ram[214] = 0;
    exp_54_ram[215] = 64;
    exp_54_ram[216] = 2;
    exp_54_ram[217] = 0;
    exp_54_ram[218] = 238;
    exp_54_ram[219] = 0;
    exp_54_ram[220] = 0;
    exp_54_ram[221] = 239;
    exp_54_ram[222] = 1;
    exp_54_ram[223] = 1;
    exp_54_ram[224] = 252;
    exp_54_ram[225] = 1;
    exp_54_ram[226] = 251;
    exp_54_ram[227] = 0;
    exp_54_ram[228] = 0;
    exp_54_ram[229] = 0;
    exp_54_ram[230] = 0;
    exp_54_ram[231] = 1;
    exp_54_ram[232] = 3;
    exp_54_ram[233] = 0;
    exp_54_ram[234] = 0;
    exp_54_ram[235] = 0;
    exp_54_ram[236] = 0;
    exp_54_ram[237] = 1;
    exp_54_ram[238] = 1;
    exp_54_ram[239] = 1;
    exp_54_ram[240] = 3;
    exp_54_ram[241] = 1;
    exp_54_ram[242] = 0;
    exp_54_ram[243] = 3;
    exp_54_ram[244] = 0;
    exp_54_ram[245] = 1;
    exp_54_ram[246] = 1;
    exp_54_ram[247] = 255;
    exp_54_ram[248] = 1;
    exp_54_ram[249] = 1;
    exp_54_ram[250] = 255;
    exp_54_ram[251] = 1;
    exp_54_ram[252] = 65;
    exp_54_ram[253] = 3;
    exp_54_ram[254] = 3;
    exp_54_ram[255] = 1;
    exp_54_ram[256] = 2;
    exp_54_ram[257] = 1;
    exp_54_ram[258] = 1;
    exp_54_ram[259] = 0;
    exp_54_ram[260] = 0;
    exp_54_ram[261] = 1;
    exp_54_ram[262] = 1;
    exp_54_ram[263] = 255;
    exp_54_ram[264] = 1;
    exp_54_ram[265] = 1;
    exp_54_ram[266] = 255;
    exp_54_ram[267] = 1;
    exp_54_ram[268] = 1;
    exp_54_ram[269] = 0;
    exp_54_ram[270] = 0;
    exp_54_ram[271] = 255;
    exp_54_ram[272] = 0;
    exp_54_ram[273] = 1;
    exp_54_ram[274] = 0;
    exp_54_ram[275] = 1;
    exp_54_ram[276] = 65;
    exp_54_ram[277] = 2;
    exp_54_ram[278] = 2;
    exp_54_ram[279] = 1;
    exp_54_ram[280] = 2;
    exp_54_ram[281] = 0;
    exp_54_ram[282] = 1;
    exp_54_ram[283] = 2;
    exp_54_ram[284] = 0;
    exp_54_ram[285] = 1;
    exp_54_ram[286] = 1;
    exp_54_ram[287] = 0;
    exp_54_ram[288] = 2;
    exp_54_ram[289] = 206;
    exp_54_ram[290] = 0;
    exp_54_ram[291] = 255;
    exp_54_ram[292] = 0;
    exp_54_ram[293] = 1;
    exp_54_ram[294] = 0;
    exp_54_ram[295] = 0;
    exp_54_ram[296] = 1;
    exp_54_ram[297] = 0;
    exp_54_ram[298] = 218;
    exp_54_ram[299] = 255;
    exp_54_ram[300] = 204;
    exp_54_ram[301] = 0;
    exp_54_ram[302] = 0;
    exp_54_ram[303] = 218;
    exp_54_ram[304] = 0;
    exp_54_ram[305] = 255;
    exp_54_ram[306] = 1;
    exp_54_ram[307] = 0;
    exp_54_ram[308] = 0;
    exp_54_ram[309] = 0;
    exp_54_ram[310] = 127;
    exp_54_ram[311] = 1;
    exp_54_ram[312] = 127;
    exp_54_ram[313] = 1;
    exp_54_ram[314] = 0;
    exp_54_ram[315] = 0;
    exp_54_ram[316] = 127;
    exp_54_ram[317] = 1;
    exp_54_ram[318] = 1;
    exp_54_ram[319] = 0;
    exp_54_ram[320] = 8;
    exp_54_ram[321] = 0;
    exp_54_ram[322] = 0;
    exp_54_ram[323] = 1;
    exp_54_ram[324] = 0;
    exp_54_ram[325] = 254;
    exp_54_ram[326] = 8;
    exp_54_ram[327] = 0;
    exp_54_ram[328] = 0;
    exp_54_ram[329] = 0;
    exp_54_ram[330] = 0;
    exp_54_ram[331] = 4;
    exp_54_ram[332] = 0;
    exp_54_ram[333] = 0;
    exp_54_ram[334] = 3;
    exp_54_ram[335] = 4;
    exp_54_ram[336] = 255;
    exp_54_ram[337] = 0;
    exp_54_ram[338] = 255;
    exp_54_ram[339] = 0;
    exp_54_ram[340] = 0;
    exp_54_ram[341] = 0;
    exp_54_ram[342] = 0;
    exp_54_ram[343] = 254;
    exp_54_ram[344] = 0;
    exp_54_ram[345] = 253;
    exp_54_ram[346] = 2;
    exp_54_ram[347] = 252;
    exp_54_ram[348] = 255;
    exp_54_ram[349] = 0;
    exp_54_ram[350] = 0;
    exp_54_ram[351] = 0;
    exp_54_ram[352] = 0;
    exp_54_ram[353] = 254;
    exp_54_ram[354] = 251;
    exp_54_ram[355] = 252;
    exp_54_ram[356] = 254;
    exp_54_ram[357] = 247;
    exp_54_ram[358] = 248;
    exp_54_ram[359] = 0;
    exp_54_ram[360] = 248;
    exp_54_ram[361] = 255;
    exp_54_ram[362] = 0;
    exp_54_ram[363] = 0;
    exp_54_ram[364] = 0;
    exp_54_ram[365] = 6;
    exp_54_ram[366] = 42;
    exp_54_ram[367] = 65;
    exp_54_ram[368] = 0;
    exp_54_ram[369] = 64;
    exp_54_ram[370] = 4;
    exp_54_ram[371] = 0;
    exp_54_ram[372] = 64;
    exp_54_ram[373] = 1;
    exp_54_ram[374] = 0;
    exp_54_ram[375] = 0;
    exp_54_ram[376] = 0;
    exp_54_ram[377] = 0;
    exp_54_ram[378] = 0;
    exp_54_ram[379] = 0;
    exp_54_ram[380] = 1;
    exp_54_ram[381] = 0;
    exp_54_ram[382] = 0;
    exp_54_ram[383] = 0;
    exp_54_ram[384] = 1;
    exp_54_ram[385] = 0;
    exp_54_ram[386] = 255;
    exp_54_ram[387] = 0;
    exp_54_ram[388] = 0;
    exp_54_ram[389] = 252;
    exp_54_ram[390] = 0;
    exp_54_ram[391] = 0;
    exp_54_ram[392] = 252;
    exp_54_ram[393] = 254;
    exp_54_ram[394] = 0;
    exp_54_ram[395] = 0;
    exp_54_ram[396] = 0;
    exp_54_ram[397] = 1;
    exp_54_ram[398] = 1;
    exp_54_ram[399] = 1;
    exp_54_ram[400] = 0;
    exp_54_ram[401] = 24;
    exp_54_ram[402] = 0;
    exp_54_ram[403] = 0;
    exp_54_ram[404] = 0;
    exp_54_ram[405] = 8;
    exp_54_ram[406] = 0;
    exp_54_ram[407] = 32;
    exp_54_ram[408] = 0;
    exp_54_ram[409] = 67;
    exp_54_ram[410] = 65;
    exp_54_ram[411] = 67;
    exp_54_ram[412] = 9;
    exp_54_ram[413] = 0;
    exp_54_ram[414] = 0;
    exp_54_ram[415] = 3;
    exp_54_ram[416] = 2;
    exp_54_ram[417] = 7;
    exp_54_ram[418] = 2;
    exp_54_ram[419] = 255;
    exp_54_ram[420] = 65;
    exp_54_ram[421] = 0;
    exp_54_ram[422] = 0;
    exp_54_ram[423] = 0;
    exp_54_ram[424] = 0;
    exp_54_ram[425] = 1;
    exp_54_ram[426] = 1;
    exp_54_ram[427] = 0;
    exp_54_ram[428] = 1;
    exp_54_ram[429] = 0;
    exp_54_ram[430] = 0;
    exp_54_ram[431] = 1;
    exp_54_ram[432] = 1;
    exp_54_ram[433] = 0;
    exp_54_ram[434] = 0;
    exp_54_ram[435] = 0;
    exp_54_ram[436] = 0;
    exp_54_ram[437] = 2;
    exp_54_ram[438] = 0;
    exp_54_ram[439] = 24;
    exp_54_ram[440] = 2;
    exp_54_ram[441] = 248;
    exp_54_ram[442] = 253;
    exp_54_ram[443] = 0;
    exp_54_ram[444] = 0;
    exp_54_ram[445] = 251;
    exp_54_ram[446] = 67;
    exp_54_ram[447] = 3;
    exp_54_ram[448] = 3;
    exp_54_ram[449] = 0;
    exp_54_ram[450] = 0;
    exp_54_ram[451] = 17;
    exp_54_ram[452] = 0;
    exp_54_ram[453] = 0;
    exp_54_ram[454] = 0;
    exp_54_ram[455] = 0;
    exp_54_ram[456] = 0;
    exp_54_ram[457] = 65;
    exp_54_ram[458] = 12;
    exp_54_ram[459] = 0;
    exp_54_ram[460] = 0;
    exp_54_ram[461] = 0;
    exp_54_ram[462] = 0;
    exp_54_ram[463] = 0;
    exp_54_ram[464] = 3;
    exp_54_ram[465] = 2;
    exp_54_ram[466] = 9;
    exp_54_ram[467] = 255;
    exp_54_ram[468] = 0;
    exp_54_ram[469] = 2;
    exp_54_ram[470] = 65;
    exp_54_ram[471] = 1;
    exp_54_ram[472] = 0;
    exp_54_ram[473] = 0;
    exp_54_ram[474] = 255;
    exp_54_ram[475] = 255;
    exp_54_ram[476] = 0;
    exp_54_ram[477] = 0;
    exp_54_ram[478] = 2;
    exp_54_ram[479] = 0;
    exp_54_ram[480] = 0;
    exp_54_ram[481] = 0;
    exp_54_ram[482] = 0;
    exp_54_ram[483] = 0;
    exp_54_ram[484] = 0;
    exp_54_ram[485] = 0;
    exp_54_ram[486] = 0;
    exp_54_ram[487] = 0;
    exp_54_ram[488] = 0;
    exp_54_ram[489] = 255;
    exp_54_ram[490] = 255;
    exp_54_ram[491] = 67;
    exp_54_ram[492] = 0;
    exp_54_ram[493] = 65;
    exp_54_ram[494] = 0;
    exp_54_ram[495] = 1;
    exp_54_ram[496] = 0;
    exp_54_ram[497] = 0;
    exp_54_ram[498] = 237;
    exp_54_ram[499] = 253;
    exp_54_ram[500] = 0;
    exp_54_ram[501] = 0;
    exp_54_ram[502] = 249;
    exp_54_ram[503] = 0;
    exp_54_ram[504] = 0;
    exp_54_ram[505] = 0;
    exp_54_ram[506] = 235;
    exp_54_ram[507] = 2;
    exp_54_ram[508] = 2;
    exp_54_ram[509] = 64;
    exp_54_ram[510] = 0;
    exp_54_ram[511] = 254;
    exp_54_ram[512] = 0;
    exp_54_ram[513] = 0;
    exp_54_ram[514] = 0;
    exp_54_ram[515] = 0;
    exp_54_ram[516] = 0;
    exp_54_ram[517] = 0;
    exp_54_ram[518] = 0;
    exp_54_ram[519] = 0;
    exp_54_ram[520] = 254;
    exp_54_ram[521] = 2;
    exp_54_ram[522] = 2;
    exp_54_ram[523] = 64;
    exp_54_ram[524] = 0;
    exp_54_ram[525] = 254;
    exp_54_ram[526] = 0;
    exp_54_ram[527] = 0;
    exp_54_ram[528] = 0;
    exp_54_ram[529] = 0;
    exp_54_ram[530] = 0;
    exp_54_ram[531] = 0;
    exp_54_ram[532] = 0;
    exp_54_ram[533] = 0;
    exp_54_ram[534] = 254;
    exp_54_ram[535] = 0;
    exp_54_ram[536] = 2;
    exp_54_ram[537] = 15;
    exp_54_ram[538] = 0;
    exp_54_ram[539] = 0;
    exp_54_ram[540] = 0;
    exp_54_ram[541] = 2;
    exp_54_ram[542] = 64;
    exp_54_ram[543] = 0;
    exp_54_ram[544] = 165;
    exp_54_ram[545] = 0;
    exp_54_ram[546] = 0;
    exp_54_ram[547] = 64;
    exp_54_ram[548] = 0;
    exp_54_ram[549] = 1;
    exp_54_ram[550] = 1;
    exp_54_ram[551] = 252;
    exp_54_ram[552] = 1;
    exp_54_ram[553] = 252;
    exp_54_ram[554] = 77;
    exp_54_ram[555] = 117;
    exp_54_ram[556] = 100;
    exp_54_ram[557] = 70;
    exp_54_ram[558] = 97;
    exp_54_ram[559] = 0;
    exp_54_ram[560] = 70;
    exp_54_ram[561] = 97;
    exp_54_ram[562] = 114;
    exp_54_ram[563] = 74;
    exp_54_ram[564] = 117;
    exp_54_ram[565] = 103;
    exp_54_ram[566] = 79;
    exp_54_ram[567] = 111;
    exp_54_ram[568] = 99;
    exp_54_ram[569] = 0;
    exp_54_ram[570] = 108;
    exp_54_ram[571] = 111;
    exp_54_ram[572] = 33;
    exp_54_ram[573] = 0;
    exp_54_ram[574] = 110;
    exp_54_ram[575] = 32;
    exp_54_ram[576] = 103;
    exp_54_ram[577] = 114;
    exp_54_ram[578] = 114;
    exp_54_ram[579] = 109;
    exp_54_ram[580] = 46;
    exp_54_ram[581] = 0;
    exp_54_ram[582] = 0;
    exp_54_ram[583] = 51;
    exp_54_ram[584] = 105;
    exp_54_ram[585] = 110;
    exp_54_ram[586] = 101;
    exp_54_ram[587] = 117;
    exp_54_ram[588] = 112;
    exp_54_ram[589] = 115;
    exp_54_ram[590] = 32;
    exp_54_ram[591] = 101;
    exp_54_ram[592] = 100;
    exp_54_ram[593] = 0;
    exp_54_ram[594] = 54;
    exp_54_ram[595] = 105;
    exp_54_ram[596] = 110;
    exp_54_ram[597] = 101;
    exp_54_ram[598] = 117;
    exp_54_ram[599] = 112;
    exp_54_ram[600] = 115;
    exp_54_ram[601] = 32;
    exp_54_ram[602] = 101;
    exp_54_ram[603] = 100;
    exp_54_ram[604] = 0;
    exp_54_ram[605] = 51;
    exp_54_ram[606] = 105;
    exp_54_ram[607] = 110;
    exp_54_ram[608] = 101;
    exp_54_ram[609] = 105;
    exp_54_ram[610] = 101;
    exp_54_ram[611] = 110;
    exp_54_ram[612] = 115;
    exp_54_ram[613] = 110;
    exp_54_ram[614] = 0;
    exp_54_ram[615] = 54;
    exp_54_ram[616] = 105;
    exp_54_ram[617] = 110;
    exp_54_ram[618] = 101;
    exp_54_ram[619] = 105;
    exp_54_ram[620] = 101;
    exp_54_ram[621] = 110;
    exp_54_ram[622] = 115;
    exp_54_ram[623] = 110;
    exp_54_ram[624] = 0;
    exp_54_ram[625] = 114;
    exp_54_ram[626] = 0;
    exp_54_ram[627] = 116;
    exp_54_ram[628] = 0;
    exp_54_ram[629] = 58;
    exp_54_ram[630] = 0;
    exp_54_ram[631] = 114;
    exp_54_ram[632] = 0;
    exp_54_ram[633] = 117;
    exp_54_ram[634] = 10;
    exp_54_ram[635] = 0;
    exp_54_ram[636] = 105;
    exp_54_ram[637] = 86;
    exp_54_ram[638] = 109;
    exp_54_ram[639] = 0;
    exp_54_ram[640] = 32;
    exp_54_ram[641] = 108;
    exp_54_ram[642] = 111;
    exp_54_ram[643] = 10;
    exp_54_ram[644] = 0;
    exp_54_ram[645] = 75;
    exp_54_ram[646] = 104;
    exp_54_ram[647] = 105;
    exp_54_ram[648] = 10;
    exp_54_ram[649] = 0;
    exp_54_ram[650] = 84;
    exp_54_ram[651] = 32;
    exp_54_ram[652] = 116;
    exp_54_ram[653] = 105;
    exp_54_ram[654] = 105;
    exp_54_ram[655] = 0;
    exp_54_ram[656] = 87;
    exp_54_ram[657] = 32;
    exp_54_ram[658] = 99;
    exp_54_ram[659] = 0;
    exp_54_ram[660] = 2;
    exp_54_ram[661] = 3;
    exp_54_ram[662] = 4;
    exp_54_ram[663] = 4;
    exp_54_ram[664] = 5;
    exp_54_ram[665] = 5;
    exp_54_ram[666] = 5;
    exp_54_ram[667] = 5;
    exp_54_ram[668] = 6;
    exp_54_ram[669] = 6;
    exp_54_ram[670] = 6;
    exp_54_ram[671] = 6;
    exp_54_ram[672] = 6;
    exp_54_ram[673] = 6;
    exp_54_ram[674] = 6;
    exp_54_ram[675] = 6;
    exp_54_ram[676] = 7;
    exp_54_ram[677] = 7;
    exp_54_ram[678] = 7;
    exp_54_ram[679] = 7;
    exp_54_ram[680] = 7;
    exp_54_ram[681] = 7;
    exp_54_ram[682] = 7;
    exp_54_ram[683] = 7;
    exp_54_ram[684] = 7;
    exp_54_ram[685] = 7;
    exp_54_ram[686] = 7;
    exp_54_ram[687] = 7;
    exp_54_ram[688] = 7;
    exp_54_ram[689] = 7;
    exp_54_ram[690] = 7;
    exp_54_ram[691] = 7;
    exp_54_ram[692] = 8;
    exp_54_ram[693] = 8;
    exp_54_ram[694] = 8;
    exp_54_ram[695] = 8;
    exp_54_ram[696] = 8;
    exp_54_ram[697] = 8;
    exp_54_ram[698] = 8;
    exp_54_ram[699] = 8;
    exp_54_ram[700] = 8;
    exp_54_ram[701] = 8;
    exp_54_ram[702] = 8;
    exp_54_ram[703] = 8;
    exp_54_ram[704] = 8;
    exp_54_ram[705] = 8;
    exp_54_ram[706] = 8;
    exp_54_ram[707] = 8;
    exp_54_ram[708] = 8;
    exp_54_ram[709] = 8;
    exp_54_ram[710] = 8;
    exp_54_ram[711] = 8;
    exp_54_ram[712] = 8;
    exp_54_ram[713] = 8;
    exp_54_ram[714] = 8;
    exp_54_ram[715] = 8;
    exp_54_ram[716] = 8;
    exp_54_ram[717] = 8;
    exp_54_ram[718] = 8;
    exp_54_ram[719] = 8;
    exp_54_ram[720] = 8;
    exp_54_ram[721] = 8;
    exp_54_ram[722] = 8;
    exp_54_ram[723] = 8;
    exp_54_ram[724] = 253;
    exp_54_ram[725] = 2;
    exp_54_ram[726] = 3;
    exp_54_ram[727] = 252;
    exp_54_ram[728] = 253;
    exp_54_ram[729] = 254;
    exp_54_ram[730] = 254;
    exp_54_ram[731] = 0;
    exp_54_ram[732] = 0;
    exp_54_ram[733] = 2;
    exp_54_ram[734] = 3;
    exp_54_ram[735] = 0;
    exp_54_ram[736] = 253;
    exp_54_ram[737] = 2;
    exp_54_ram[738] = 3;
    exp_54_ram[739] = 252;
    exp_54_ram[740] = 252;
    exp_54_ram[741] = 253;
    exp_54_ram[742] = 254;
    exp_54_ram[743] = 253;
    exp_54_ram[744] = 254;
    exp_54_ram[745] = 0;
    exp_54_ram[746] = 253;
    exp_54_ram[747] = 0;
    exp_54_ram[748] = 2;
    exp_54_ram[749] = 3;
    exp_54_ram[750] = 0;
    exp_54_ram[751] = 255;
    exp_54_ram[752] = 0;
    exp_54_ram[753] = 0;
    exp_54_ram[754] = 1;
    exp_54_ram[755] = 0;
    exp_54_ram[756] = 13;
    exp_54_ram[757] = 0;
    exp_54_ram[758] = 247;
    exp_54_ram[759] = 0;
    exp_54_ram[760] = 0;
    exp_54_ram[761] = 0;
    exp_54_ram[762] = 0;
    exp_54_ram[763] = 1;
    exp_54_ram[764] = 0;
    exp_54_ram[765] = 253;
    exp_54_ram[766] = 2;
    exp_54_ram[767] = 2;
    exp_54_ram[768] = 3;
    exp_54_ram[769] = 252;
    exp_54_ram[770] = 252;
    exp_54_ram[771] = 254;
    exp_54_ram[772] = 2;
    exp_54_ram[773] = 254;
    exp_54_ram[774] = 0;
    exp_54_ram[775] = 254;
    exp_54_ram[776] = 253;
    exp_54_ram[777] = 0;
    exp_54_ram[778] = 0;
    exp_54_ram[779] = 253;
    exp_54_ram[780] = 0;
    exp_54_ram[781] = 244;
    exp_54_ram[782] = 253;
    exp_54_ram[783] = 254;
    exp_54_ram[784] = 0;
    exp_54_ram[785] = 0;
    exp_54_ram[786] = 252;
    exp_54_ram[787] = 254;
    exp_54_ram[788] = 0;
    exp_54_ram[789] = 2;
    exp_54_ram[790] = 2;
    exp_54_ram[791] = 3;
    exp_54_ram[792] = 0;
    exp_54_ram[793] = 254;
    exp_54_ram[794] = 0;
    exp_54_ram[795] = 0;
    exp_54_ram[796] = 2;
    exp_54_ram[797] = 254;
    exp_54_ram[798] = 0;
    exp_54_ram[799] = 13;
    exp_54_ram[800] = 0;
    exp_54_ram[801] = 254;
    exp_54_ram[802] = 246;
    exp_54_ram[803] = 0;
    exp_54_ram[804] = 13;
    exp_54_ram[805] = 0;
    exp_54_ram[806] = 0;
    exp_54_ram[807] = 238;
    exp_54_ram[808] = 0;
    exp_54_ram[809] = 0;
    exp_54_ram[810] = 1;
    exp_54_ram[811] = 1;
    exp_54_ram[812] = 2;
    exp_54_ram[813] = 0;
    exp_54_ram[814] = 254;
    exp_54_ram[815] = 0;
    exp_54_ram[816] = 2;
    exp_54_ram[817] = 0;
    exp_54_ram[818] = 254;
    exp_54_ram[819] = 254;
    exp_54_ram[820] = 254;
    exp_54_ram[821] = 254;
    exp_54_ram[822] = 0;
    exp_54_ram[823] = 1;
    exp_54_ram[824] = 2;
    exp_54_ram[825] = 0;
    exp_54_ram[826] = 254;
    exp_54_ram[827] = 0;
    exp_54_ram[828] = 0;
    exp_54_ram[829] = 2;
    exp_54_ram[830] = 0;
    exp_54_ram[831] = 254;
    exp_54_ram[832] = 254;
    exp_54_ram[833] = 254;
    exp_54_ram[834] = 254;
    exp_54_ram[835] = 254;
    exp_54_ram[836] = 0;
    exp_54_ram[837] = 254;
    exp_54_ram[838] = 0;
    exp_54_ram[839] = 31;
    exp_54_ram[840] = 0;
    exp_54_ram[841] = 1;
    exp_54_ram[842] = 1;
    exp_54_ram[843] = 2;
    exp_54_ram[844] = 0;
    exp_54_ram[845] = 253;
    exp_54_ram[846] = 2;
    exp_54_ram[847] = 3;
    exp_54_ram[848] = 252;
    exp_54_ram[849] = 252;
    exp_54_ram[850] = 253;
    exp_54_ram[851] = 254;
    exp_54_ram[852] = 1;
    exp_54_ram[853] = 254;
    exp_54_ram[854] = 0;
    exp_54_ram[855] = 254;
    exp_54_ram[856] = 254;
    exp_54_ram[857] = 0;
    exp_54_ram[858] = 0;
    exp_54_ram[859] = 253;
    exp_54_ram[860] = 255;
    exp_54_ram[861] = 252;
    exp_54_ram[862] = 252;
    exp_54_ram[863] = 254;
    exp_54_ram[864] = 253;
    exp_54_ram[865] = 64;
    exp_54_ram[866] = 0;
    exp_54_ram[867] = 2;
    exp_54_ram[868] = 3;
    exp_54_ram[869] = 0;
    exp_54_ram[870] = 254;
    exp_54_ram[871] = 0;
    exp_54_ram[872] = 2;
    exp_54_ram[873] = 0;
    exp_54_ram[874] = 254;
    exp_54_ram[875] = 254;
    exp_54_ram[876] = 2;
    exp_54_ram[877] = 0;
    exp_54_ram[878] = 254;
    exp_54_ram[879] = 3;
    exp_54_ram[880] = 0;
    exp_54_ram[881] = 0;
    exp_54_ram[882] = 0;
    exp_54_ram[883] = 0;
    exp_54_ram[884] = 0;
    exp_54_ram[885] = 15;
    exp_54_ram[886] = 0;
    exp_54_ram[887] = 1;
    exp_54_ram[888] = 2;
    exp_54_ram[889] = 0;
    exp_54_ram[890] = 253;
    exp_54_ram[891] = 2;
    exp_54_ram[892] = 2;
    exp_54_ram[893] = 3;
    exp_54_ram[894] = 252;
    exp_54_ram[895] = 254;
    exp_54_ram[896] = 4;
    exp_54_ram[897] = 254;
    exp_54_ram[898] = 0;
    exp_54_ram[899] = 0;
    exp_54_ram[900] = 0;
    exp_54_ram[901] = 0;
    exp_54_ram[902] = 0;
    exp_54_ram[903] = 253;
    exp_54_ram[904] = 0;
    exp_54_ram[905] = 0;
    exp_54_ram[906] = 253;
    exp_54_ram[907] = 0;
    exp_54_ram[908] = 0;
    exp_54_ram[909] = 0;
    exp_54_ram[910] = 253;
    exp_54_ram[911] = 254;
    exp_54_ram[912] = 253;
    exp_54_ram[913] = 0;
    exp_54_ram[914] = 0;
    exp_54_ram[915] = 0;
    exp_54_ram[916] = 244;
    exp_54_ram[917] = 0;
    exp_54_ram[918] = 250;
    exp_54_ram[919] = 254;
    exp_54_ram[920] = 0;
    exp_54_ram[921] = 2;
    exp_54_ram[922] = 2;
    exp_54_ram[923] = 3;
    exp_54_ram[924] = 0;
    exp_54_ram[925] = 252;
    exp_54_ram[926] = 2;
    exp_54_ram[927] = 2;
    exp_54_ram[928] = 4;
    exp_54_ram[929] = 252;
    exp_54_ram[930] = 252;
    exp_54_ram[931] = 252;
    exp_54_ram[932] = 252;
    exp_54_ram[933] = 252;
    exp_54_ram[934] = 252;
    exp_54_ram[935] = 253;
    exp_54_ram[936] = 253;
    exp_54_ram[937] = 253;
    exp_54_ram[938] = 254;
    exp_54_ram[939] = 252;
    exp_54_ram[940] = 0;
    exp_54_ram[941] = 8;
    exp_54_ram[942] = 252;
    exp_54_ram[943] = 0;
    exp_54_ram[944] = 8;
    exp_54_ram[945] = 252;
    exp_54_ram[946] = 254;
    exp_54_ram[947] = 3;
    exp_54_ram[948] = 253;
    exp_54_ram[949] = 0;
    exp_54_ram[950] = 252;
    exp_54_ram[951] = 253;
    exp_54_ram[952] = 253;
    exp_54_ram[953] = 0;
    exp_54_ram[954] = 253;
    exp_54_ram[955] = 2;
    exp_54_ram[956] = 0;
    exp_54_ram[957] = 254;
    exp_54_ram[958] = 0;
    exp_54_ram[959] = 254;
    exp_54_ram[960] = 254;
    exp_54_ram[961] = 252;
    exp_54_ram[962] = 252;
    exp_54_ram[963] = 4;
    exp_54_ram[964] = 252;
    exp_54_ram[965] = 255;
    exp_54_ram[966] = 252;
    exp_54_ram[967] = 252;
    exp_54_ram[968] = 252;
    exp_54_ram[969] = 0;
    exp_54_ram[970] = 0;
    exp_54_ram[971] = 253;
    exp_54_ram[972] = 0;
    exp_54_ram[973] = 252;
    exp_54_ram[974] = 253;
    exp_54_ram[975] = 253;
    exp_54_ram[976] = 0;
    exp_54_ram[977] = 253;
    exp_54_ram[978] = 0;
    exp_54_ram[979] = 252;
    exp_54_ram[980] = 252;
    exp_54_ram[981] = 252;
    exp_54_ram[982] = 0;
    exp_54_ram[983] = 4;
    exp_54_ram[984] = 2;
    exp_54_ram[985] = 253;
    exp_54_ram[986] = 0;
    exp_54_ram[987] = 252;
    exp_54_ram[988] = 253;
    exp_54_ram[989] = 253;
    exp_54_ram[990] = 0;
    exp_54_ram[991] = 253;
    exp_54_ram[992] = 2;
    exp_54_ram[993] = 0;
    exp_54_ram[994] = 253;
    exp_54_ram[995] = 254;
    exp_54_ram[996] = 64;
    exp_54_ram[997] = 252;
    exp_54_ram[998] = 252;
    exp_54_ram[999] = 253;
    exp_54_ram[1000] = 0;
    exp_54_ram[1001] = 3;
    exp_54_ram[1002] = 3;
    exp_54_ram[1003] = 4;
    exp_54_ram[1004] = 0;
    exp_54_ram[1005] = 253;
    exp_54_ram[1006] = 2;
    exp_54_ram[1007] = 2;
    exp_54_ram[1008] = 3;
    exp_54_ram[1009] = 254;
    exp_54_ram[1010] = 254;
    exp_54_ram[1011] = 254;
    exp_54_ram[1012] = 254;
    exp_54_ram[1013] = 252;
    exp_54_ram[1014] = 252;
    exp_54_ram[1015] = 0;
    exp_54_ram[1016] = 253;
    exp_54_ram[1017] = 252;
    exp_54_ram[1018] = 0;
    exp_54_ram[1019] = 0;
    exp_54_ram[1020] = 10;
    exp_54_ram[1021] = 0;
    exp_54_ram[1022] = 4;
    exp_54_ram[1023] = 0;
    exp_54_ram[1024] = 0;
    exp_54_ram[1025] = 4;
    exp_54_ram[1026] = 253;
    exp_54_ram[1027] = 0;
    exp_54_ram[1028] = 0;
    exp_54_ram[1029] = 0;
    exp_54_ram[1030] = 2;
    exp_54_ram[1031] = 0;
    exp_54_ram[1032] = 255;
    exp_54_ram[1033] = 0;
    exp_54_ram[1034] = 2;
    exp_54_ram[1035] = 253;
    exp_54_ram[1036] = 0;
    exp_54_ram[1037] = 252;
    exp_54_ram[1038] = 253;
    exp_54_ram[1039] = 0;
    exp_54_ram[1040] = 3;
    exp_54_ram[1041] = 0;
    exp_54_ram[1042] = 253;
    exp_54_ram[1043] = 0;
    exp_54_ram[1044] = 2;
    exp_54_ram[1045] = 253;
    exp_54_ram[1046] = 1;
    exp_54_ram[1047] = 252;
    exp_54_ram[1048] = 2;
    exp_54_ram[1049] = 253;
    exp_54_ram[1050] = 0;
    exp_54_ram[1051] = 252;
    exp_54_ram[1052] = 253;
    exp_54_ram[1053] = 0;
    exp_54_ram[1054] = 3;
    exp_54_ram[1055] = 0;
    exp_54_ram[1056] = 0;
    exp_54_ram[1057] = 0;
    exp_54_ram[1058] = 0;
    exp_54_ram[1059] = 253;
    exp_54_ram[1060] = 0;
    exp_54_ram[1061] = 0;
    exp_54_ram[1062] = 253;
    exp_54_ram[1063] = 1;
    exp_54_ram[1064] = 252;
    exp_54_ram[1065] = 0;
    exp_54_ram[1066] = 1;
    exp_54_ram[1067] = 20;
    exp_54_ram[1068] = 0;
    exp_54_ram[1069] = 64;
    exp_54_ram[1070] = 4;
    exp_54_ram[1071] = 253;
    exp_54_ram[1072] = 4;
    exp_54_ram[1073] = 253;
    exp_54_ram[1074] = 0;
    exp_54_ram[1075] = 0;
    exp_54_ram[1076] = 253;
    exp_54_ram[1077] = 0;
    exp_54_ram[1078] = 2;
    exp_54_ram[1079] = 253;
    exp_54_ram[1080] = 255;
    exp_54_ram[1081] = 252;
    exp_54_ram[1082] = 253;
    exp_54_ram[1083] = 0;
    exp_54_ram[1084] = 253;
    exp_54_ram[1085] = 1;
    exp_54_ram[1086] = 0;
    exp_54_ram[1087] = 253;
    exp_54_ram[1088] = 255;
    exp_54_ram[1089] = 252;
    exp_54_ram[1090] = 253;
    exp_54_ram[1091] = 1;
    exp_54_ram[1092] = 2;
    exp_54_ram[1093] = 0;
    exp_54_ram[1094] = 2;
    exp_54_ram[1095] = 2;
    exp_54_ram[1096] = 253;
    exp_54_ram[1097] = 1;
    exp_54_ram[1098] = 2;
    exp_54_ram[1099] = 253;
    exp_54_ram[1100] = 0;
    exp_54_ram[1101] = 252;
    exp_54_ram[1102] = 253;
    exp_54_ram[1103] = 0;
    exp_54_ram[1104] = 7;
    exp_54_ram[1105] = 0;
    exp_54_ram[1106] = 7;
    exp_54_ram[1107] = 253;
    exp_54_ram[1108] = 1;
    exp_54_ram[1109] = 2;
    exp_54_ram[1110] = 0;
    exp_54_ram[1111] = 2;
    exp_54_ram[1112] = 2;
    exp_54_ram[1113] = 253;
    exp_54_ram[1114] = 1;
    exp_54_ram[1115] = 2;
    exp_54_ram[1116] = 253;
    exp_54_ram[1117] = 0;
    exp_54_ram[1118] = 252;
    exp_54_ram[1119] = 253;
    exp_54_ram[1120] = 0;
    exp_54_ram[1121] = 5;
    exp_54_ram[1122] = 0;
    exp_54_ram[1123] = 3;
    exp_54_ram[1124] = 253;
    exp_54_ram[1125] = 0;
    exp_54_ram[1126] = 2;
    exp_54_ram[1127] = 253;
    exp_54_ram[1128] = 1;
    exp_54_ram[1129] = 2;
    exp_54_ram[1130] = 253;
    exp_54_ram[1131] = 0;
    exp_54_ram[1132] = 252;
    exp_54_ram[1133] = 253;
    exp_54_ram[1134] = 0;
    exp_54_ram[1135] = 6;
    exp_54_ram[1136] = 0;
    exp_54_ram[1137] = 253;
    exp_54_ram[1138] = 1;
    exp_54_ram[1139] = 2;
    exp_54_ram[1140] = 253;
    exp_54_ram[1141] = 0;
    exp_54_ram[1142] = 252;
    exp_54_ram[1143] = 253;
    exp_54_ram[1144] = 0;
    exp_54_ram[1145] = 3;
    exp_54_ram[1146] = 0;
    exp_54_ram[1147] = 253;
    exp_54_ram[1148] = 1;
    exp_54_ram[1149] = 8;
    exp_54_ram[1150] = 253;
    exp_54_ram[1151] = 2;
    exp_54_ram[1152] = 253;
    exp_54_ram[1153] = 0;
    exp_54_ram[1154] = 252;
    exp_54_ram[1155] = 253;
    exp_54_ram[1156] = 0;
    exp_54_ram[1157] = 2;
    exp_54_ram[1158] = 0;
    exp_54_ram[1159] = 5;
    exp_54_ram[1160] = 0;
    exp_54_ram[1161] = 0;
    exp_54_ram[1162] = 2;
    exp_54_ram[1163] = 253;
    exp_54_ram[1164] = 0;
    exp_54_ram[1165] = 252;
    exp_54_ram[1166] = 253;
    exp_54_ram[1167] = 0;
    exp_54_ram[1168] = 2;
    exp_54_ram[1169] = 0;
    exp_54_ram[1170] = 2;
    exp_54_ram[1171] = 0;
    exp_54_ram[1172] = 0;
    exp_54_ram[1173] = 2;
    exp_54_ram[1174] = 253;
    exp_54_ram[1175] = 0;
    exp_54_ram[1176] = 252;
    exp_54_ram[1177] = 253;
    exp_54_ram[1178] = 0;
    exp_54_ram[1179] = 2;
    exp_54_ram[1180] = 0;
    exp_54_ram[1181] = 0;
    exp_54_ram[1182] = 0;
    exp_54_ram[1183] = 253;
    exp_54_ram[1184] = 253;
    exp_54_ram[1185] = 254;
    exp_54_ram[1186] = 254;
    exp_54_ram[1187] = 254;
    exp_54_ram[1188] = 254;
    exp_54_ram[1189] = 190;
    exp_54_ram[1190] = 0;
    exp_54_ram[1191] = 0;
    exp_54_ram[1192] = 2;
    exp_54_ram[1193] = 2;
    exp_54_ram[1194] = 3;
    exp_54_ram[1195] = 0;
    exp_54_ram[1196] = 249;
    exp_54_ram[1197] = 6;
    exp_54_ram[1198] = 6;
    exp_54_ram[1199] = 7;
    exp_54_ram[1200] = 250;
    exp_54_ram[1201] = 250;
    exp_54_ram[1202] = 250;
    exp_54_ram[1203] = 250;
    exp_54_ram[1204] = 250;
    exp_54_ram[1205] = 251;
    exp_54_ram[1206] = 251;
    exp_54_ram[1207] = 250;
    exp_54_ram[1208] = 254;
    exp_54_ram[1209] = 250;
    exp_54_ram[1210] = 0;
    exp_54_ram[1211] = 0;
    exp_54_ram[1212] = 254;
    exp_54_ram[1213] = 0;
    exp_54_ram[1214] = 0;
    exp_54_ram[1215] = 64;
    exp_54_ram[1216] = 0;
    exp_54_ram[1217] = 250;
    exp_54_ram[1218] = 8;
    exp_54_ram[1219] = 250;
    exp_54_ram[1220] = 250;
    exp_54_ram[1221] = 2;
    exp_54_ram[1222] = 254;
    exp_54_ram[1223] = 254;
    exp_54_ram[1224] = 0;
    exp_54_ram[1225] = 0;
    exp_54_ram[1226] = 254;
    exp_54_ram[1227] = 3;
    exp_54_ram[1228] = 15;
    exp_54_ram[1229] = 3;
    exp_54_ram[1230] = 0;
    exp_54_ram[1231] = 2;
    exp_54_ram[1232] = 0;
    exp_54_ram[1233] = 4;
    exp_54_ram[1234] = 0;
    exp_54_ram[1235] = 6;
    exp_54_ram[1236] = 254;
    exp_54_ram[1237] = 0;
    exp_54_ram[1238] = 15;
    exp_54_ram[1239] = 255;
    exp_54_ram[1240] = 15;
    exp_54_ram[1241] = 254;
    exp_54_ram[1242] = 0;
    exp_54_ram[1243] = 254;
    exp_54_ram[1244] = 255;
    exp_54_ram[1245] = 0;
    exp_54_ram[1246] = 252;
    exp_54_ram[1247] = 250;
    exp_54_ram[1248] = 250;
    exp_54_ram[1249] = 2;
    exp_54_ram[1250] = 250;
    exp_54_ram[1251] = 250;
    exp_54_ram[1252] = 0;
    exp_54_ram[1253] = 254;
    exp_54_ram[1254] = 1;
    exp_54_ram[1255] = 246;
    exp_54_ram[1256] = 250;
    exp_54_ram[1257] = 252;
    exp_54_ram[1258] = 0;
    exp_54_ram[1259] = 0;
    exp_54_ram[1260] = 0;
    exp_54_ram[1261] = 0;
    exp_54_ram[1262] = 250;
    exp_54_ram[1263] = 0;
    exp_54_ram[1264] = 250;
    exp_54_ram[1265] = 0;
    exp_54_ram[1266] = 254;
    exp_54_ram[1267] = 251;
    exp_54_ram[1268] = 251;
    exp_54_ram[1269] = 251;
    exp_54_ram[1270] = 251;
    exp_54_ram[1271] = 189;
    exp_54_ram[1272] = 0;
    exp_54_ram[1273] = 0;
    exp_54_ram[1274] = 6;
    exp_54_ram[1275] = 6;
    exp_54_ram[1276] = 7;
    exp_54_ram[1277] = 0;
    exp_54_ram[1278] = 248;
    exp_54_ram[1279] = 6;
    exp_54_ram[1280] = 6;
    exp_54_ram[1281] = 8;
    exp_54_ram[1282] = 250;
    exp_54_ram[1283] = 250;
    exp_54_ram[1284] = 250;
    exp_54_ram[1285] = 250;
    exp_54_ram[1286] = 248;
    exp_54_ram[1287] = 252;
    exp_54_ram[1288] = 250;
    exp_54_ram[1289] = 32;
    exp_54_ram[1290] = 0;
    exp_54_ram[1291] = 203;
    exp_54_ram[1292] = 250;
    exp_54_ram[1293] = 32;
    exp_54_ram[1294] = 250;
    exp_54_ram[1295] = 0;
    exp_54_ram[1296] = 2;
    exp_54_ram[1297] = 2;
    exp_54_ram[1298] = 250;
    exp_54_ram[1299] = 0;
    exp_54_ram[1300] = 253;
    exp_54_ram[1301] = 0;
    exp_54_ram[1302] = 252;
    exp_54_ram[1303] = 250;
    exp_54_ram[1304] = 250;
    exp_54_ram[1305] = 0;
    exp_54_ram[1306] = 250;
    exp_54_ram[1307] = 0;
    exp_54_ram[1308] = 250;
    exp_54_ram[1309] = 0;
    exp_54_ram[1310] = 250;
    exp_54_ram[1311] = 28;
    exp_54_ram[1312] = 250;
    exp_54_ram[1313] = 0;
    exp_54_ram[1314] = 250;
    exp_54_ram[1315] = 254;
    exp_54_ram[1316] = 250;
    exp_54_ram[1317] = 0;
    exp_54_ram[1318] = 254;
    exp_54_ram[1319] = 1;
    exp_54_ram[1320] = 12;
    exp_54_ram[1321] = 0;
    exp_54_ram[1322] = 0;
    exp_54_ram[1323] = 14;
    exp_54_ram[1324] = 0;
    exp_54_ram[1325] = 0;
    exp_54_ram[1326] = 0;
    exp_54_ram[1327] = 254;
    exp_54_ram[1328] = 0;
    exp_54_ram[1329] = 254;
    exp_54_ram[1330] = 250;
    exp_54_ram[1331] = 0;
    exp_54_ram[1332] = 250;
    exp_54_ram[1333] = 0;
    exp_54_ram[1334] = 254;
    exp_54_ram[1335] = 9;
    exp_54_ram[1336] = 254;
    exp_54_ram[1337] = 0;
    exp_54_ram[1338] = 254;
    exp_54_ram[1339] = 250;
    exp_54_ram[1340] = 0;
    exp_54_ram[1341] = 250;
    exp_54_ram[1342] = 0;
    exp_54_ram[1343] = 254;
    exp_54_ram[1344] = 7;
    exp_54_ram[1345] = 254;
    exp_54_ram[1346] = 0;
    exp_54_ram[1347] = 254;
    exp_54_ram[1348] = 250;
    exp_54_ram[1349] = 0;
    exp_54_ram[1350] = 250;
    exp_54_ram[1351] = 0;
    exp_54_ram[1352] = 254;
    exp_54_ram[1353] = 5;
    exp_54_ram[1354] = 254;
    exp_54_ram[1355] = 0;
    exp_54_ram[1356] = 254;
    exp_54_ram[1357] = 250;
    exp_54_ram[1358] = 0;
    exp_54_ram[1359] = 250;
    exp_54_ram[1360] = 0;
    exp_54_ram[1361] = 254;
    exp_54_ram[1362] = 3;
    exp_54_ram[1363] = 254;
    exp_54_ram[1364] = 1;
    exp_54_ram[1365] = 254;
    exp_54_ram[1366] = 250;
    exp_54_ram[1367] = 0;
    exp_54_ram[1368] = 250;
    exp_54_ram[1369] = 0;
    exp_54_ram[1370] = 254;
    exp_54_ram[1371] = 0;
    exp_54_ram[1372] = 254;
    exp_54_ram[1373] = 0;
    exp_54_ram[1374] = 254;
    exp_54_ram[1375] = 240;
    exp_54_ram[1376] = 254;
    exp_54_ram[1377] = 250;
    exp_54_ram[1378] = 0;
    exp_54_ram[1379] = 0;
    exp_54_ram[1380] = 128;
    exp_54_ram[1381] = 0;
    exp_54_ram[1382] = 0;
    exp_54_ram[1383] = 250;
    exp_54_ram[1384] = 0;
    exp_54_ram[1385] = 132;
    exp_54_ram[1386] = 254;
    exp_54_ram[1387] = 6;
    exp_54_ram[1388] = 250;
    exp_54_ram[1389] = 0;
    exp_54_ram[1390] = 2;
    exp_54_ram[1391] = 4;
    exp_54_ram[1392] = 249;
    exp_54_ram[1393] = 0;
    exp_54_ram[1394] = 248;
    exp_54_ram[1395] = 0;
    exp_54_ram[1396] = 252;
    exp_54_ram[1397] = 252;
    exp_54_ram[1398] = 2;
    exp_54_ram[1399] = 254;
    exp_54_ram[1400] = 0;
    exp_54_ram[1401] = 254;
    exp_54_ram[1402] = 252;
    exp_54_ram[1403] = 64;
    exp_54_ram[1404] = 254;
    exp_54_ram[1405] = 0;
    exp_54_ram[1406] = 252;
    exp_54_ram[1407] = 254;
    exp_54_ram[1408] = 250;
    exp_54_ram[1409] = 0;
    exp_54_ram[1410] = 250;
    exp_54_ram[1411] = 254;
    exp_54_ram[1412] = 250;
    exp_54_ram[1413] = 0;
    exp_54_ram[1414] = 2;
    exp_54_ram[1415] = 8;
    exp_54_ram[1416] = 254;
    exp_54_ram[1417] = 64;
    exp_54_ram[1418] = 254;
    exp_54_ram[1419] = 250;
    exp_54_ram[1420] = 0;
    exp_54_ram[1421] = 250;
    exp_54_ram[1422] = 250;
    exp_54_ram[1423] = 0;
    exp_54_ram[1424] = 0;
    exp_54_ram[1425] = 245;
    exp_54_ram[1426] = 0;
    exp_54_ram[1427] = 0;
    exp_54_ram[1428] = 250;
    exp_54_ram[1429] = 0;
    exp_54_ram[1430] = 249;
    exp_54_ram[1431] = 254;
    exp_54_ram[1432] = 4;
    exp_54_ram[1433] = 250;
    exp_54_ram[1434] = 0;
    exp_54_ram[1435] = 2;
    exp_54_ram[1436] = 2;
    exp_54_ram[1437] = 249;
    exp_54_ram[1438] = 0;
    exp_54_ram[1439] = 248;
    exp_54_ram[1440] = 0;
    exp_54_ram[1441] = 252;
    exp_54_ram[1442] = 252;
    exp_54_ram[1443] = 0;
    exp_54_ram[1444] = 0;
    exp_54_ram[1445] = 254;
    exp_54_ram[1446] = 250;
    exp_54_ram[1447] = 0;
    exp_54_ram[1448] = 250;
    exp_54_ram[1449] = 250;
    exp_54_ram[1450] = 0;
    exp_54_ram[1451] = 249;
    exp_54_ram[1452] = 1;
    exp_54_ram[1453] = 14;
    exp_54_ram[1454] = 0;
    exp_54_ram[1455] = 0;
    exp_54_ram[1456] = 18;
    exp_54_ram[1457] = 0;
    exp_54_ram[1458] = 0;
    exp_54_ram[1459] = 0;
    exp_54_ram[1460] = 254;
    exp_54_ram[1461] = 16;
    exp_54_ram[1462] = 254;
    exp_54_ram[1463] = 250;
    exp_54_ram[1464] = 0;
    exp_54_ram[1465] = 250;
    exp_54_ram[1466] = 250;
    exp_54_ram[1467] = 0;
    exp_54_ram[1468] = 6;
    exp_54_ram[1469] = 12;
    exp_54_ram[1470] = 254;
    exp_54_ram[1471] = 32;
    exp_54_ram[1472] = 254;
    exp_54_ram[1473] = 250;
    exp_54_ram[1474] = 0;
    exp_54_ram[1475] = 250;
    exp_54_ram[1476] = 10;
    exp_54_ram[1477] = 254;
    exp_54_ram[1478] = 8;
    exp_54_ram[1479] = 254;
    exp_54_ram[1480] = 250;
    exp_54_ram[1481] = 0;
    exp_54_ram[1482] = 250;
    exp_54_ram[1483] = 250;
    exp_54_ram[1484] = 0;
    exp_54_ram[1485] = 6;
    exp_54_ram[1486] = 8;
    exp_54_ram[1487] = 254;
    exp_54_ram[1488] = 4;
    exp_54_ram[1489] = 254;
    exp_54_ram[1490] = 250;
    exp_54_ram[1491] = 0;
    exp_54_ram[1492] = 250;
    exp_54_ram[1493] = 6;
    exp_54_ram[1494] = 254;
    exp_54_ram[1495] = 16;
    exp_54_ram[1496] = 254;
    exp_54_ram[1497] = 250;
    exp_54_ram[1498] = 0;
    exp_54_ram[1499] = 250;
    exp_54_ram[1500] = 5;
    exp_54_ram[1501] = 254;
    exp_54_ram[1502] = 32;
    exp_54_ram[1503] = 254;
    exp_54_ram[1504] = 250;
    exp_54_ram[1505] = 0;
    exp_54_ram[1506] = 250;
    exp_54_ram[1507] = 3;
    exp_54_ram[1508] = 254;
    exp_54_ram[1509] = 16;
    exp_54_ram[1510] = 254;
    exp_54_ram[1511] = 250;
    exp_54_ram[1512] = 0;
    exp_54_ram[1513] = 250;
    exp_54_ram[1514] = 1;
    exp_54_ram[1515] = 0;
    exp_54_ram[1516] = 1;
    exp_54_ram[1517] = 0;
    exp_54_ram[1518] = 0;
    exp_54_ram[1519] = 0;
    exp_54_ram[1520] = 250;
    exp_54_ram[1521] = 0;
    exp_54_ram[1522] = 253;
    exp_54_ram[1523] = 5;
    exp_54_ram[1524] = 98;
    exp_54_ram[1525] = 0;
    exp_54_ram[1526] = 0;
    exp_54_ram[1527] = 23;
    exp_54_ram[1528] = 0;
    exp_54_ram[1529] = 0;
    exp_54_ram[1530] = 0;
    exp_54_ram[1531] = 250;
    exp_54_ram[1532] = 0;
    exp_54_ram[1533] = 7;
    exp_54_ram[1534] = 0;
    exp_54_ram[1535] = 250;
    exp_54_ram[1536] = 0;
    exp_54_ram[1537] = 5;
    exp_54_ram[1538] = 0;
    exp_54_ram[1539] = 1;
    exp_54_ram[1540] = 252;
    exp_54_ram[1541] = 5;
    exp_54_ram[1542] = 250;
    exp_54_ram[1543] = 0;
    exp_54_ram[1544] = 6;
    exp_54_ram[1545] = 0;
    exp_54_ram[1546] = 0;
    exp_54_ram[1547] = 252;
    exp_54_ram[1548] = 3;
    exp_54_ram[1549] = 250;
    exp_54_ram[1550] = 0;
    exp_54_ram[1551] = 6;
    exp_54_ram[1552] = 0;
    exp_54_ram[1553] = 0;
    exp_54_ram[1554] = 252;
    exp_54_ram[1555] = 1;
    exp_54_ram[1556] = 0;
    exp_54_ram[1557] = 252;
    exp_54_ram[1558] = 254;
    exp_54_ram[1559] = 254;
    exp_54_ram[1560] = 254;
    exp_54_ram[1561] = 250;
    exp_54_ram[1562] = 0;
    exp_54_ram[1563] = 5;
    exp_54_ram[1564] = 0;
    exp_54_ram[1565] = 254;
    exp_54_ram[1566] = 2;
    exp_54_ram[1567] = 254;
    exp_54_ram[1568] = 250;
    exp_54_ram[1569] = 0;
    exp_54_ram[1570] = 6;
    exp_54_ram[1571] = 2;
    exp_54_ram[1572] = 250;
    exp_54_ram[1573] = 0;
    exp_54_ram[1574] = 6;
    exp_54_ram[1575] = 0;
    exp_54_ram[1576] = 254;
    exp_54_ram[1577] = 255;
    exp_54_ram[1578] = 254;
    exp_54_ram[1579] = 254;
    exp_54_ram[1580] = 64;
    exp_54_ram[1581] = 0;
    exp_54_ram[1582] = 254;
    exp_54_ram[1583] = 255;
    exp_54_ram[1584] = 254;
    exp_54_ram[1585] = 250;
    exp_54_ram[1586] = 0;
    exp_54_ram[1587] = 6;
    exp_54_ram[1588] = 0;
    exp_54_ram[1589] = 250;
    exp_54_ram[1590] = 0;
    exp_54_ram[1591] = 6;
    exp_54_ram[1592] = 20;
    exp_54_ram[1593] = 254;
    exp_54_ram[1594] = 32;
    exp_54_ram[1595] = 34;
    exp_54_ram[1596] = 254;
    exp_54_ram[1597] = 16;
    exp_54_ram[1598] = 6;
    exp_54_ram[1599] = 249;
    exp_54_ram[1600] = 0;
    exp_54_ram[1601] = 248;
    exp_54_ram[1602] = 0;
    exp_54_ram[1603] = 250;
    exp_54_ram[1604] = 251;
    exp_54_ram[1605] = 65;
    exp_54_ram[1606] = 251;
    exp_54_ram[1607] = 0;
    exp_54_ram[1608] = 64;
    exp_54_ram[1609] = 0;
    exp_54_ram[1610] = 251;
    exp_54_ram[1611] = 1;
    exp_54_ram[1612] = 15;
    exp_54_ram[1613] = 254;
    exp_54_ram[1614] = 0;
    exp_54_ram[1615] = 254;
    exp_54_ram[1616] = 0;
    exp_54_ram[1617] = 254;
    exp_54_ram[1618] = 253;
    exp_54_ram[1619] = 0;
    exp_54_ram[1620] = 0;
    exp_54_ram[1621] = 250;
    exp_54_ram[1622] = 253;
    exp_54_ram[1623] = 250;
    exp_54_ram[1624] = 250;
    exp_54_ram[1625] = 148;
    exp_54_ram[1626] = 252;
    exp_54_ram[1627] = 27;
    exp_54_ram[1628] = 254;
    exp_54_ram[1629] = 4;
    exp_54_ram[1630] = 0;
    exp_54_ram[1631] = 249;
    exp_54_ram[1632] = 0;
    exp_54_ram[1633] = 248;
    exp_54_ram[1634] = 0;
    exp_54_ram[1635] = 15;
    exp_54_ram[1636] = 3;
    exp_54_ram[1637] = 254;
    exp_54_ram[1638] = 8;
    exp_54_ram[1639] = 2;
    exp_54_ram[1640] = 249;
    exp_54_ram[1641] = 0;
    exp_54_ram[1642] = 248;
    exp_54_ram[1643] = 0;
    exp_54_ram[1644] = 1;
    exp_54_ram[1645] = 65;
    exp_54_ram[1646] = 1;
    exp_54_ram[1647] = 249;
    exp_54_ram[1648] = 0;
    exp_54_ram[1649] = 248;
    exp_54_ram[1650] = 0;
    exp_54_ram[1651] = 250;
    exp_54_ram[1652] = 251;
    exp_54_ram[1653] = 65;
    exp_54_ram[1654] = 251;
    exp_54_ram[1655] = 0;
    exp_54_ram[1656] = 64;
    exp_54_ram[1657] = 0;
    exp_54_ram[1658] = 251;
    exp_54_ram[1659] = 1;
    exp_54_ram[1660] = 15;
    exp_54_ram[1661] = 254;
    exp_54_ram[1662] = 0;
    exp_54_ram[1663] = 254;
    exp_54_ram[1664] = 0;
    exp_54_ram[1665] = 254;
    exp_54_ram[1666] = 253;
    exp_54_ram[1667] = 0;
    exp_54_ram[1668] = 0;
    exp_54_ram[1669] = 250;
    exp_54_ram[1670] = 253;
    exp_54_ram[1671] = 250;
    exp_54_ram[1672] = 250;
    exp_54_ram[1673] = 136;
    exp_54_ram[1674] = 252;
    exp_54_ram[1675] = 15;
    exp_54_ram[1676] = 254;
    exp_54_ram[1677] = 32;
    exp_54_ram[1678] = 14;
    exp_54_ram[1679] = 254;
    exp_54_ram[1680] = 16;
    exp_54_ram[1681] = 4;
    exp_54_ram[1682] = 249;
    exp_54_ram[1683] = 0;
    exp_54_ram[1684] = 248;
    exp_54_ram[1685] = 0;
    exp_54_ram[1686] = 254;
    exp_54_ram[1687] = 0;
    exp_54_ram[1688] = 254;
    exp_54_ram[1689] = 0;
    exp_54_ram[1690] = 254;
    exp_54_ram[1691] = 253;
    exp_54_ram[1692] = 0;
    exp_54_ram[1693] = 250;
    exp_54_ram[1694] = 253;
    exp_54_ram[1695] = 250;
    exp_54_ram[1696] = 250;
    exp_54_ram[1697] = 130;
    exp_54_ram[1698] = 252;
    exp_54_ram[1699] = 9;
    exp_54_ram[1700] = 254;
    exp_54_ram[1701] = 4;
    exp_54_ram[1702] = 0;
    exp_54_ram[1703] = 249;
    exp_54_ram[1704] = 0;
    exp_54_ram[1705] = 248;
    exp_54_ram[1706] = 0;
    exp_54_ram[1707] = 15;
    exp_54_ram[1708] = 3;
    exp_54_ram[1709] = 254;
    exp_54_ram[1710] = 8;
    exp_54_ram[1711] = 2;
    exp_54_ram[1712] = 249;
    exp_54_ram[1713] = 0;
    exp_54_ram[1714] = 248;
    exp_54_ram[1715] = 0;
    exp_54_ram[1716] = 1;
    exp_54_ram[1717] = 1;
    exp_54_ram[1718] = 1;
    exp_54_ram[1719] = 249;
    exp_54_ram[1720] = 0;
    exp_54_ram[1721] = 248;
    exp_54_ram[1722] = 0;
    exp_54_ram[1723] = 252;
    exp_54_ram[1724] = 254;
    exp_54_ram[1725] = 0;
    exp_54_ram[1726] = 254;
    exp_54_ram[1727] = 0;
    exp_54_ram[1728] = 254;
    exp_54_ram[1729] = 253;
    exp_54_ram[1730] = 0;
    exp_54_ram[1731] = 252;
    exp_54_ram[1732] = 250;
    exp_54_ram[1733] = 253;
    exp_54_ram[1734] = 250;
    exp_54_ram[1735] = 250;
    exp_54_ram[1736] = 249;
    exp_54_ram[1737] = 252;
    exp_54_ram[1738] = 250;
    exp_54_ram[1739] = 0;
    exp_54_ram[1740] = 250;
    exp_54_ram[1741] = 48;
    exp_54_ram[1742] = 0;
    exp_54_ram[1743] = 252;
    exp_54_ram[1744] = 254;
    exp_54_ram[1745] = 0;
    exp_54_ram[1746] = 4;
    exp_54_ram[1747] = 2;
    exp_54_ram[1748] = 253;
    exp_54_ram[1749] = 0;
    exp_54_ram[1750] = 252;
    exp_54_ram[1751] = 250;
    exp_54_ram[1752] = 250;
    exp_54_ram[1753] = 0;
    exp_54_ram[1754] = 250;
    exp_54_ram[1755] = 2;
    exp_54_ram[1756] = 0;
    exp_54_ram[1757] = 253;
    exp_54_ram[1758] = 0;
    exp_54_ram[1759] = 252;
    exp_54_ram[1760] = 254;
    exp_54_ram[1761] = 252;
    exp_54_ram[1762] = 249;
    exp_54_ram[1763] = 0;
    exp_54_ram[1764] = 248;
    exp_54_ram[1765] = 0;
    exp_54_ram[1766] = 15;
    exp_54_ram[1767] = 253;
    exp_54_ram[1768] = 0;
    exp_54_ram[1769] = 252;
    exp_54_ram[1770] = 250;
    exp_54_ram[1771] = 250;
    exp_54_ram[1772] = 0;
    exp_54_ram[1773] = 250;
    exp_54_ram[1774] = 0;
    exp_54_ram[1775] = 254;
    exp_54_ram[1776] = 0;
    exp_54_ram[1777] = 4;
    exp_54_ram[1778] = 2;
    exp_54_ram[1779] = 253;
    exp_54_ram[1780] = 0;
    exp_54_ram[1781] = 252;
    exp_54_ram[1782] = 250;
    exp_54_ram[1783] = 250;
    exp_54_ram[1784] = 0;
    exp_54_ram[1785] = 250;
    exp_54_ram[1786] = 2;
    exp_54_ram[1787] = 0;
    exp_54_ram[1788] = 253;
    exp_54_ram[1789] = 0;
    exp_54_ram[1790] = 252;
    exp_54_ram[1791] = 254;
    exp_54_ram[1792] = 252;
    exp_54_ram[1793] = 250;
    exp_54_ram[1794] = 0;
    exp_54_ram[1795] = 250;
    exp_54_ram[1796] = 35;
    exp_54_ram[1797] = 249;
    exp_54_ram[1798] = 0;
    exp_54_ram[1799] = 248;
    exp_54_ram[1800] = 0;
    exp_54_ram[1801] = 252;
    exp_54_ram[1802] = 254;
    exp_54_ram[1803] = 0;
    exp_54_ram[1804] = 254;
    exp_54_ram[1805] = 0;
    exp_54_ram[1806] = 255;
    exp_54_ram[1807] = 0;
    exp_54_ram[1808] = 253;
    exp_54_ram[1809] = 143;
    exp_54_ram[1810] = 252;
    exp_54_ram[1811] = 254;
    exp_54_ram[1812] = 64;
    exp_54_ram[1813] = 0;
    exp_54_ram[1814] = 252;
    exp_54_ram[1815] = 254;
    exp_54_ram[1816] = 0;
    exp_54_ram[1817] = 0;
    exp_54_ram[1818] = 252;
    exp_54_ram[1819] = 254;
    exp_54_ram[1820] = 0;
    exp_54_ram[1821] = 6;
    exp_54_ram[1822] = 2;
    exp_54_ram[1823] = 253;
    exp_54_ram[1824] = 0;
    exp_54_ram[1825] = 252;
    exp_54_ram[1826] = 250;
    exp_54_ram[1827] = 250;
    exp_54_ram[1828] = 0;
    exp_54_ram[1829] = 250;
    exp_54_ram[1830] = 2;
    exp_54_ram[1831] = 0;
    exp_54_ram[1832] = 252;
    exp_54_ram[1833] = 0;
    exp_54_ram[1834] = 252;
    exp_54_ram[1835] = 254;
    exp_54_ram[1836] = 252;
    exp_54_ram[1837] = 3;
    exp_54_ram[1838] = 253;
    exp_54_ram[1839] = 0;
    exp_54_ram[1840] = 252;
    exp_54_ram[1841] = 0;
    exp_54_ram[1842] = 253;
    exp_54_ram[1843] = 0;
    exp_54_ram[1844] = 252;
    exp_54_ram[1845] = 250;
    exp_54_ram[1846] = 250;
    exp_54_ram[1847] = 0;
    exp_54_ram[1848] = 250;
    exp_54_ram[1849] = 0;
    exp_54_ram[1850] = 253;
    exp_54_ram[1851] = 0;
    exp_54_ram[1852] = 2;
    exp_54_ram[1853] = 254;
    exp_54_ram[1854] = 64;
    exp_54_ram[1855] = 250;
    exp_54_ram[1856] = 254;
    exp_54_ram[1857] = 255;
    exp_54_ram[1858] = 254;
    exp_54_ram[1859] = 250;
    exp_54_ram[1860] = 254;
    exp_54_ram[1861] = 0;
    exp_54_ram[1862] = 4;
    exp_54_ram[1863] = 2;
    exp_54_ram[1864] = 253;
    exp_54_ram[1865] = 0;
    exp_54_ram[1866] = 252;
    exp_54_ram[1867] = 250;
    exp_54_ram[1868] = 250;
    exp_54_ram[1869] = 0;
    exp_54_ram[1870] = 250;
    exp_54_ram[1871] = 2;
    exp_54_ram[1872] = 0;
    exp_54_ram[1873] = 252;
    exp_54_ram[1874] = 0;
    exp_54_ram[1875] = 252;
    exp_54_ram[1876] = 254;
    exp_54_ram[1877] = 252;
    exp_54_ram[1878] = 250;
    exp_54_ram[1879] = 0;
    exp_54_ram[1880] = 250;
    exp_54_ram[1881] = 13;
    exp_54_ram[1882] = 0;
    exp_54_ram[1883] = 254;
    exp_54_ram[1884] = 254;
    exp_54_ram[1885] = 2;
    exp_54_ram[1886] = 254;
    exp_54_ram[1887] = 249;
    exp_54_ram[1888] = 0;
    exp_54_ram[1889] = 248;
    exp_54_ram[1890] = 0;
    exp_54_ram[1891] = 0;
    exp_54_ram[1892] = 254;
    exp_54_ram[1893] = 0;
    exp_54_ram[1894] = 254;
    exp_54_ram[1895] = 0;
    exp_54_ram[1896] = 254;
    exp_54_ram[1897] = 1;
    exp_54_ram[1898] = 0;
    exp_54_ram[1899] = 250;
    exp_54_ram[1900] = 253;
    exp_54_ram[1901] = 250;
    exp_54_ram[1902] = 250;
    exp_54_ram[1903] = 207;
    exp_54_ram[1904] = 252;
    exp_54_ram[1905] = 250;
    exp_54_ram[1906] = 0;
    exp_54_ram[1907] = 250;
    exp_54_ram[1908] = 7;
    exp_54_ram[1909] = 253;
    exp_54_ram[1910] = 0;
    exp_54_ram[1911] = 252;
    exp_54_ram[1912] = 250;
    exp_54_ram[1913] = 250;
    exp_54_ram[1914] = 0;
    exp_54_ram[1915] = 250;
    exp_54_ram[1916] = 2;
    exp_54_ram[1917] = 0;
    exp_54_ram[1918] = 250;
    exp_54_ram[1919] = 0;
    exp_54_ram[1920] = 250;
    exp_54_ram[1921] = 3;
    exp_54_ram[1922] = 250;
    exp_54_ram[1923] = 0;
    exp_54_ram[1924] = 253;
    exp_54_ram[1925] = 0;
    exp_54_ram[1926] = 252;
    exp_54_ram[1927] = 250;
    exp_54_ram[1928] = 250;
    exp_54_ram[1929] = 0;
    exp_54_ram[1930] = 250;
    exp_54_ram[1931] = 0;
    exp_54_ram[1932] = 250;
    exp_54_ram[1933] = 0;
    exp_54_ram[1934] = 250;
    exp_54_ram[1935] = 0;
    exp_54_ram[1936] = 250;
    exp_54_ram[1937] = 0;
    exp_54_ram[1938] = 222;
    exp_54_ram[1939] = 253;
    exp_54_ram[1940] = 250;
    exp_54_ram[1941] = 0;
    exp_54_ram[1942] = 250;
    exp_54_ram[1943] = 255;
    exp_54_ram[1944] = 0;
    exp_54_ram[1945] = 253;
    exp_54_ram[1946] = 250;
    exp_54_ram[1947] = 250;
    exp_54_ram[1948] = 0;
    exp_54_ram[1949] = 250;
    exp_54_ram[1950] = 0;
    exp_54_ram[1951] = 0;
    exp_54_ram[1952] = 253;
    exp_54_ram[1953] = 0;
    exp_54_ram[1954] = 7;
    exp_54_ram[1955] = 7;
    exp_54_ram[1956] = 8;
    exp_54_ram[1957] = 0;
    exp_54_ram[1958] = 251;
    exp_54_ram[1959] = 2;
    exp_54_ram[1960] = 2;
    exp_54_ram[1961] = 3;
    exp_54_ram[1962] = 252;
    exp_54_ram[1963] = 0;
    exp_54_ram[1964] = 0;
    exp_54_ram[1965] = 0;
    exp_54_ram[1966] = 0;
    exp_54_ram[1967] = 0;
    exp_54_ram[1968] = 1;
    exp_54_ram[1969] = 1;
    exp_54_ram[1970] = 2;
    exp_54_ram[1971] = 252;
    exp_54_ram[1972] = 253;
    exp_54_ram[1973] = 254;
    exp_54_ram[1974] = 254;
    exp_54_ram[1975] = 254;
    exp_54_ram[1976] = 254;
    exp_54_ram[1977] = 253;
    exp_54_ram[1978] = 255;
    exp_54_ram[1979] = 0;
    exp_54_ram[1980] = 0;
    exp_54_ram[1981] = 206;
    exp_54_ram[1982] = 208;
    exp_54_ram[1983] = 254;
    exp_54_ram[1984] = 254;
    exp_54_ram[1985] = 0;
    exp_54_ram[1986] = 2;
    exp_54_ram[1987] = 2;
    exp_54_ram[1988] = 5;
    exp_54_ram[1989] = 0;
    exp_54_ram[1990] = 254;
    exp_54_ram[1991] = 0;
    exp_54_ram[1992] = 0;
    exp_54_ram[1993] = 2;
    exp_54_ram[1994] = 0;
    exp_54_ram[1995] = 254;
    exp_54_ram[1996] = 254;
    exp_54_ram[1997] = 0;
    exp_54_ram[1998] = 13;
    exp_54_ram[1999] = 0;
    exp_54_ram[2000] = 0;
    exp_54_ram[2001] = 195;
    exp_54_ram[2002] = 0;
    exp_54_ram[2003] = 1;
    exp_54_ram[2004] = 1;
    exp_54_ram[2005] = 2;
    exp_54_ram[2006] = 0;
    exp_54_ram[2007] = 246;
    exp_54_ram[2008] = 8;
    exp_54_ram[2009] = 8;
    exp_54_ram[2010] = 8;
    exp_54_ram[2011] = 10;
    exp_54_ram[2012] = 0;
    exp_54_ram[2013] = 1;
    exp_54_ram[2014] = 252;
    exp_54_ram[2015] = 0;
    exp_54_ram[2016] = 252;
    exp_54_ram[2017] = 1;
    exp_54_ram[2018] = 252;
    exp_54_ram[2019] = 0;
    exp_54_ram[2020] = 250;
    exp_54_ram[2021] = 250;
    exp_54_ram[2022] = 250;
    exp_54_ram[2023] = 252;
    exp_54_ram[2024] = 251;
    exp_54_ram[2025] = 251;
    exp_54_ram[2026] = 251;
    exp_54_ram[2027] = 252;
    exp_54_ram[2028] = 252;
    exp_54_ram[2029] = 252;
    exp_54_ram[2030] = 252;
    exp_54_ram[2031] = 253;
    exp_54_ram[2032] = 253;
    exp_54_ram[2033] = 246;
    exp_54_ram[2034] = 247;
    exp_54_ram[2035] = 247;
    exp_54_ram[2036] = 246;
    exp_54_ram[2037] = 246;
    exp_54_ram[2038] = 246;
    exp_54_ram[2039] = 246;
    exp_54_ram[2040] = 246;
    exp_54_ram[2041] = 248;
    exp_54_ram[2042] = 246;
    exp_54_ram[2043] = 0;
    exp_54_ram[2044] = 80;
    exp_54_ram[2045] = 254;
    exp_54_ram[2046] = 254;
    exp_54_ram[2047] = 251;
    exp_54_ram[2048] = 254;
    exp_54_ram[2049] = 254;
    exp_54_ram[2050] = 0;
    exp_54_ram[2051] = 12;
    exp_54_ram[2052] = 252;
    exp_54_ram[2053] = 252;
    exp_54_ram[2054] = 64;
    exp_54_ram[2055] = 252;
    exp_54_ram[2056] = 251;
    exp_54_ram[2057] = 251;
    exp_54_ram[2058] = 251;
    exp_54_ram[2059] = 252;
    exp_54_ram[2060] = 252;
    exp_54_ram[2061] = 252;
    exp_54_ram[2062] = 252;
    exp_54_ram[2063] = 253;
    exp_54_ram[2064] = 253;
    exp_54_ram[2065] = 246;
    exp_54_ram[2066] = 247;
    exp_54_ram[2067] = 247;
    exp_54_ram[2068] = 246;
    exp_54_ram[2069] = 246;
    exp_54_ram[2070] = 246;
    exp_54_ram[2071] = 246;
    exp_54_ram[2072] = 246;
    exp_54_ram[2073] = 248;
    exp_54_ram[2074] = 246;
    exp_54_ram[2075] = 0;
    exp_54_ram[2076] = 72;
    exp_54_ram[2077] = 254;
    exp_54_ram[2078] = 254;
    exp_54_ram[2079] = 1;
    exp_54_ram[2080] = 250;
    exp_54_ram[2081] = 0;
    exp_54_ram[2082] = 250;
    exp_54_ram[2083] = 1;
    exp_54_ram[2084] = 248;
    exp_54_ram[2085] = 0;
    exp_54_ram[2086] = 248;
    exp_54_ram[2087] = 248;
    exp_54_ram[2088] = 248;
    exp_54_ram[2089] = 252;
    exp_54_ram[2090] = 249;
    exp_54_ram[2091] = 249;
    exp_54_ram[2092] = 249;
    exp_54_ram[2093] = 249;
    exp_54_ram[2094] = 250;
    exp_54_ram[2095] = 250;
    exp_54_ram[2096] = 250;
    exp_54_ram[2097] = 250;
    exp_54_ram[2098] = 251;
    exp_54_ram[2099] = 246;
    exp_54_ram[2100] = 247;
    exp_54_ram[2101] = 247;
    exp_54_ram[2102] = 246;
    exp_54_ram[2103] = 246;
    exp_54_ram[2104] = 246;
    exp_54_ram[2105] = 246;
    exp_54_ram[2106] = 246;
    exp_54_ram[2107] = 248;
    exp_54_ram[2108] = 246;
    exp_54_ram[2109] = 0;
    exp_54_ram[2110] = 63;
    exp_54_ram[2111] = 254;
    exp_54_ram[2112] = 254;
    exp_54_ram[2113] = 249;
    exp_54_ram[2114] = 254;
    exp_54_ram[2115] = 254;
    exp_54_ram[2116] = 0;
    exp_54_ram[2117] = 123;
    exp_54_ram[2118] = 249;
    exp_54_ram[2119] = 250;
    exp_54_ram[2120] = 64;
    exp_54_ram[2121] = 248;
    exp_54_ram[2122] = 249;
    exp_54_ram[2123] = 249;
    exp_54_ram[2124] = 249;
    exp_54_ram[2125] = 249;
    exp_54_ram[2126] = 250;
    exp_54_ram[2127] = 250;
    exp_54_ram[2128] = 250;
    exp_54_ram[2129] = 250;
    exp_54_ram[2130] = 251;
    exp_54_ram[2131] = 246;
    exp_54_ram[2132] = 247;
    exp_54_ram[2133] = 247;
    exp_54_ram[2134] = 246;
    exp_54_ram[2135] = 246;
    exp_54_ram[2136] = 246;
    exp_54_ram[2137] = 246;
    exp_54_ram[2138] = 246;
    exp_54_ram[2139] = 248;
    exp_54_ram[2140] = 246;
    exp_54_ram[2141] = 0;
    exp_54_ram[2142] = 55;
    exp_54_ram[2143] = 254;
    exp_54_ram[2144] = 254;
    exp_54_ram[2145] = 0;
    exp_54_ram[2146] = 0;
    exp_54_ram[2147] = 0;
    exp_54_ram[2148] = 0;
    exp_54_ram[2149] = 1;
    exp_54_ram[2150] = 1;
    exp_54_ram[2151] = 1;
    exp_54_ram[2152] = 1;
    exp_54_ram[2153] = 2;
    exp_54_ram[2154] = 246;
    exp_54_ram[2155] = 247;
    exp_54_ram[2156] = 247;
    exp_54_ram[2157] = 246;
    exp_54_ram[2158] = 246;
    exp_54_ram[2159] = 246;
    exp_54_ram[2160] = 246;
    exp_54_ram[2161] = 246;
    exp_54_ram[2162] = 248;
    exp_54_ram[2163] = 246;
    exp_54_ram[2164] = 0;
    exp_54_ram[2165] = 50;
    exp_54_ram[2166] = 252;
    exp_54_ram[2167] = 252;
    exp_54_ram[2168] = 254;
    exp_54_ram[2169] = 253;
    exp_54_ram[2170] = 4;
    exp_54_ram[2171] = 254;
    exp_54_ram[2172] = 253;
    exp_54_ram[2173] = 0;
    exp_54_ram[2174] = 254;
    exp_54_ram[2175] = 253;
    exp_54_ram[2176] = 2;
    exp_54_ram[2177] = 254;
    exp_54_ram[2178] = 253;
    exp_54_ram[2179] = 0;
    exp_54_ram[2180] = 254;
    exp_54_ram[2181] = 253;
    exp_54_ram[2182] = 0;
    exp_54_ram[2183] = 254;
    exp_54_ram[2184] = 253;
    exp_54_ram[2185] = 0;
    exp_54_ram[2186] = 0;
    exp_54_ram[2187] = 0;
    exp_54_ram[2188] = 0;
    exp_54_ram[2189] = 0;
    exp_54_ram[2190] = 9;
    exp_54_ram[2191] = 9;
    exp_54_ram[2192] = 9;
    exp_54_ram[2193] = 10;
    exp_54_ram[2194] = 0;
    exp_54_ram[2195] = 248;
    exp_54_ram[2196] = 6;
    exp_54_ram[2197] = 6;
    exp_54_ram[2198] = 8;
    exp_54_ram[2199] = 250;
    exp_54_ram[2200] = 250;
    exp_54_ram[2201] = 252;
    exp_54_ram[2202] = 251;
    exp_54_ram[2203] = 251;
    exp_54_ram[2204] = 0;
    exp_54_ram[2205] = 101;
    exp_54_ram[2206] = 252;
    exp_54_ram[2207] = 253;
    exp_54_ram[2208] = 253;
    exp_54_ram[2209] = 253;
    exp_54_ram[2210] = 253;
    exp_54_ram[2211] = 254;
    exp_54_ram[2212] = 254;
    exp_54_ram[2213] = 254;
    exp_54_ram[2214] = 254;
    exp_54_ram[2215] = 248;
    exp_54_ram[2216] = 249;
    exp_54_ram[2217] = 249;
    exp_54_ram[2218] = 248;
    exp_54_ram[2219] = 248;
    exp_54_ram[2220] = 248;
    exp_54_ram[2221] = 248;
    exp_54_ram[2222] = 248;
    exp_54_ram[2223] = 250;
    exp_54_ram[2224] = 248;
    exp_54_ram[2225] = 0;
    exp_54_ram[2226] = 201;
    exp_54_ram[2227] = 0;
    exp_54_ram[2228] = 0;
    exp_54_ram[2229] = 7;
    exp_54_ram[2230] = 7;
    exp_54_ram[2231] = 8;
    exp_54_ram[2232] = 0;
    exp_54_ram[2233] = 254;
    exp_54_ram[2234] = 0;
    exp_54_ram[2235] = 2;
    exp_54_ram[2236] = 128;
    exp_54_ram[2237] = 254;
    exp_54_ram[2238] = 128;
    exp_54_ram[2239] = 0;
    exp_54_ram[2240] = 254;
    exp_54_ram[2241] = 254;
    exp_54_ram[2242] = 0;
    exp_54_ram[2243] = 0;
    exp_54_ram[2244] = 254;
    exp_54_ram[2245] = 0;
    exp_54_ram[2246] = 0;
    exp_54_ram[2247] = 0;
    exp_54_ram[2248] = 0;
    exp_54_ram[2249] = 0;
    exp_54_ram[2250] = 0;
    exp_54_ram[2251] = 0;
    exp_54_ram[2252] = 0;
    exp_54_ram[2253] = 0;
    exp_54_ram[2254] = 0;
    exp_54_ram[2255] = 1;
    exp_54_ram[2256] = 2;
    exp_54_ram[2257] = 0;
    exp_54_ram[2258] = 254;
    exp_54_ram[2259] = 0;
    exp_54_ram[2260] = 0;
    exp_54_ram[2261] = 2;
    exp_54_ram[2262] = 254;
    exp_54_ram[2263] = 254;
    exp_54_ram[2264] = 254;
    exp_54_ram[2265] = 254;
    exp_54_ram[2266] = 254;
    exp_54_ram[2267] = 254;
    exp_54_ram[2268] = 254;
    exp_54_ram[2269] = 254;
    exp_54_ram[2270] = 64;
    exp_54_ram[2271] = 0;
    exp_54_ram[2272] = 1;
    exp_54_ram[2273] = 64;
    exp_54_ram[2274] = 65;
    exp_54_ram[2275] = 0;
    exp_54_ram[2276] = 0;
    exp_54_ram[2277] = 0;
    exp_54_ram[2278] = 0;
    exp_54_ram[2279] = 0;
    exp_54_ram[2280] = 168;
    exp_54_ram[2281] = 0;
    exp_54_ram[2282] = 0;
    exp_54_ram[2283] = 0;
    exp_54_ram[2284] = 0;
    exp_54_ram[2285] = 1;
    exp_54_ram[2286] = 1;
    exp_54_ram[2287] = 2;
    exp_54_ram[2288] = 0;
    exp_54_ram[2289] = 254;
    exp_54_ram[2290] = 0;
    exp_54_ram[2291] = 2;
    exp_54_ram[2292] = 254;
    exp_54_ram[2293] = 254;
    exp_54_ram[2294] = 0;
    exp_54_ram[2295] = 2;
    exp_54_ram[2296] = 254;
    exp_54_ram[2297] = 6;
    exp_54_ram[2298] = 2;
    exp_54_ram[2299] = 0;
    exp_54_ram[2300] = 254;
    exp_54_ram[2301] = 25;
    exp_54_ram[2302] = 2;
    exp_54_ram[2303] = 0;
    exp_54_ram[2304] = 0;
    exp_54_ram[2305] = 0;
    exp_54_ram[2306] = 0;
    exp_54_ram[2307] = 0;
    exp_54_ram[2308] = 1;
    exp_54_ram[2309] = 2;
    exp_54_ram[2310] = 0;
    exp_54_ram[2311] = 254;
    exp_54_ram[2312] = 0;
    exp_54_ram[2313] = 0;
    exp_54_ram[2314] = 2;
    exp_54_ram[2315] = 254;
    exp_54_ram[2316] = 254;
    exp_54_ram[2317] = 249;
    exp_54_ram[2318] = 0;
    exp_54_ram[2319] = 0;
    exp_54_ram[2320] = 22;
    exp_54_ram[2321] = 0;
    exp_54_ram[2322] = 22;
    exp_54_ram[2323] = 0;
    exp_54_ram[2324] = 1;
    exp_54_ram[2325] = 1;
    exp_54_ram[2326] = 2;
    exp_54_ram[2327] = 0;
    exp_54_ram[2328] = 254;
    exp_54_ram[2329] = 0;
    exp_54_ram[2330] = 0;
    exp_54_ram[2331] = 2;
    exp_54_ram[2332] = 254;
    exp_54_ram[2333] = 254;
    exp_54_ram[2334] = 254;
    exp_54_ram[2335] = 0;
    exp_54_ram[2336] = 2;
    exp_54_ram[2337] = 254;
    exp_54_ram[2338] = 0;
    exp_54_ram[2339] = 0;
    exp_54_ram[2340] = 254;
    exp_54_ram[2341] = 0;
    exp_54_ram[2342] = 0;
    exp_54_ram[2343] = 254;
    exp_54_ram[2344] = 0;
    exp_54_ram[2345] = 0;
    exp_54_ram[2346] = 1;
    exp_54_ram[2347] = 3;
    exp_54_ram[2348] = 254;
    exp_54_ram[2349] = 0;
    exp_54_ram[2350] = 2;
    exp_54_ram[2351] = 254;
    exp_54_ram[2352] = 240;
    exp_54_ram[2353] = 0;
    exp_54_ram[2354] = 0;
    exp_54_ram[2355] = 1;
    exp_54_ram[2356] = 1;
    exp_54_ram[2357] = 1;
    exp_54_ram[2358] = 0;
    exp_54_ram[2359] = 1;
    exp_54_ram[2360] = 0;
    exp_54_ram[2361] = 1;
    exp_54_ram[2362] = 1;
    exp_54_ram[2363] = 2;
    exp_54_ram[2364] = 0;
    exp_54_ram[2365] = 249;
    exp_54_ram[2366] = 6;
    exp_54_ram[2367] = 6;
    exp_54_ram[2368] = 6;
    exp_54_ram[2369] = 7;
    exp_54_ram[2370] = 5;
    exp_54_ram[2371] = 5;
    exp_54_ram[2372] = 5;
    exp_54_ram[2373] = 5;
    exp_54_ram[2374] = 5;
    exp_54_ram[2375] = 5;
    exp_54_ram[2376] = 5;
    exp_54_ram[2377] = 5;
    exp_54_ram[2378] = 3;
    exp_54_ram[2379] = 7;
    exp_54_ram[2380] = 0;
    exp_54_ram[2381] = 0;
    exp_54_ram[2382] = 0;
    exp_54_ram[2383] = 250;
    exp_54_ram[2384] = 251;
    exp_54_ram[2385] = 123;
    exp_54_ram[2386] = 250;
    exp_54_ram[2387] = 1;
    exp_54_ram[2388] = 250;
    exp_54_ram[2389] = 250;
    exp_54_ram[2390] = 118;
    exp_54_ram[2391] = 251;
    exp_54_ram[2392] = 6;
    exp_54_ram[2393] = 251;
    exp_54_ram[2394] = 235;
    exp_54_ram[2395] = 0;
    exp_54_ram[2396] = 0;
    exp_54_ram[2397] = 24;
    exp_54_ram[2398] = 2;
    exp_54_ram[2399] = 248;
    exp_54_ram[2400] = 248;
    exp_54_ram[2401] = 251;
    exp_54_ram[2402] = 251;
    exp_54_ram[2403] = 249;
    exp_54_ram[2404] = 249;
    exp_54_ram[2405] = 0;
    exp_54_ram[2406] = 0;
    exp_54_ram[2407] = 0;
    exp_54_ram[2408] = 0;
    exp_54_ram[2409] = 0;
    exp_54_ram[2410] = 0;
    exp_54_ram[2411] = 0;
    exp_54_ram[2412] = 0;
    exp_54_ram[2413] = 250;
    exp_54_ram[2414] = 250;
    exp_54_ram[2415] = 251;
    exp_54_ram[2416] = 0;
    exp_54_ram[2417] = 250;
    exp_54_ram[2418] = 248;
    exp_54_ram[2419] = 0;
    exp_54_ram[2420] = 250;
    exp_54_ram[2421] = 1;
    exp_54_ram[2422] = 0;
    exp_54_ram[2423] = 251;
    exp_54_ram[2424] = 6;
    exp_54_ram[2425] = 251;
    exp_54_ram[2426] = 251;
    exp_54_ram[2427] = 231;
    exp_54_ram[2428] = 0;
    exp_54_ram[2429] = 0;
    exp_54_ram[2430] = 24;
    exp_54_ram[2431] = 2;
    exp_54_ram[2432] = 0;
    exp_54_ram[2433] = 0;
    exp_54_ram[2434] = 251;
    exp_54_ram[2435] = 251;
    exp_54_ram[2436] = 1;
    exp_54_ram[2437] = 0;
    exp_54_ram[2438] = 0;
    exp_54_ram[2439] = 1;
    exp_54_ram[2440] = 0;
    exp_54_ram[2441] = 0;
    exp_54_ram[2442] = 250;
    exp_54_ram[2443] = 250;
    exp_54_ram[2444] = 251;
    exp_54_ram[2445] = 0;
    exp_54_ram[2446] = 250;
    exp_54_ram[2447] = 249;
    exp_54_ram[2448] = 0;
    exp_54_ram[2449] = 0;
    exp_54_ram[2450] = 255;
    exp_54_ram[2451] = 0;
    exp_54_ram[2452] = 24;
    exp_54_ram[2453] = 2;
    exp_54_ram[2454] = 0;
    exp_54_ram[2455] = 65;
    exp_54_ram[2456] = 0;
    exp_54_ram[2457] = 251;
    exp_54_ram[2458] = 251;
    exp_54_ram[2459] = 1;
    exp_54_ram[2460] = 0;
    exp_54_ram[2461] = 0;
    exp_54_ram[2462] = 1;
    exp_54_ram[2463] = 0;
    exp_54_ram[2464] = 0;
    exp_54_ram[2465] = 250;
    exp_54_ram[2466] = 250;
    exp_54_ram[2467] = 0;
    exp_54_ram[2468] = 0;
    exp_54_ram[2469] = 225;
    exp_54_ram[2470] = 2;
    exp_54_ram[2471] = 0;
    exp_54_ram[2472] = 65;
    exp_54_ram[2473] = 0;
    exp_54_ram[2474] = 251;
    exp_54_ram[2475] = 251;
    exp_54_ram[2476] = 1;
    exp_54_ram[2477] = 0;
    exp_54_ram[2478] = 0;
    exp_54_ram[2479] = 1;
    exp_54_ram[2480] = 0;
    exp_54_ram[2481] = 0;
    exp_54_ram[2482] = 250;
    exp_54_ram[2483] = 250;
    exp_54_ram[2484] = 0;
    exp_54_ram[2485] = 0;
    exp_54_ram[2486] = 0;
    exp_54_ram[2487] = 64;
    exp_54_ram[2488] = 0;
    exp_54_ram[2489] = 0;
    exp_54_ram[2490] = 65;
    exp_54_ram[2491] = 0;
    exp_54_ram[2492] = 251;
    exp_54_ram[2493] = 251;
    exp_54_ram[2494] = 1;
    exp_54_ram[2495] = 0;
    exp_54_ram[2496] = 0;
    exp_54_ram[2497] = 1;
    exp_54_ram[2498] = 0;
    exp_54_ram[2499] = 0;
    exp_54_ram[2500] = 250;
    exp_54_ram[2501] = 250;
    exp_54_ram[2502] = 0;
    exp_54_ram[2503] = 0;
    exp_54_ram[2504] = 65;
    exp_54_ram[2505] = 0;
    exp_54_ram[2506] = 251;
    exp_54_ram[2507] = 251;
    exp_54_ram[2508] = 1;
    exp_54_ram[2509] = 0;
    exp_54_ram[2510] = 0;
    exp_54_ram[2511] = 1;
    exp_54_ram[2512] = 0;
    exp_54_ram[2513] = 0;
    exp_54_ram[2514] = 250;
    exp_54_ram[2515] = 250;
    exp_54_ram[2516] = 251;
    exp_54_ram[2517] = 251;
    exp_54_ram[2518] = 0;
    exp_54_ram[2519] = 0;
    exp_54_ram[2520] = 6;
    exp_54_ram[2521] = 6;
    exp_54_ram[2522] = 6;
    exp_54_ram[2523] = 6;
    exp_54_ram[2524] = 5;
    exp_54_ram[2525] = 5;
    exp_54_ram[2526] = 5;
    exp_54_ram[2527] = 5;
    exp_54_ram[2528] = 4;
    exp_54_ram[2529] = 4;
    exp_54_ram[2530] = 4;
    exp_54_ram[2531] = 4;
    exp_54_ram[2532] = 3;
    exp_54_ram[2533] = 7;
    exp_54_ram[2534] = 0;
    exp_54_ram[2535] = 246;
    exp_54_ram[2536] = 8;
    exp_54_ram[2537] = 8;
    exp_54_ram[2538] = 8;
    exp_54_ram[2539] = 9;
    exp_54_ram[2540] = 9;
    exp_54_ram[2541] = 10;
    exp_54_ram[2542] = 248;
    exp_54_ram[2543] = 249;
    exp_54_ram[2544] = 0;
    exp_54_ram[2545] = 0;
    exp_54_ram[2546] = 0;
    exp_54_ram[2547] = 0;
    exp_54_ram[2548] = 1;
    exp_54_ram[2549] = 1;
    exp_54_ram[2550] = 1;
    exp_54_ram[2551] = 1;
    exp_54_ram[2552] = 2;
    exp_54_ram[2553] = 250;
    exp_54_ram[2554] = 251;
    exp_54_ram[2555] = 251;
    exp_54_ram[2556] = 250;
    exp_54_ram[2557] = 250;
    exp_54_ram[2558] = 252;
    exp_54_ram[2559] = 252;
    exp_54_ram[2560] = 252;
    exp_54_ram[2561] = 252;
    exp_54_ram[2562] = 250;
    exp_54_ram[2563] = 251;
    exp_54_ram[2564] = 251;
    exp_54_ram[2565] = 251;
    exp_54_ram[2566] = 251;
    exp_54_ram[2567] = 252;
    exp_54_ram[2568] = 252;
    exp_54_ram[2569] = 252;
    exp_54_ram[2570] = 252;
    exp_54_ram[2571] = 246;
    exp_54_ram[2572] = 247;
    exp_54_ram[2573] = 247;
    exp_54_ram[2574] = 246;
    exp_54_ram[2575] = 246;
    exp_54_ram[2576] = 246;
    exp_54_ram[2577] = 246;
    exp_54_ram[2578] = 246;
    exp_54_ram[2579] = 248;
    exp_54_ram[2580] = 246;
    exp_54_ram[2581] = 0;
    exp_54_ram[2582] = 201;
    exp_54_ram[2583] = 252;
    exp_54_ram[2584] = 252;
    exp_54_ram[2585] = 252;
    exp_54_ram[2586] = 2;
    exp_54_ram[2587] = 253;
    exp_54_ram[2588] = 253;
    exp_54_ram[2589] = 255;
    exp_54_ram[2590] = 31;
    exp_54_ram[2591] = 255;
    exp_54_ram[2592] = 0;
    exp_54_ram[2593] = 0;
    exp_54_ram[2594] = 0;
    exp_54_ram[2595] = 0;
    exp_54_ram[2596] = 0;
    exp_54_ram[2597] = 0;
    exp_54_ram[2598] = 252;
    exp_54_ram[2599] = 252;
    exp_54_ram[2600] = 11;
    exp_54_ram[2601] = 252;
    exp_54_ram[2602] = 10;
    exp_54_ram[2603] = 250;
    exp_54_ram[2604] = 251;
    exp_54_ram[2605] = 251;
    exp_54_ram[2606] = 251;
    exp_54_ram[2607] = 251;
    exp_54_ram[2608] = 252;
    exp_54_ram[2609] = 252;
    exp_54_ram[2610] = 252;
    exp_54_ram[2611] = 252;
    exp_54_ram[2612] = 246;
    exp_54_ram[2613] = 247;
    exp_54_ram[2614] = 247;
    exp_54_ram[2615] = 246;
    exp_54_ram[2616] = 246;
    exp_54_ram[2617] = 246;
    exp_54_ram[2618] = 246;
    exp_54_ram[2619] = 246;
    exp_54_ram[2620] = 248;
    exp_54_ram[2621] = 246;
    exp_54_ram[2622] = 0;
    exp_54_ram[2623] = 230;
    exp_54_ram[2624] = 0;
    exp_54_ram[2625] = 0;
    exp_54_ram[2626] = 0;
    exp_54_ram[2627] = 225;
    exp_54_ram[2628] = 0;
    exp_54_ram[2629] = 0;
    exp_54_ram[2630] = 0;
    exp_54_ram[2631] = 0;
    exp_54_ram[2632] = 253;
    exp_54_ram[2633] = 253;
    exp_54_ram[2634] = 64;
    exp_54_ram[2635] = 0;
    exp_54_ram[2636] = 1;
    exp_54_ram[2637] = 64;
    exp_54_ram[2638] = 65;
    exp_54_ram[2639] = 0;
    exp_54_ram[2640] = 252;
    exp_54_ram[2641] = 252;
    exp_54_ram[2642] = 1;
    exp_54_ram[2643] = 253;
    exp_54_ram[2644] = 253;
    exp_54_ram[2645] = 252;
    exp_54_ram[2646] = 252;
    exp_54_ram[2647] = 0;
    exp_54_ram[2648] = 44;
    exp_54_ram[2649] = 0;
    exp_54_ram[2650] = 65;
    exp_54_ram[2651] = 0;
    exp_54_ram[2652] = 253;
    exp_54_ram[2653] = 253;
    exp_54_ram[2654] = 65;
    exp_54_ram[2655] = 0;
    exp_54_ram[2656] = 0;
    exp_54_ram[2657] = 65;
    exp_54_ram[2658] = 64;
    exp_54_ram[2659] = 0;
    exp_54_ram[2660] = 252;
    exp_54_ram[2661] = 252;
    exp_54_ram[2662] = 249;
    exp_54_ram[2663] = 246;
    exp_54_ram[2664] = 253;
    exp_54_ram[2665] = 253;
    exp_54_ram[2666] = 0;
    exp_54_ram[2667] = 114;
    exp_54_ram[2668] = 246;
    exp_54_ram[2669] = 246;
    exp_54_ram[2670] = 246;
    exp_54_ram[2671] = 246;
    exp_54_ram[2672] = 247;
    exp_54_ram[2673] = 247;
    exp_54_ram[2674] = 247;
    exp_54_ram[2675] = 247;
    exp_54_ram[2676] = 248;
    exp_54_ram[2677] = 0;
    exp_54_ram[2678] = 1;
    exp_54_ram[2679] = 1;
    exp_54_ram[2680] = 0;
    exp_54_ram[2681] = 0;
    exp_54_ram[2682] = 0;
    exp_54_ram[2683] = 0;
    exp_54_ram[2684] = 0;
    exp_54_ram[2685] = 2;
    exp_54_ram[2686] = 252;
    exp_54_ram[2687] = 0;
    exp_54_ram[2688] = 249;
    exp_54_ram[2689] = 0;
    exp_54_ram[2690] = 2;
    exp_54_ram[2691] = 7;
    exp_54_ram[2692] = 252;
    exp_54_ram[2693] = 6;
    exp_54_ram[2694] = 250;
    exp_54_ram[2695] = 251;
    exp_54_ram[2696] = 251;
    exp_54_ram[2697] = 251;
    exp_54_ram[2698] = 251;
    exp_54_ram[2699] = 252;
    exp_54_ram[2700] = 252;
    exp_54_ram[2701] = 252;
    exp_54_ram[2702] = 252;
    exp_54_ram[2703] = 246;
    exp_54_ram[2704] = 247;
    exp_54_ram[2705] = 247;
    exp_54_ram[2706] = 246;
    exp_54_ram[2707] = 246;
    exp_54_ram[2708] = 246;
    exp_54_ram[2709] = 246;
    exp_54_ram[2710] = 246;
    exp_54_ram[2711] = 248;
    exp_54_ram[2712] = 246;
    exp_54_ram[2713] = 0;
    exp_54_ram[2714] = 207;
    exp_54_ram[2715] = 0;
    exp_54_ram[2716] = 249;
    exp_54_ram[2717] = 2;
    exp_54_ram[2718] = 0;
    exp_54_ram[2719] = 249;
    exp_54_ram[2720] = 2;
    exp_54_ram[2721] = 253;
    exp_54_ram[2722] = 253;
    exp_54_ram[2723] = 0;
    exp_54_ram[2724] = 0;
    exp_54_ram[2725] = 9;
    exp_54_ram[2726] = 9;
    exp_54_ram[2727] = 9;
    exp_54_ram[2728] = 9;
    exp_54_ram[2729] = 8;
    exp_54_ram[2730] = 10;
    exp_54_ram[2731] = 0;
    exp_54_ram[2732] = 252;
    exp_54_ram[2733] = 2;
    exp_54_ram[2734] = 2;
    exp_54_ram[2735] = 3;
    exp_54_ram[2736] = 3;
    exp_54_ram[2737] = 3;
    exp_54_ram[2738] = 3;
    exp_54_ram[2739] = 3;
    exp_54_ram[2740] = 3;
    exp_54_ram[2741] = 4;
    exp_54_ram[2742] = 252;
    exp_54_ram[2743] = 128;
    exp_54_ram[2744] = 0;
    exp_54_ram[2745] = 0;
    exp_54_ram[2746] = 0;
    exp_54_ram[2747] = 13;
    exp_54_ram[2748] = 0;
    exp_54_ram[2749] = 0;
    exp_54_ram[2750] = 0;
    exp_54_ram[2751] = 0;
    exp_54_ram[2752] = 0;
    exp_54_ram[2753] = 0;
    exp_54_ram[2754] = 216;
    exp_54_ram[2755] = 0;
    exp_54_ram[2756] = 0;
    exp_54_ram[2757] = 252;
    exp_54_ram[2758] = 0;
    exp_54_ram[2759] = 44;
    exp_54_ram[2760] = 44;
    exp_54_ram[2761] = 253;
    exp_54_ram[2762] = 0;
    exp_54_ram[2763] = 252;
    exp_54_ram[2764] = 252;
    exp_54_ram[2765] = 0;
    exp_54_ram[2766] = 253;
    exp_54_ram[2767] = 0;
    exp_54_ram[2768] = 0;
    exp_54_ram[2769] = 252;
    exp_54_ram[2770] = 1;
    exp_54_ram[2771] = 1;
    exp_54_ram[2772] = 253;
    exp_54_ram[2773] = 0;
    exp_54_ram[2774] = 0;
    exp_54_ram[2775] = 0;
    exp_54_ram[2776] = 0;
    exp_54_ram[2777] = 0;
    exp_54_ram[2778] = 0;
    exp_54_ram[2779] = 3;
    exp_54_ram[2780] = 3;
    exp_54_ram[2781] = 3;
    exp_54_ram[2782] = 3;
    exp_54_ram[2783] = 2;
    exp_54_ram[2784] = 2;
    exp_54_ram[2785] = 2;
    exp_54_ram[2786] = 2;
    exp_54_ram[2787] = 4;
    exp_54_ram[2788] = 0;
    exp_54_ram[2789] = 253;
    exp_54_ram[2790] = 2;
    exp_54_ram[2791] = 2;
    exp_54_ram[2792] = 3;
    exp_54_ram[2793] = 3;
    exp_54_ram[2794] = 3;
    exp_54_ram[2795] = 252;
    exp_54_ram[2796] = 252;
    exp_54_ram[2797] = 243;
    exp_54_ram[2798] = 0;
    exp_54_ram[2799] = 0;
    exp_54_ram[2800] = 0;
    exp_54_ram[2801] = 13;
    exp_54_ram[2802] = 0;
    exp_54_ram[2803] = 0;
    exp_54_ram[2804] = 0;
    exp_54_ram[2805] = 0;
    exp_54_ram[2806] = 0;
    exp_54_ram[2807] = 0;
    exp_54_ram[2808] = 202;
    exp_54_ram[2809] = 0;
    exp_54_ram[2810] = 0;
    exp_54_ram[2811] = 254;
    exp_54_ram[2812] = 254;
    exp_54_ram[2813] = 253;
    exp_54_ram[2814] = 253;
    exp_54_ram[2815] = 254;
    exp_54_ram[2816] = 254;
    exp_54_ram[2817] = 64;
    exp_54_ram[2818] = 0;
    exp_54_ram[2819] = 1;
    exp_54_ram[2820] = 64;
    exp_54_ram[2821] = 65;
    exp_54_ram[2822] = 0;
    exp_54_ram[2823] = 0;
    exp_54_ram[2824] = 0;
    exp_54_ram[2825] = 0;
    exp_54_ram[2826] = 44;
    exp_54_ram[2827] = 44;
    exp_54_ram[2828] = 0;
    exp_54_ram[2829] = 2;
    exp_54_ram[2830] = 2;
    exp_54_ram[2831] = 2;
    exp_54_ram[2832] = 2;
    exp_54_ram[2833] = 3;
    exp_54_ram[2834] = 0;
    exp_54_ram[2835] = 249;
    exp_54_ram[2836] = 6;
    exp_54_ram[2837] = 6;
    exp_54_ram[2838] = 7;
    exp_54_ram[2839] = 248;
    exp_54_ram[2840] = 0;
    exp_54_ram[2841] = 138;
    exp_54_ram[2842] = 0;
    exp_54_ram[2843] = 0;
    exp_54_ram[2844] = 0;
    exp_54_ram[2845] = 0;
    exp_54_ram[2846] = 1;
    exp_54_ram[2847] = 252;
    exp_54_ram[2848] = 252;
    exp_54_ram[2849] = 252;
    exp_54_ram[2850] = 254;
    exp_54_ram[2851] = 254;
    exp_54_ram[2852] = 1;
    exp_54_ram[2853] = 254;
    exp_54_ram[2854] = 0;
    exp_54_ram[2855] = 140;
    exp_54_ram[2856] = 0;
    exp_54_ram[2857] = 0;
    exp_54_ram[2858] = 0;
    exp_54_ram[2859] = 0;
    exp_54_ram[2860] = 1;
    exp_54_ram[2861] = 1;
    exp_54_ram[2862] = 1;
    exp_54_ram[2863] = 1;
    exp_54_ram[2864] = 2;
    exp_54_ram[2865] = 251;
    exp_54_ram[2866] = 250;
    exp_54_ram[2867] = 251;
    exp_54_ram[2868] = 251;
    exp_54_ram[2869] = 250;
    exp_54_ram[2870] = 252;
    exp_54_ram[2871] = 252;
    exp_54_ram[2872] = 252;
    exp_54_ram[2873] = 252;
    exp_54_ram[2874] = 2;
    exp_54_ram[2875] = 252;
    exp_54_ram[2876] = 254;
    exp_54_ram[2877] = 4;
    exp_54_ram[2878] = 249;
    exp_54_ram[2879] = 1;
    exp_54_ram[2880] = 0;
    exp_54_ram[2881] = 0;
    exp_54_ram[2882] = 0;
    exp_54_ram[2883] = 254;
    exp_54_ram[2884] = 0;
    exp_54_ram[2885] = 255;
    exp_54_ram[2886] = 0;
    exp_54_ram[2887] = 254;
    exp_54_ram[2888] = 0;
    exp_54_ram[2889] = 45;
    exp_54_ram[2890] = 254;
    exp_54_ram[2891] = 0;
    exp_54_ram[2892] = 0;
    exp_54_ram[2893] = 254;
    exp_54_ram[2894] = 0;
    exp_54_ram[2895] = 254;
    exp_54_ram[2896] = 254;
    exp_54_ram[2897] = 0;
    exp_54_ram[2898] = 250;
    exp_54_ram[2899] = 0;
    exp_54_ram[2900] = 45;
    exp_54_ram[2901] = 2;
    exp_54_ram[2902] = 0;
    exp_54_ram[2903] = 254;
    exp_54_ram[2904] = 5;
    exp_54_ram[2905] = 249;
    exp_54_ram[2906] = 1;
    exp_54_ram[2907] = 0;
    exp_54_ram[2908] = 0;
    exp_54_ram[2909] = 0;
    exp_54_ram[2910] = 254;
    exp_54_ram[2911] = 0;
    exp_54_ram[2912] = 254;
    exp_54_ram[2913] = 0;
    exp_54_ram[2914] = 255;
    exp_54_ram[2915] = 0;
    exp_54_ram[2916] = 251;
    exp_54_ram[2917] = 0;
    exp_54_ram[2918] = 45;
    exp_54_ram[2919] = 0;
    exp_54_ram[2920] = 0;
    exp_54_ram[2921] = 254;
    exp_54_ram[2922] = 0;
    exp_54_ram[2923] = 254;
    exp_54_ram[2924] = 254;
    exp_54_ram[2925] = 0;
    exp_54_ram[2926] = 250;
    exp_54_ram[2927] = 0;
    exp_54_ram[2928] = 45;
    exp_54_ram[2929] = 2;
    exp_54_ram[2930] = 0;
    exp_54_ram[2931] = 249;
    exp_54_ram[2932] = 0;
    exp_54_ram[2933] = 0;
    exp_54_ram[2934] = 0;
    exp_54_ram[2935] = 43;
    exp_54_ram[2936] = 0;
    exp_54_ram[2937] = 0;
    exp_54_ram[2938] = 250;
    exp_54_ram[2939] = 250;
    exp_54_ram[2940] = 250;
    exp_54_ram[2941] = 15;
    exp_54_ram[2942] = 3;
    exp_54_ram[2943] = 15;
    exp_54_ram[2944] = 0;
    exp_54_ram[2945] = 45;
    exp_54_ram[2946] = 0;
    exp_54_ram[2947] = 250;
    exp_54_ram[2948] = 15;
    exp_54_ram[2949] = 3;
    exp_54_ram[2950] = 15;
    exp_54_ram[2951] = 0;
    exp_54_ram[2952] = 45;
    exp_54_ram[2953] = 0;
    exp_54_ram[2954] = 0;
    exp_54_ram[2955] = 45;
    exp_54_ram[2956] = 2;
    exp_54_ram[2957] = 0;
    exp_54_ram[2958] = 249;
    exp_54_ram[2959] = 0;
    exp_54_ram[2960] = 0;
    exp_54_ram[2961] = 0;
    exp_54_ram[2962] = 36;
    exp_54_ram[2963] = 0;
    exp_54_ram[2964] = 0;
    exp_54_ram[2965] = 250;
    exp_54_ram[2966] = 250;
    exp_54_ram[2967] = 250;
    exp_54_ram[2968] = 15;
    exp_54_ram[2969] = 3;
    exp_54_ram[2970] = 15;
    exp_54_ram[2971] = 0;
    exp_54_ram[2972] = 45;
    exp_54_ram[2973] = 0;
    exp_54_ram[2974] = 250;
    exp_54_ram[2975] = 15;
    exp_54_ram[2976] = 3;
    exp_54_ram[2977] = 15;
    exp_54_ram[2978] = 0;
    exp_54_ram[2979] = 45;
    exp_54_ram[2980] = 0;
    exp_54_ram[2981] = 0;
    exp_54_ram[2982] = 45;
    exp_54_ram[2983] = 3;
    exp_54_ram[2984] = 0;
    exp_54_ram[2985] = 249;
    exp_54_ram[2986] = 0;
    exp_54_ram[2987] = 0;
    exp_54_ram[2988] = 0;
    exp_54_ram[2989] = 30;
    exp_54_ram[2990] = 0;
    exp_54_ram[2991] = 0;
    exp_54_ram[2992] = 250;
    exp_54_ram[2993] = 250;
    exp_54_ram[2994] = 250;
    exp_54_ram[2995] = 15;
    exp_54_ram[2996] = 3;
    exp_54_ram[2997] = 15;
    exp_54_ram[2998] = 0;
    exp_54_ram[2999] = 45;
    exp_54_ram[3000] = 0;
    exp_54_ram[3001] = 250;
    exp_54_ram[3002] = 15;
    exp_54_ram[3003] = 3;
    exp_54_ram[3004] = 15;
    exp_54_ram[3005] = 0;
    exp_54_ram[3006] = 45;
    exp_54_ram[3007] = 0;
    exp_54_ram[3008] = 0;
    exp_54_ram[3009] = 45;
    exp_54_ram[3010] = 3;
    exp_54_ram[3011] = 0;
    exp_54_ram[3012] = 249;
    exp_54_ram[3013] = 0;
    exp_54_ram[3014] = 0;
    exp_54_ram[3015] = 0;
    exp_54_ram[3016] = 23;
    exp_54_ram[3017] = 0;
    exp_54_ram[3018] = 0;
    exp_54_ram[3019] = 250;
    exp_54_ram[3020] = 250;
    exp_54_ram[3021] = 250;
    exp_54_ram[3022] = 15;
    exp_54_ram[3023] = 3;
    exp_54_ram[3024] = 15;
    exp_54_ram[3025] = 0;
    exp_54_ram[3026] = 45;
    exp_54_ram[3027] = 0;
    exp_54_ram[3028] = 250;
    exp_54_ram[3029] = 15;
    exp_54_ram[3030] = 3;
    exp_54_ram[3031] = 15;
    exp_54_ram[3032] = 0;
    exp_54_ram[3033] = 45;
    exp_54_ram[3034] = 0;
    exp_54_ram[3035] = 0;
    exp_54_ram[3036] = 45;
    exp_54_ram[3037] = 2;
    exp_54_ram[3038] = 0;
    exp_54_ram[3039] = 249;
    exp_54_ram[3040] = 1;
    exp_54_ram[3041] = 118;
    exp_54_ram[3042] = 62;
    exp_54_ram[3043] = 0;
    exp_54_ram[3044] = 16;
    exp_54_ram[3045] = 0;
    exp_54_ram[3046] = 0;
    exp_54_ram[3047] = 250;
    exp_54_ram[3048] = 250;
    exp_54_ram[3049] = 250;
    exp_54_ram[3050] = 15;
    exp_54_ram[3051] = 3;
    exp_54_ram[3052] = 15;
    exp_54_ram[3053] = 0;
    exp_54_ram[3054] = 45;
    exp_54_ram[3055] = 0;
    exp_54_ram[3056] = 250;
    exp_54_ram[3057] = 6;
    exp_54_ram[3058] = 0;
    exp_54_ram[3059] = 12;
    exp_54_ram[3060] = 0;
    exp_54_ram[3061] = 0;
    exp_54_ram[3062] = 250;
    exp_54_ram[3063] = 250;
    exp_54_ram[3064] = 250;
    exp_54_ram[3065] = 15;
    exp_54_ram[3066] = 3;
    exp_54_ram[3067] = 15;
    exp_54_ram[3068] = 0;
    exp_54_ram[3069] = 45;
    exp_54_ram[3070] = 0;
    exp_54_ram[3071] = 250;
    exp_54_ram[3072] = 0;
    exp_54_ram[3073] = 0;
    exp_54_ram[3074] = 8;
    exp_54_ram[3075] = 0;
    exp_54_ram[3076] = 0;
    exp_54_ram[3077] = 250;
    exp_54_ram[3078] = 250;
    exp_54_ram[3079] = 250;
    exp_54_ram[3080] = 15;
    exp_54_ram[3081] = 3;
    exp_54_ram[3082] = 15;
    exp_54_ram[3083] = 0;
    exp_54_ram[3084] = 45;
    exp_54_ram[3085] = 0;
    exp_54_ram[3086] = 250;
    exp_54_ram[3087] = 15;
    exp_54_ram[3088] = 3;
    exp_54_ram[3089] = 15;
    exp_54_ram[3090] = 0;
    exp_54_ram[3091] = 45;
    exp_54_ram[3092] = 0;
    exp_54_ram[3093] = 0;
    exp_54_ram[3094] = 45;
    exp_54_ram[3095] = 0;
    exp_54_ram[3096] = 0;
    exp_54_ram[3097] = 0;
    exp_54_ram[3098] = 45;
    exp_54_ram[3099] = 0;
    exp_54_ram[3100] = 0;
    exp_54_ram[3101] = 45;
    exp_54_ram[3102] = 0;
    exp_54_ram[3103] = 6;
    exp_54_ram[3104] = 6;
    exp_54_ram[3105] = 7;
    exp_54_ram[3106] = 0;
    exp_54_ram[3107] = 254;
    exp_54_ram[3108] = 0;
    exp_54_ram[3109] = 0;
    exp_54_ram[3110] = 2;
    exp_54_ram[3111] = 254;
    exp_54_ram[3112] = 254;
    exp_54_ram[3113] = 55;
    exp_54_ram[3114] = 0;
    exp_54_ram[3115] = 0;
    exp_54_ram[3116] = 185;
    exp_54_ram[3117] = 0;
    exp_54_ram[3118] = 0;
    exp_54_ram[3119] = 1;
    exp_54_ram[3120] = 1;
    exp_54_ram[3121] = 2;
    exp_54_ram[3122] = 0;
    exp_54_ram[3123] = 248;
    exp_54_ram[3124] = 6;
    exp_54_ram[3125] = 6;
    exp_54_ram[3126] = 7;
    exp_54_ram[3127] = 7;
    exp_54_ram[3128] = 7;
    exp_54_ram[3129] = 7;
    exp_54_ram[3130] = 7;
    exp_54_ram[3131] = 7;
    exp_54_ram[3132] = 5;
    exp_54_ram[3133] = 5;
    exp_54_ram[3134] = 8;
    exp_54_ram[3135] = 248;
    exp_54_ram[3136] = 248;
    exp_54_ram[3137] = 248;
    exp_54_ram[3138] = 123;
    exp_54_ram[3139] = 250;
    exp_54_ram[3140] = 0;
    exp_54_ram[3141] = 250;
    exp_54_ram[3142] = 251;
    exp_54_ram[3143] = 0;
    exp_54_ram[3144] = 175;
    exp_54_ram[3145] = 252;
    exp_54_ram[3146] = 252;
    exp_54_ram[3147] = 0;
    exp_54_ram[3148] = 24;
    exp_54_ram[3149] = 2;
    exp_54_ram[3150] = 252;
    exp_54_ram[3151] = 252;
    exp_54_ram[3152] = 0;
    exp_54_ram[3153] = 0;
    exp_54_ram[3154] = 248;
    exp_54_ram[3155] = 0;
    exp_54_ram[3156] = 6;
    exp_54_ram[3157] = 248;
    exp_54_ram[3158] = 0;
    exp_54_ram[3159] = 0;
    exp_54_ram[3160] = 248;
    exp_54_ram[3161] = 0;
    exp_54_ram[3162] = 4;
    exp_54_ram[3163] = 251;
    exp_54_ram[3164] = 0;
    exp_54_ram[3165] = 250;
    exp_54_ram[3166] = 251;
    exp_54_ram[3167] = 0;
    exp_54_ram[3168] = 252;
    exp_54_ram[3169] = 0;
    exp_54_ram[3170] = 250;
    exp_54_ram[3171] = 252;
    exp_54_ram[3172] = 0;
    exp_54_ram[3173] = 0;
    exp_54_ram[3174] = 248;
    exp_54_ram[3175] = 248;
    exp_54_ram[3176] = 65;
    exp_54_ram[3177] = 0;
    exp_54_ram[3178] = 0;
    exp_54_ram[3179] = 65;
    exp_54_ram[3180] = 64;
    exp_54_ram[3181] = 0;
    exp_54_ram[3182] = 248;
    exp_54_ram[3183] = 248;
    exp_54_ram[3184] = 245;
    exp_54_ram[3185] = 0;
    exp_54_ram[3186] = 250;
    exp_54_ram[3187] = 252;
    exp_54_ram[3188] = 251;
    exp_54_ram[3189] = 0;
    exp_54_ram[3190] = 251;
    exp_54_ram[3191] = 0;
    exp_54_ram[3192] = 0;
    exp_54_ram[3193] = 167;
    exp_54_ram[3194] = 252;
    exp_54_ram[3195] = 252;
    exp_54_ram[3196] = 0;
    exp_54_ram[3197] = 24;
    exp_54_ram[3198] = 2;
    exp_54_ram[3199] = 252;
    exp_54_ram[3200] = 252;
    exp_54_ram[3201] = 0;
    exp_54_ram[3202] = 0;
    exp_54_ram[3203] = 248;
    exp_54_ram[3204] = 0;
    exp_54_ram[3205] = 8;
    exp_54_ram[3206] = 248;
    exp_54_ram[3207] = 0;
    exp_54_ram[3208] = 0;
    exp_54_ram[3209] = 248;
    exp_54_ram[3210] = 0;
    exp_54_ram[3211] = 6;
    exp_54_ram[3212] = 251;
    exp_54_ram[3213] = 0;
    exp_54_ram[3214] = 250;
    exp_54_ram[3215] = 251;
    exp_54_ram[3216] = 0;
    exp_54_ram[3217] = 252;
    exp_54_ram[3218] = 0;
    exp_54_ram[3219] = 250;
    exp_54_ram[3220] = 252;
    exp_54_ram[3221] = 0;
    exp_54_ram[3222] = 252;
    exp_54_ram[3223] = 0;
    exp_54_ram[3224] = 252;
    exp_54_ram[3225] = 252;
    exp_54_ram[3226] = 0;
    exp_54_ram[3227] = 0;
    exp_54_ram[3228] = 248;
    exp_54_ram[3229] = 248;
    exp_54_ram[3230] = 65;
    exp_54_ram[3231] = 0;
    exp_54_ram[3232] = 0;
    exp_54_ram[3233] = 65;
    exp_54_ram[3234] = 64;
    exp_54_ram[3235] = 0;
    exp_54_ram[3236] = 248;
    exp_54_ram[3237] = 248;
    exp_54_ram[3238] = 243;
    exp_54_ram[3239] = 0;
    exp_54_ram[3240] = 251;
    exp_54_ram[3241] = 137;
    exp_54_ram[3242] = 250;
    exp_54_ram[3243] = 248;
    exp_54_ram[3244] = 0;
    exp_54_ram[3245] = 24;
    exp_54_ram[3246] = 0;
    exp_54_ram[3247] = 93;
    exp_54_ram[3248] = 0;
    exp_54_ram[3249] = 0;
    exp_54_ram[3250] = 248;
    exp_54_ram[3251] = 250;
    exp_54_ram[3252] = 249;
    exp_54_ram[3253] = 0;
    exp_54_ram[3254] = 250;
    exp_54_ram[3255] = 251;
    exp_54_ram[3256] = 249;
    exp_54_ram[3257] = 0;
    exp_54_ram[3258] = 250;
    exp_54_ram[3259] = 251;
    exp_54_ram[3260] = 0;
    exp_54_ram[3261] = 2;
    exp_54_ram[3262] = 250;
    exp_54_ram[3263] = 252;
    exp_54_ram[3264] = 249;
    exp_54_ram[3265] = 0;
    exp_54_ram[3266] = 252;
    exp_54_ram[3267] = 250;
    exp_54_ram[3268] = 248;
    exp_54_ram[3269] = 65;
    exp_54_ram[3270] = 248;
    exp_54_ram[3271] = 248;
    exp_54_ram[3272] = 0;
    exp_54_ram[3273] = 225;
    exp_54_ram[3274] = 0;
    exp_54_ram[3275] = 86;
    exp_54_ram[3276] = 0;
    exp_54_ram[3277] = 0;
    exp_54_ram[3278] = 248;
    exp_54_ram[3279] = 250;
    exp_54_ram[3280] = 249;
    exp_54_ram[3281] = 250;
    exp_54_ram[3282] = 250;
    exp_54_ram[3283] = 248;
    exp_54_ram[3284] = 65;
    exp_54_ram[3285] = 248;
    exp_54_ram[3286] = 248;
    exp_54_ram[3287] = 3;
    exp_54_ram[3288] = 0;
    exp_54_ram[3289] = 83;
    exp_54_ram[3290] = 0;
    exp_54_ram[3291] = 0;
    exp_54_ram[3292] = 248;
    exp_54_ram[3293] = 250;
    exp_54_ram[3294] = 249;
    exp_54_ram[3295] = 250;
    exp_54_ram[3296] = 250;
    exp_54_ram[3297] = 248;
    exp_54_ram[3298] = 65;
    exp_54_ram[3299] = 248;
    exp_54_ram[3300] = 248;
    exp_54_ram[3301] = 250;
    exp_54_ram[3302] = 248;
    exp_54_ram[3303] = 250;
    exp_54_ram[3304] = 250;
    exp_54_ram[3305] = 250;
    exp_54_ram[3306] = 251;
    exp_54_ram[3307] = 251;
    exp_54_ram[3308] = 251;
    exp_54_ram[3309] = 251;
    exp_54_ram[3310] = 252;
    exp_54_ram[3311] = 252;
    exp_54_ram[3312] = 1;
    exp_54_ram[3313] = 0;
    exp_54_ram[3314] = 1;
    exp_54_ram[3315] = 1;
    exp_54_ram[3316] = 0;
    exp_54_ram[3317] = 0;
    exp_54_ram[3318] = 0;
    exp_54_ram[3319] = 0;
    exp_54_ram[3320] = 2;
    exp_54_ram[3321] = 248;
    exp_54_ram[3322] = 7;
    exp_54_ram[3323] = 7;
    exp_54_ram[3324] = 7;
    exp_54_ram[3325] = 7;
    exp_54_ram[3326] = 6;
    exp_54_ram[3327] = 6;
    exp_54_ram[3328] = 6;
    exp_54_ram[3329] = 6;
    exp_54_ram[3330] = 5;
    exp_54_ram[3331] = 5;
    exp_54_ram[3332] = 8;
    exp_54_ram[3333] = 0;
    exp_54_ram[3334] = 246;
    exp_54_ram[3335] = 8;
    exp_54_ram[3336] = 8;
    exp_54_ram[3337] = 8;
    exp_54_ram[3338] = 9;
    exp_54_ram[3339] = 9;
    exp_54_ram[3340] = 10;
    exp_54_ram[3341] = 248;
    exp_54_ram[3342] = 0;
    exp_54_ram[3343] = 0;
    exp_54_ram[3344] = 252;
    exp_54_ram[3345] = 253;
    exp_54_ram[3346] = 249;
    exp_54_ram[3347] = 0;
    exp_54_ram[3348] = 0;
    exp_54_ram[3349] = 252;
    exp_54_ram[3350] = 252;
    exp_54_ram[3351] = 253;
    exp_54_ram[3352] = 253;
    exp_54_ram[3353] = 222;
    exp_54_ram[3354] = 0;
    exp_54_ram[3355] = 0;
    exp_54_ram[3356] = 0;
    exp_54_ram[3357] = 225;
    exp_54_ram[3358] = 0;
    exp_54_ram[3359] = 252;
    exp_54_ram[3360] = 252;
    exp_54_ram[3361] = 0;
    exp_54_ram[3362] = 44;
    exp_54_ram[3363] = 0;
    exp_54_ram[3364] = 65;
    exp_54_ram[3365] = 0;
    exp_54_ram[3366] = 253;
    exp_54_ram[3367] = 253;
    exp_54_ram[3368] = 0;
    exp_54_ram[3369] = 0;
    exp_54_ram[3370] = 1;
    exp_54_ram[3371] = 0;
    exp_54_ram[3372] = 0;
    exp_54_ram[3373] = 0;
    exp_54_ram[3374] = 0;
    exp_54_ram[3375] = 0;
    exp_54_ram[3376] = 253;
    exp_54_ram[3377] = 253;
    exp_54_ram[3378] = 0;
    exp_54_ram[3379] = 0;
    exp_54_ram[3380] = 0;
    exp_54_ram[3381] = 0;
    exp_54_ram[3382] = 0;
    exp_54_ram[3383] = 0;
    exp_54_ram[3384] = 252;
    exp_54_ram[3385] = 252;
    exp_54_ram[3386] = 0;
    exp_54_ram[3387] = 46;
    exp_54_ram[3388] = 246;
    exp_54_ram[3389] = 252;
    exp_54_ram[3390] = 252;
    exp_54_ram[3391] = 0;
    exp_54_ram[3392] = 188;
    exp_54_ram[3393] = 246;
    exp_54_ram[3394] = 246;
    exp_54_ram[3395] = 246;
    exp_54_ram[3396] = 246;
    exp_54_ram[3397] = 247;
    exp_54_ram[3398] = 247;
    exp_54_ram[3399] = 247;
    exp_54_ram[3400] = 247;
    exp_54_ram[3401] = 248;
    exp_54_ram[3402] = 0;
    exp_54_ram[3403] = 1;
    exp_54_ram[3404] = 1;
    exp_54_ram[3405] = 0;
    exp_54_ram[3406] = 0;
    exp_54_ram[3407] = 0;
    exp_54_ram[3408] = 0;
    exp_54_ram[3409] = 0;
    exp_54_ram[3410] = 2;
    exp_54_ram[3411] = 253;
    exp_54_ram[3412] = 253;
    exp_54_ram[3413] = 207;
    exp_54_ram[3414] = 0;
    exp_54_ram[3415] = 0;
    exp_54_ram[3416] = 46;
    exp_54_ram[3417] = 2;
    exp_54_ram[3418] = 0;
    exp_54_ram[3419] = 46;
    exp_54_ram[3420] = 0;
    exp_54_ram[3421] = 9;
    exp_54_ram[3422] = 9;
    exp_54_ram[3423] = 9;
    exp_54_ram[3424] = 9;
    exp_54_ram[3425] = 8;
    exp_54_ram[3426] = 10;
    exp_54_ram[3427] = 0;
    exp_54_ram[3428] = 253;
    exp_54_ram[3429] = 2;
    exp_54_ram[3430] = 2;
    exp_54_ram[3431] = 3;
    exp_54_ram[3432] = 252;
    exp_54_ram[3433] = 254;
    exp_54_ram[3434] = 253;
    exp_54_ram[3435] = 218;
    exp_54_ram[3436] = 0;
    exp_54_ram[3437] = 254;
    exp_54_ram[3438] = 254;
    exp_54_ram[3439] = 253;
    exp_54_ram[3440] = 0;
    exp_54_ram[3441] = 2;
    exp_54_ram[3442] = 254;
    exp_54_ram[3443] = 0;
    exp_54_ram[3444] = 0;
    exp_54_ram[3445] = 0;
    exp_54_ram[3446] = 0;
    exp_54_ram[3447] = 254;
    exp_54_ram[3448] = 254;
    exp_54_ram[3449] = 254;
    exp_54_ram[3450] = 0;
    exp_54_ram[3451] = 253;
    exp_54_ram[3452] = 254;
    exp_54_ram[3453] = 251;
    exp_54_ram[3454] = 0;
    exp_54_ram[3455] = 254;
    exp_54_ram[3456] = 0;
    exp_54_ram[3457] = 2;
    exp_54_ram[3458] = 2;
    exp_54_ram[3459] = 3;
    exp_54_ram[3460] = 0;
    exp_54_ram[3461] = 255;
    exp_54_ram[3462] = 0;
    exp_54_ram[3463] = 0;
    exp_54_ram[3464] = 1;
    exp_54_ram[3465] = 0;
    exp_54_ram[3466] = 13;
    exp_54_ram[3467] = 0;
    exp_54_ram[3468] = 246;
    exp_54_ram[3469] = 0;
    exp_54_ram[3470] = 0;
    exp_54_ram[3471] = 0;
    exp_54_ram[3472] = 0;
    exp_54_ram[3473] = 1;
    exp_54_ram[3474] = 0;
    exp_54_ram[3475] = 253;
    exp_54_ram[3476] = 2;
    exp_54_ram[3477] = 2;
    exp_54_ram[3478] = 3;
    exp_54_ram[3479] = 3;
    exp_54_ram[3480] = 3;
    exp_54_ram[3481] = 252;
    exp_54_ram[3482] = 199;
    exp_54_ram[3483] = 254;
    exp_54_ram[3484] = 254;
    exp_54_ram[3485] = 0;
    exp_54_ram[3486] = 198;
    exp_54_ram[3487] = 0;
    exp_54_ram[3488] = 0;
    exp_54_ram[3489] = 254;
    exp_54_ram[3490] = 254;
    exp_54_ram[3491] = 64;
    exp_54_ram[3492] = 0;
    exp_54_ram[3493] = 1;
    exp_54_ram[3494] = 64;
    exp_54_ram[3495] = 65;
    exp_54_ram[3496] = 0;
    exp_54_ram[3497] = 253;
    exp_54_ram[3498] = 0;
    exp_54_ram[3499] = 0;
    exp_54_ram[3500] = 0;
    exp_54_ram[3501] = 0;
    exp_54_ram[3502] = 252;
    exp_54_ram[3503] = 0;
    exp_54_ram[3504] = 0;
    exp_54_ram[3505] = 0;
    exp_54_ram[3506] = 0;
    exp_54_ram[3507] = 0;
    exp_54_ram[3508] = 250;
    exp_54_ram[3509] = 0;
    exp_54_ram[3510] = 0;
    exp_54_ram[3511] = 2;
    exp_54_ram[3512] = 2;
    exp_54_ram[3513] = 2;
    exp_54_ram[3514] = 2;
    exp_54_ram[3515] = 3;
    exp_54_ram[3516] = 0;
    exp_54_ram[3517] = 255;
    exp_54_ram[3518] = 0;
    exp_54_ram[3519] = 0;
    exp_54_ram[3520] = 1;
    exp_54_ram[3521] = 0;
    exp_54_ram[3522] = 142;
    exp_54_ram[3523] = 248;
    exp_54_ram[3524] = 0;
    exp_54_ram[3525] = 0;
    exp_54_ram[3526] = 0;
    exp_54_ram[3527] = 1;
    exp_54_ram[3528] = 0;
    exp_54_ram[3529] = 254;
    exp_54_ram[3530] = 0;
    exp_54_ram[3531] = 0;
    exp_54_ram[3532] = 2;
    exp_54_ram[3533] = 0;
    exp_54_ram[3534] = 143;
    exp_54_ram[3535] = 245;
    exp_54_ram[3536] = 0;
    exp_54_ram[3537] = 254;
    exp_54_ram[3538] = 254;
    exp_54_ram[3539] = 11;
    exp_54_ram[3540] = 254;
    exp_54_ram[3541] = 0;
    exp_54_ram[3542] = 145;
    exp_54_ram[3543] = 243;
    exp_54_ram[3544] = 3;
    exp_54_ram[3545] = 254;
    exp_54_ram[3546] = 0;
    exp_54_ram[3547] = 254;
    exp_54_ram[3548] = 0;
    exp_54_ram[3549] = 13;
    exp_54_ram[3550] = 0;
    exp_54_ram[3551] = 254;
    exp_54_ram[3552] = 192;
    exp_54_ram[3553] = 0;
    exp_54_ram[3554] = 13;
    exp_54_ram[3555] = 0;
    exp_54_ram[3556] = 2;
    exp_54_ram[3557] = 0;
    exp_54_ram[3558] = 235;
    exp_54_ram[3559] = 254;
    exp_54_ram[3560] = 7;
    exp_54_ram[3561] = 252;
    exp_54_ram[3562] = 3;
    exp_54_ram[3563] = 254;
    exp_54_ram[3564] = 64;
    exp_54_ram[3565] = 254;
    exp_54_ram[3566] = 0;
    exp_54_ram[3567] = 13;
    exp_54_ram[3568] = 0;
    exp_54_ram[3569] = 254;
    exp_54_ram[3570] = 187;
    exp_54_ram[3571] = 0;
    exp_54_ram[3572] = 13;
    exp_54_ram[3573] = 0;
    exp_54_ram[3574] = 2;
    exp_54_ram[3575] = 0;
    exp_54_ram[3576] = 230;
    exp_54_ram[3577] = 254;
    exp_54_ram[3578] = 0;
    exp_54_ram[3579] = 252;
    exp_54_ram[3580] = 254;
    exp_54_ram[3581] = 0;
    exp_54_ram[3582] = 254;
    exp_54_ram[3583] = 254;
    exp_54_ram[3584] = 0;
    exp_54_ram[3585] = 244;
    exp_54_ram[3586] = 0;
    exp_54_ram[3587] = 13;
    exp_54_ram[3588] = 0;
    exp_54_ram[3589] = 0;
    exp_54_ram[3590] = 182;
    exp_54_ram[3591] = 0;
    exp_54_ram[3592] = 1;
    exp_54_ram[3593] = 1;
    exp_54_ram[3594] = 2;
    exp_54_ram[3595] = 0;
    exp_54_ram[3596] = 249;
    exp_54_ram[3597] = 6;
    exp_54_ram[3598] = 6;
    exp_54_ram[3599] = 7;
    exp_54_ram[3600] = 7;
    exp_54_ram[3601] = 5;
    exp_54_ram[3602] = 5;
    exp_54_ram[3603] = 5;
    exp_54_ram[3604] = 5;
    exp_54_ram[3605] = 5;
    exp_54_ram[3606] = 5;
    exp_54_ram[3607] = 5;
    exp_54_ram[3608] = 5;
    exp_54_ram[3609] = 7;
    exp_54_ram[3610] = 0;
    exp_54_ram[3611] = 250;
    exp_54_ram[3612] = 0;
    exp_54_ram[3613] = 0;
    exp_54_ram[3614] = 250;
    exp_54_ram[3615] = 250;
    exp_54_ram[3616] = 166;
    exp_54_ram[3617] = 252;
    exp_54_ram[3618] = 252;
    exp_54_ram[3619] = 252;
    exp_54_ram[3620] = 6;
    exp_54_ram[3621] = 251;
    exp_54_ram[3622] = 18;
    exp_54_ram[3623] = 103;
    exp_54_ram[3624] = 2;
    exp_54_ram[3625] = 250;
    exp_54_ram[3626] = 251;
    exp_54_ram[3627] = 18;
    exp_54_ram[3628] = 103;
    exp_54_ram[3629] = 2;
    exp_54_ram[3630] = 250;
    exp_54_ram[3631] = 251;
    exp_54_ram[3632] = 18;
    exp_54_ram[3633] = 103;
    exp_54_ram[3634] = 2;
    exp_54_ram[3635] = 250;
    exp_54_ram[3636] = 251;
    exp_54_ram[3637] = 18;
    exp_54_ram[3638] = 103;
    exp_54_ram[3639] = 2;
    exp_54_ram[3640] = 250;
    exp_54_ram[3641] = 252;
    exp_54_ram[3642] = 0;
    exp_54_ram[3643] = 252;
    exp_54_ram[3644] = 159;
    exp_54_ram[3645] = 0;
    exp_54_ram[3646] = 0;
    exp_54_ram[3647] = 252;
    exp_54_ram[3648] = 252;
    exp_54_ram[3649] = 64;
    exp_54_ram[3650] = 0;
    exp_54_ram[3651] = 1;
    exp_54_ram[3652] = 64;
    exp_54_ram[3653] = 65;
    exp_54_ram[3654] = 0;
    exp_54_ram[3655] = 0;
    exp_54_ram[3656] = 13;
    exp_54_ram[3657] = 250;
    exp_54_ram[3658] = 250;
    exp_54_ram[3659] = 250;
    exp_54_ram[3660] = 250;
    exp_54_ram[3661] = 0;
    exp_54_ram[3662] = 0;
    exp_54_ram[3663] = 244;
    exp_54_ram[3664] = 0;
    exp_54_ram[3665] = 0;
    exp_54_ram[3666] = 0;
    exp_54_ram[3667] = 0;
    exp_54_ram[3668] = 0;
    exp_54_ram[3669] = 244;
    exp_54_ram[3670] = 252;
    exp_54_ram[3671] = 0;
    exp_54_ram[3672] = 145;
    exp_54_ram[3673] = 211;
    exp_54_ram[3674] = 151;
    exp_54_ram[3675] = 252;
    exp_54_ram[3676] = 252;
    exp_54_ram[3677] = 252;
    exp_54_ram[3678] = 18;
    exp_54_ram[3679] = 251;
    exp_54_ram[3680] = 251;
    exp_54_ram[3681] = 18;
    exp_54_ram[3682] = 103;
    exp_54_ram[3683] = 2;
    exp_54_ram[3684] = 0;
    exp_54_ram[3685] = 2;
    exp_54_ram[3686] = 0;
    exp_54_ram[3687] = 18;
    exp_54_ram[3688] = 103;
    exp_54_ram[3689] = 2;
    exp_54_ram[3690] = 2;
    exp_54_ram[3691] = 0;
    exp_54_ram[3692] = 1;
    exp_54_ram[3693] = 0;
    exp_54_ram[3694] = 251;
    exp_54_ram[3695] = 251;
    exp_54_ram[3696] = 251;
    exp_54_ram[3697] = 251;
    exp_54_ram[3698] = 18;
    exp_54_ram[3699] = 103;
    exp_54_ram[3700] = 2;
    exp_54_ram[3701] = 0;
    exp_54_ram[3702] = 2;
    exp_54_ram[3703] = 0;
    exp_54_ram[3704] = 18;
    exp_54_ram[3705] = 103;
    exp_54_ram[3706] = 2;
    exp_54_ram[3707] = 2;
    exp_54_ram[3708] = 0;
    exp_54_ram[3709] = 1;
    exp_54_ram[3710] = 0;
    exp_54_ram[3711] = 251;
    exp_54_ram[3712] = 251;
    exp_54_ram[3713] = 251;
    exp_54_ram[3714] = 251;
    exp_54_ram[3715] = 18;
    exp_54_ram[3716] = 103;
    exp_54_ram[3717] = 2;
    exp_54_ram[3718] = 0;
    exp_54_ram[3719] = 2;
    exp_54_ram[3720] = 0;
    exp_54_ram[3721] = 18;
    exp_54_ram[3722] = 103;
    exp_54_ram[3723] = 2;
    exp_54_ram[3724] = 2;
    exp_54_ram[3725] = 0;
    exp_54_ram[3726] = 1;
    exp_54_ram[3727] = 0;
    exp_54_ram[3728] = 251;
    exp_54_ram[3729] = 251;
    exp_54_ram[3730] = 251;
    exp_54_ram[3731] = 251;
    exp_54_ram[3732] = 18;
    exp_54_ram[3733] = 103;
    exp_54_ram[3734] = 2;
    exp_54_ram[3735] = 0;
    exp_54_ram[3736] = 2;
    exp_54_ram[3737] = 0;
    exp_54_ram[3738] = 18;
    exp_54_ram[3739] = 103;
    exp_54_ram[3740] = 2;
    exp_54_ram[3741] = 2;
    exp_54_ram[3742] = 0;
    exp_54_ram[3743] = 1;
    exp_54_ram[3744] = 0;
    exp_54_ram[3745] = 251;
    exp_54_ram[3746] = 251;
    exp_54_ram[3747] = 252;
    exp_54_ram[3748] = 0;
    exp_54_ram[3749] = 252;
    exp_54_ram[3750] = 132;
    exp_54_ram[3751] = 0;
    exp_54_ram[3752] = 0;
    exp_54_ram[3753] = 252;
    exp_54_ram[3754] = 252;
    exp_54_ram[3755] = 64;
    exp_54_ram[3756] = 0;
    exp_54_ram[3757] = 1;
    exp_54_ram[3758] = 64;
    exp_54_ram[3759] = 65;
    exp_54_ram[3760] = 0;
    exp_54_ram[3761] = 0;
    exp_54_ram[3762] = 13;
    exp_54_ram[3763] = 250;
    exp_54_ram[3764] = 250;
    exp_54_ram[3765] = 250;
    exp_54_ram[3766] = 250;
    exp_54_ram[3767] = 0;
    exp_54_ram[3768] = 0;
    exp_54_ram[3769] = 232;
    exp_54_ram[3770] = 0;
    exp_54_ram[3771] = 0;
    exp_54_ram[3772] = 0;
    exp_54_ram[3773] = 0;
    exp_54_ram[3774] = 0;
    exp_54_ram[3775] = 232;
    exp_54_ram[3776] = 252;
    exp_54_ram[3777] = 0;
    exp_54_ram[3778] = 148;
    exp_54_ram[3779] = 184;
    exp_54_ram[3780] = 253;
    exp_54_ram[3781] = 252;
    exp_54_ram[3782] = 252;
    exp_54_ram[3783] = 252;
    exp_54_ram[3784] = 6;
    exp_54_ram[3785] = 251;
    exp_54_ram[3786] = 18;
    exp_54_ram[3787] = 103;
    exp_54_ram[3788] = 2;
    exp_54_ram[3789] = 250;
    exp_54_ram[3790] = 251;
    exp_54_ram[3791] = 18;
    exp_54_ram[3792] = 103;
    exp_54_ram[3793] = 2;
    exp_54_ram[3794] = 250;
    exp_54_ram[3795] = 251;
    exp_54_ram[3796] = 18;
    exp_54_ram[3797] = 103;
    exp_54_ram[3798] = 2;
    exp_54_ram[3799] = 250;
    exp_54_ram[3800] = 251;
    exp_54_ram[3801] = 18;
    exp_54_ram[3802] = 103;
    exp_54_ram[3803] = 2;
    exp_54_ram[3804] = 250;
    exp_54_ram[3805] = 252;
    exp_54_ram[3806] = 0;
    exp_54_ram[3807] = 252;
    exp_54_ram[3808] = 246;
    exp_54_ram[3809] = 0;
    exp_54_ram[3810] = 0;
    exp_54_ram[3811] = 252;
    exp_54_ram[3812] = 252;
    exp_54_ram[3813] = 64;
    exp_54_ram[3814] = 0;
    exp_54_ram[3815] = 1;
    exp_54_ram[3816] = 64;
    exp_54_ram[3817] = 65;
    exp_54_ram[3818] = 0;
    exp_54_ram[3819] = 0;
    exp_54_ram[3820] = 13;
    exp_54_ram[3821] = 248;
    exp_54_ram[3822] = 248;
    exp_54_ram[3823] = 249;
    exp_54_ram[3824] = 249;
    exp_54_ram[3825] = 0;
    exp_54_ram[3826] = 0;
    exp_54_ram[3827] = 244;
    exp_54_ram[3828] = 0;
    exp_54_ram[3829] = 0;
    exp_54_ram[3830] = 0;
    exp_54_ram[3831] = 0;
    exp_54_ram[3832] = 0;
    exp_54_ram[3833] = 244;
    exp_54_ram[3834] = 252;
    exp_54_ram[3835] = 0;
    exp_54_ram[3836] = 151;
    exp_54_ram[3837] = 170;
    exp_54_ram[3838] = 238;
    exp_54_ram[3839] = 252;
    exp_54_ram[3840] = 252;
    exp_54_ram[3841] = 252;
    exp_54_ram[3842] = 13;
    exp_54_ram[3843] = 251;
    exp_54_ram[3844] = 251;
    exp_54_ram[3845] = 18;
    exp_54_ram[3846] = 103;
    exp_54_ram[3847] = 0;
    exp_54_ram[3848] = 0;
    exp_54_ram[3849] = 0;
    exp_54_ram[3850] = 198;
    exp_54_ram[3851] = 0;
    exp_54_ram[3852] = 0;
    exp_54_ram[3853] = 250;
    exp_54_ram[3854] = 250;
    exp_54_ram[3855] = 251;
    exp_54_ram[3856] = 251;
    exp_54_ram[3857] = 18;
    exp_54_ram[3858] = 103;
    exp_54_ram[3859] = 0;
    exp_54_ram[3860] = 0;
    exp_54_ram[3861] = 0;
    exp_54_ram[3862] = 195;
    exp_54_ram[3863] = 0;
    exp_54_ram[3864] = 0;
    exp_54_ram[3865] = 250;
    exp_54_ram[3866] = 250;
    exp_54_ram[3867] = 251;
    exp_54_ram[3868] = 251;
    exp_54_ram[3869] = 18;
    exp_54_ram[3870] = 103;
    exp_54_ram[3871] = 0;
    exp_54_ram[3872] = 0;
    exp_54_ram[3873] = 0;
    exp_54_ram[3874] = 192;
    exp_54_ram[3875] = 0;
    exp_54_ram[3876] = 0;
    exp_54_ram[3877] = 250;
    exp_54_ram[3878] = 250;
    exp_54_ram[3879] = 251;
    exp_54_ram[3880] = 251;
    exp_54_ram[3881] = 18;
    exp_54_ram[3882] = 103;
    exp_54_ram[3883] = 0;
    exp_54_ram[3884] = 0;
    exp_54_ram[3885] = 0;
    exp_54_ram[3886] = 189;
    exp_54_ram[3887] = 0;
    exp_54_ram[3888] = 0;
    exp_54_ram[3889] = 250;
    exp_54_ram[3890] = 250;
    exp_54_ram[3891] = 252;
    exp_54_ram[3892] = 0;
    exp_54_ram[3893] = 252;
    exp_54_ram[3894] = 224;
    exp_54_ram[3895] = 0;
    exp_54_ram[3896] = 0;
    exp_54_ram[3897] = 252;
    exp_54_ram[3898] = 252;
    exp_54_ram[3899] = 64;
    exp_54_ram[3900] = 0;
    exp_54_ram[3901] = 1;
    exp_54_ram[3902] = 64;
    exp_54_ram[3903] = 65;
    exp_54_ram[3904] = 0;
    exp_54_ram[3905] = 0;
    exp_54_ram[3906] = 13;
    exp_54_ram[3907] = 0;
    exp_54_ram[3908] = 0;
    exp_54_ram[3909] = 0;
    exp_54_ram[3910] = 0;
    exp_54_ram[3911] = 238;
    exp_54_ram[3912] = 0;
    exp_54_ram[3913] = 0;
    exp_54_ram[3914] = 0;
    exp_54_ram[3915] = 0;
    exp_54_ram[3916] = 0;
    exp_54_ram[3917] = 236;
    exp_54_ram[3918] = 252;
    exp_54_ram[3919] = 0;
    exp_54_ram[3920] = 153;
    exp_54_ram[3921] = 149;
    exp_54_ram[3922] = 0;
    exp_54_ram[3923] = 6;
    exp_54_ram[3924] = 6;
    exp_54_ram[3925] = 6;
    exp_54_ram[3926] = 6;
    exp_54_ram[3927] = 5;
    exp_54_ram[3928] = 5;
    exp_54_ram[3929] = 5;
    exp_54_ram[3930] = 5;
    exp_54_ram[3931] = 4;
    exp_54_ram[3932] = 4;
    exp_54_ram[3933] = 4;
    exp_54_ram[3934] = 4;
    exp_54_ram[3935] = 7;
    exp_54_ram[3936] = 0;
    exp_54_ram[3937] = 250;
    exp_54_ram[3938] = 4;
    exp_54_ram[3939] = 4;
    exp_54_ram[3940] = 5;
    exp_54_ram[3941] = 5;
    exp_54_ram[3942] = 5;
    exp_54_ram[3943] = 5;
    exp_54_ram[3944] = 6;
    exp_54_ram[3945] = 0;
    exp_54_ram[3946] = 156;
    exp_54_ram[3947] = 142;
    exp_54_ram[3948] = 134;
    exp_54_ram[3949] = 0;
    exp_54_ram[3950] = 137;
    exp_54_ram[3951] = 252;
    exp_54_ram[3952] = 0;
    exp_54_ram[3953] = 156;
    exp_54_ram[3954] = 141;
    exp_54_ram[3955] = 132;
    exp_54_ram[3956] = 0;
    exp_54_ram[3957] = 255;
    exp_54_ram[3958] = 252;
    exp_54_ram[3959] = 0;
    exp_54_ram[3960] = 157;
    exp_54_ram[3961] = 139;
    exp_54_ram[3962] = 130;
    exp_54_ram[3963] = 0;
    exp_54_ram[3964] = 250;
    exp_54_ram[3965] = 0;
    exp_54_ram[3966] = 157;
    exp_54_ram[3967] = 137;
    exp_54_ram[3968] = 129;
    exp_54_ram[3969] = 0;
    exp_54_ram[3970] = 250;
    exp_54_ram[3971] = 0;
    exp_54_ram[3972] = 158;
    exp_54_ram[3973] = 136;
    exp_54_ram[3974] = 255;
    exp_54_ram[3975] = 0;
    exp_54_ram[3976] = 250;
    exp_54_ram[3977] = 3;
    exp_54_ram[3978] = 250;
    exp_54_ram[3979] = 0;
    exp_54_ram[3980] = 252;
    exp_54_ram[3981] = 251;
    exp_54_ram[3982] = 0;
    exp_54_ram[3983] = 150;
    exp_54_ram[3984] = 0;
    exp_54_ram[3985] = 0;
    exp_54_ram[3986] = 250;
    exp_54_ram[3987] = 250;
    exp_54_ram[3988] = 251;
    exp_54_ram[3989] = 0;
    exp_54_ram[3990] = 223;
    exp_54_ram[3991] = 0;
    exp_54_ram[3992] = 0;
    exp_54_ram[3993] = 224;
    exp_54_ram[3994] = 250;
    exp_54_ram[3995] = 0;
    exp_54_ram[3996] = 161;
    exp_54_ram[3997] = 0;
    exp_54_ram[3998] = 0;
    exp_54_ram[3999] = 222;
    exp_54_ram[4000] = 250;
    exp_54_ram[4001] = 250;
    exp_54_ram[4002] = 0;
    exp_54_ram[4003] = 0;
    exp_54_ram[4004] = 208;
    exp_54_ram[4005] = 0;
    exp_54_ram[4006] = 193;
    exp_54_ram[4007] = 0;
    exp_54_ram[4008] = 0;
    exp_54_ram[4009] = 250;
    exp_54_ram[4010] = 250;
    exp_54_ram[4011] = 250;
    exp_54_ram[4012] = 0;
    exp_54_ram[4013] = 157;
    exp_54_ram[4014] = 0;
    exp_54_ram[4015] = 0;
    exp_54_ram[4016] = 218;
    exp_54_ram[4017] = 194;
    exp_54_ram[4018] = 252;
    exp_54_ram[4019] = 252;
    exp_54_ram[4020] = 252;
    exp_54_ram[4021] = 13;
    exp_54_ram[4022] = 0;
    exp_54_ram[4023] = 192;
    exp_54_ram[4024] = 0;
    exp_54_ram[4025] = 0;
    exp_54_ram[4026] = 253;
    exp_54_ram[4027] = 253;
    exp_54_ram[4028] = 0;
    exp_54_ram[4029] = 0;
    exp_54_ram[4030] = 197;
    exp_54_ram[4031] = 0;
    exp_54_ram[4032] = 0;
    exp_54_ram[4033] = 0;
    exp_54_ram[4034] = 13;
    exp_54_ram[4035] = 0;
    exp_54_ram[4036] = 233;
    exp_54_ram[4037] = 0;
    exp_54_ram[4038] = 0;
    exp_54_ram[4039] = 0;
    exp_54_ram[4040] = 0;
    exp_54_ram[4041] = 0;
    exp_54_ram[4042] = 0;
    exp_54_ram[4043] = 217;
    exp_54_ram[4044] = 0;
    exp_54_ram[4045] = 250;
    exp_54_ram[4046] = 0;
    exp_54_ram[4047] = 13;
    exp_54_ram[4048] = 0;
    exp_54_ram[4049] = 0;
    exp_54_ram[4050] = 253;
    exp_54_ram[4051] = 253;
    exp_54_ram[4052] = 1;
    exp_54_ram[4053] = 0;
    exp_54_ram[4054] = 0;
    exp_54_ram[4055] = 1;
    exp_54_ram[4056] = 0;
    exp_54_ram[4057] = 0;
    exp_54_ram[4058] = 252;
    exp_54_ram[4059] = 252;
    exp_54_ram[4060] = 0;
    exp_54_ram[4061] = 179;
    exp_54_ram[4062] = 0;
    exp_54_ram[4063] = 0;
    exp_54_ram[4064] = 250;
    exp_54_ram[4065] = 250;
    exp_54_ram[4066] = 250;
    exp_54_ram[4067] = 0;
    exp_54_ram[4068] = 143;
    exp_54_ram[4069] = 0;
    exp_54_ram[4070] = 0;
    exp_54_ram[4071] = 204;
    exp_54_ram[4072] = 253;
    exp_54_ram[4073] = 0;
    exp_54_ram[4074] = 252;
    exp_54_ram[4075] = 253;
    exp_54_ram[4076] = 6;
    exp_54_ram[4077] = 242;
    exp_54_ram[4078] = 0;
    exp_54_ram[4079] = 0;
    exp_54_ram[4080] = 5;
    exp_54_ram[4081] = 5;
    exp_54_ram[4082] = 5;
    exp_54_ram[4083] = 5;
    exp_54_ram[4084] = 4;
    exp_54_ram[4085] = 4;
    exp_54_ram[4086] = 6;
    exp_54_ram[4087] = 0;
    exp_54_ram[4088] = 254;
    exp_54_ram[4089] = 0;
    exp_54_ram[4090] = 0;
    exp_54_ram[4091] = 2;
    exp_54_ram[4092] = 0;
    exp_54_ram[4093] = 159;
    exp_54_ram[4094] = 234;
    exp_54_ram[4095] = 0;
    exp_54_ram[4096] = 160;
    exp_54_ram[4097] = 233;
    exp_54_ram[4098] = 0;
    exp_54_ram[4099] = 161;
    exp_54_ram[4100] = 232;
    exp_54_ram[4101] = 0;
    exp_54_ram[4102] = 162;
    exp_54_ram[4103] = 231;
    exp_54_ram[4104] = 0;
    exp_54_ram[4105] = 164;
    exp_54_ram[4106] = 231;
    exp_54_ram[4107] = 185;
    exp_54_ram[4108] = 0;
    exp_54_ram[4109] = 254;
    exp_54_ram[4110] = 254;
    exp_54_ram[4111] = 6;
    exp_54_ram[4112] = 4;
    exp_54_ram[4113] = 6;
    exp_54_ram[4114] = 250;
    exp_54_ram[4115] = 6;
    exp_54_ram[4116] = 2;
    exp_54_ram[4117] = 6;
    exp_54_ram[4118] = 248;
    exp_54_ram[4119] = 6;
    exp_54_ram[4120] = 0;
    exp_54_ram[4121] = 6;
    exp_54_ram[4122] = 0;
    exp_54_ram[4123] = 2;
    exp_54_ram[4124] = 232;
    exp_54_ram[4125] = 1;
    exp_54_ram[4126] = 234;
    exp_54_ram[4127] = 1;
    exp_54_ram[4128] = 251;
    exp_54_ram[4129] = 0;
    exp_54_ram[4130] = 207;
    exp_54_ram[4131] = 0;
    exp_54_ram[4132] = 246;
    exp_54_ram[4133] = 0;
    exp_54_ram[4134] = 0;
    exp_54_ram[4135] = 2;
    exp_54_ram[4136] = 255;
    exp_54_ram[4137] = 2;
    exp_54_ram[4138] = 0;
    exp_54_ram[4139] = 0;
    exp_54_ram[4140] = 0;
    exp_54_ram[4141] = 64;
    exp_54_ram[4142] = 1;
    exp_54_ram[4143] = 0;
    exp_54_ram[4144] = 254;
    exp_54_ram[4145] = 255;
    exp_54_ram[4146] = 0;
    exp_54_ram[4147] = 254;
    exp_54_ram[4148] = 2;
    exp_54_ram[4149] = 128;
    exp_54_ram[4150] = 128;
    exp_54_ram[4151] = 128;
    exp_54_ram[4152] = 0;
    exp_54_ram[4153] = 0;
    exp_54_ram[4154] = 0;
    exp_54_ram[4155] = 0;
    exp_54_ram[4156] = 0;
    exp_54_ram[4157] = 0;
    exp_54_ram[4158] = 0;
    exp_54_ram[4159] = 0;
    exp_54_ram[4160] = 0;
    exp_54_ram[4161] = 0;
    exp_54_ram[4162] = 0;
    exp_54_ram[4163] = 0;
    exp_54_ram[4164] = 0;
    exp_54_ram[4165] = 0;
    exp_54_ram[4166] = 0;
    exp_54_ram[4167] = 0;
    exp_54_ram[4168] = 0;
    exp_54_ram[4169] = 0;
    exp_54_ram[4170] = 0;
    exp_54_ram[4171] = 0;
    exp_54_ram[4172] = 0;
    exp_54_ram[4173] = 0;
    exp_54_ram[4174] = 0;
    exp_54_ram[4175] = 0;
    exp_54_ram[4176] = 0;
    exp_54_ram[4177] = 0;
    exp_54_ram[4178] = 0;
    exp_54_ram[4179] = 0;
    exp_54_ram[4180] = 0;
    exp_54_ram[4181] = 0;
    exp_54_ram[4182] = 0;
    exp_54_ram[4183] = 0;
    exp_54_ram[4184] = 0;
    exp_54_ram[4185] = 0;
    exp_54_ram[4186] = 0;
    exp_54_ram[4187] = 0;
    exp_54_ram[4188] = 0;
    exp_54_ram[4189] = 0;
    exp_54_ram[4190] = 0;
    exp_54_ram[4191] = 0;
    exp_54_ram[4192] = 0;
    exp_54_ram[4193] = 0;
    exp_54_ram[4194] = 0;
    exp_54_ram[4195] = 0;
    exp_54_ram[4196] = 0;
    exp_54_ram[4197] = 0;
    exp_54_ram[4198] = 0;
    exp_54_ram[4199] = 0;
    exp_54_ram[4200] = 0;
    exp_54_ram[4201] = 0;
    exp_54_ram[4202] = 0;
    exp_54_ram[4203] = 0;
    exp_54_ram[4204] = 0;
    exp_54_ram[4205] = 0;
    exp_54_ram[4206] = 0;
    exp_54_ram[4207] = 0;
    exp_54_ram[4208] = 0;
    exp_54_ram[4209] = 0;
    exp_54_ram[4210] = 0;
    exp_54_ram[4211] = 0;
    exp_54_ram[4212] = 0;
    exp_54_ram[4213] = 0;
    exp_54_ram[4214] = 0;
    exp_54_ram[4215] = 0;
    exp_54_ram[4216] = 0;
    exp_54_ram[4217] = 0;
    exp_54_ram[4218] = 0;
    exp_54_ram[4219] = 0;
    exp_54_ram[4220] = 0;
    exp_54_ram[4221] = 0;
    exp_54_ram[4222] = 0;
    exp_54_ram[4223] = 0;
    exp_54_ram[4224] = 0;
    exp_54_ram[4225] = 0;
    exp_54_ram[4226] = 0;
    exp_54_ram[4227] = 0;
    exp_54_ram[4228] = 0;
    exp_54_ram[4229] = 0;
    exp_54_ram[4230] = 0;
    exp_54_ram[4231] = 0;
    exp_54_ram[4232] = 0;
    exp_54_ram[4233] = 0;
    exp_54_ram[4234] = 0;
    exp_54_ram[4235] = 0;
    exp_54_ram[4236] = 0;
    exp_54_ram[4237] = 0;
    exp_54_ram[4238] = 0;
    exp_54_ram[4239] = 0;
    exp_54_ram[4240] = 0;
    exp_54_ram[4241] = 0;
    exp_54_ram[4242] = 0;
    exp_54_ram[4243] = 0;
    exp_54_ram[4244] = 0;
    exp_54_ram[4245] = 0;
    exp_54_ram[4246] = 0;
    exp_54_ram[4247] = 0;
    exp_54_ram[4248] = 0;
    exp_54_ram[4249] = 0;
    exp_54_ram[4250] = 0;
    exp_54_ram[4251] = 0;
    exp_54_ram[4252] = 0;
    exp_54_ram[4253] = 0;
    exp_54_ram[4254] = 0;
    exp_54_ram[4255] = 0;
    exp_54_ram[4256] = 0;
    exp_54_ram[4257] = 0;
    exp_54_ram[4258] = 0;
    exp_54_ram[4259] = 0;
    exp_54_ram[4260] = 0;
    exp_54_ram[4261] = 0;
    exp_54_ram[4262] = 0;
    exp_54_ram[4263] = 0;
    exp_54_ram[4264] = 0;
    exp_54_ram[4265] = 0;
    exp_54_ram[4266] = 0;
    exp_54_ram[4267] = 0;
    exp_54_ram[4268] = 0;
    exp_54_ram[4269] = 0;
    exp_54_ram[4270] = 0;
    exp_54_ram[4271] = 0;
    exp_54_ram[4272] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_398;
  assign exp_398 = exp_679;

  reg [3:0] exp_679_reg;
  always@(*) begin
    case (exp_531)
      0:exp_679_reg <= exp_666;
      1:exp_679_reg <= exp_671;
      2:exp_679_reg <= exp_672;
      3:exp_679_reg <= exp_673;
      4:exp_679_reg <= exp_674;
      5:exp_679_reg <= exp_675;
      6:exp_679_reg <= exp_676;
      7:exp_679_reg <= exp_677;
      default:exp_679_reg <= exp_678;
    endcase
  end
  assign exp_679 = exp_679_reg;
  assign exp_678 = 0;
  assign exp_666 = exp_662 << exp_665;
  assign exp_662 = 1;
  assign exp_665 = exp_664 + exp_663;
  assign exp_664 = 0;
  assign exp_663 = exp_599[1:0];
  assign exp_671 = exp_667 << exp_670;
  assign exp_667 = 3;
  assign exp_670 = exp_669 + exp_668;
  assign exp_669 = 0;
  assign exp_668 = exp_599[1:1];
  assign exp_672 = 15;
  assign exp_673 = 0;
  assign exp_674 = 0;
  assign exp_675 = 0;
  assign exp_676 = 0;
  assign exp_677 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_393;
  assign exp_393 = exp_661;

  reg [31:0] exp_661_reg;
  always@(*) begin
    case (exp_531)
      0:exp_661_reg <= exp_648;
      1:exp_661_reg <= exp_652;
      2:exp_661_reg <= exp_654;
      3:exp_661_reg <= exp_655;
      4:exp_661_reg <= exp_656;
      5:exp_661_reg <= exp_657;
      6:exp_661_reg <= exp_658;
      7:exp_661_reg <= exp_659;
      default:exp_661_reg <= exp_660;
    endcase
  end
  assign exp_661 = exp_661_reg;
  assign exp_660 = 0;

  reg [31:0] exp_648_reg;
  always@(*) begin
    case (exp_602)
      0:exp_648_reg <= exp_634;
      1:exp_648_reg <= exp_642;
      2:exp_648_reg <= exp_644;
      3:exp_648_reg <= exp_646;
      default:exp_648_reg <= exp_647;
    endcase
  end
  assign exp_648 = exp_648_reg;
  assign exp_647 = 0;
  assign exp_634 = exp_633;
  assign exp_633 = exp_632 + exp_631;
  assign exp_632 = 0;
  assign exp_631 = exp_521[7:0];

      reg [31:0] exp_521_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_521_reg <= exp_464;
        end
      end
      assign exp_521 = exp_521_reg;
      assign exp_642 = exp_634 << exp_641;
  assign exp_641 = 8;
  assign exp_644 = exp_634 << exp_643;
  assign exp_643 = 16;
  assign exp_646 = exp_634 << exp_645;
  assign exp_645 = 24;

  reg [31:0] exp_652_reg;
  always@(*) begin
    case (exp_605)
      0:exp_652_reg <= exp_638;
      1:exp_652_reg <= exp_650;
      default:exp_652_reg <= exp_651;
    endcase
  end
  assign exp_652 = exp_652_reg;
  assign exp_605 = exp_604 + exp_603;
  assign exp_604 = 0;
  assign exp_603 = exp_599[1:1];
  assign exp_651 = 0;
  assign exp_638 = exp_637;
  assign exp_637 = exp_636 + exp_635;
  assign exp_636 = 0;
  assign exp_635 = exp_521[15:0];
  assign exp_650 = exp_638 << exp_649;
  assign exp_649 = 16;
  assign exp_654 = exp_653 + exp_640;
  assign exp_653 = 0;
  assign exp_640 = exp_639 + exp_521;
  assign exp_639 = 0;
  assign exp_655 = 0;
  assign exp_656 = 0;
  assign exp_657 = 0;
  assign exp_658 = 0;
  assign exp_659 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 0;
    exp_47_ram[32] = 1;
    exp_47_ram[33] = 208;
    exp_47_ram[34] = 0;
    exp_47_ram[35] = 5;
    exp_47_ram[36] = 5;
    exp_47_ram[37] = 6;
    exp_47_ram[38] = 6;
    exp_47_ram[39] = 8;
    exp_47_ram[40] = 6;
    exp_47_ram[41] = 0;
    exp_47_ram[42] = 6;
    exp_47_ram[43] = 197;
    exp_47_ram[44] = 1;
    exp_47_ram[45] = 230;
    exp_47_ram[46] = 240;
    exp_47_ram[47] = 199;
    exp_47_ram[48] = 55;
    exp_47_ram[49] = 230;
    exp_47_ram[50] = 166;
    exp_47_ram[51] = 6;
    exp_47_ram[52] = 0;
    exp_47_ram[53] = 230;
    exp_47_ram[54] = 229;
    exp_47_ram[55] = 229;
    exp_47_ram[56] = 215;
    exp_47_ram[57] = 232;
    exp_47_ram[58] = 214;
    exp_47_ram[59] = 183;
    exp_47_ram[60] = 216;
    exp_47_ram[61] = 8;
    exp_47_ram[62] = 21;
    exp_47_ram[63] = 8;
    exp_47_ram[64] = 6;
    exp_47_ram[65] = 3;
    exp_47_ram[66] = 21;
    exp_47_ram[67] = 6;
    exp_47_ram[68] = 214;
    exp_47_ram[69] = 7;
    exp_47_ram[70] = 247;
    exp_47_ram[71] = 183;
    exp_47_ram[72] = 7;
    exp_47_ram[73] = 246;
    exp_47_ram[74] = 7;
    exp_47_ram[75] = 183;
    exp_47_ram[76] = 230;
    exp_47_ram[77] = 7;
    exp_47_ram[78] = 183;
    exp_47_ram[79] = 23;
    exp_47_ram[80] = 3;
    exp_47_ram[81] = 3;
    exp_47_ram[82] = 23;
    exp_47_ram[83] = 7;
    exp_47_ram[84] = 103;
    exp_47_ram[85] = 246;
    exp_47_ram[86] = 7;
    exp_47_ram[87] = 211;
    exp_47_ram[88] = 104;
    exp_47_ram[89] = 247;
    exp_47_ram[90] = 3;
    exp_47_ram[91] = 211;
    exp_47_ram[92] = 231;
    exp_47_ram[93] = 5;
    exp_47_ram[94] = 197;
    exp_47_ram[95] = 0;
    exp_47_ram[96] = 64;
    exp_47_ram[97] = 0;
    exp_47_ram[98] = 0;
    exp_47_ram[99] = 166;
    exp_47_ram[100] = 128;
    exp_47_ram[101] = 31;
    exp_47_ram[102] = 6;
    exp_47_ram[103] = 16;
    exp_47_ram[104] = 199;
    exp_47_ram[105] = 1;
    exp_47_ram[106] = 232;
    exp_47_ram[107] = 240;
    exp_47_ram[108] = 7;
    exp_47_ram[109] = 128;
    exp_47_ram[110] = 168;
    exp_47_ram[111] = 230;
    exp_47_ram[112] = 6;
    exp_47_ram[113] = 0;
    exp_47_ram[114] = 167;
    exp_47_ram[115] = 230;
    exp_47_ram[116] = 230;
    exp_47_ram[117] = 7;
    exp_47_ram[118] = 16;
    exp_47_ram[119] = 8;
    exp_47_ram[120] = 8;
    exp_47_ram[121] = 6;
    exp_47_ram[122] = 3;
    exp_47_ram[123] = 23;
    exp_47_ram[124] = 23;
    exp_47_ram[125] = 6;
    exp_47_ram[126] = 230;
    exp_47_ram[127] = 246;
    exp_47_ram[128] = 7;
    exp_47_ram[129] = 199;
    exp_47_ram[130] = 7;
    exp_47_ram[131] = 247;
    exp_47_ram[132] = 7;
    exp_47_ram[133] = 199;
    exp_47_ram[134] = 231;
    exp_47_ram[135] = 7;
    exp_47_ram[136] = 199;
    exp_47_ram[137] = 23;
    exp_47_ram[138] = 3;
    exp_47_ram[139] = 3;
    exp_47_ram[140] = 23;
    exp_47_ram[141] = 7;
    exp_47_ram[142] = 103;
    exp_47_ram[143] = 230;
    exp_47_ram[144] = 7;
    exp_47_ram[145] = 211;
    exp_47_ram[146] = 104;
    exp_47_ram[147] = 247;
    exp_47_ram[148] = 3;
    exp_47_ram[149] = 211;
    exp_47_ram[150] = 231;
    exp_47_ram[151] = 5;
    exp_47_ram[152] = 197;
    exp_47_ram[153] = 0;
    exp_47_ram[154] = 0;
    exp_47_ram[155] = 0;
    exp_47_ram[156] = 232;
    exp_47_ram[157] = 128;
    exp_47_ram[158] = 31;
    exp_47_ram[159] = 216;
    exp_47_ram[160] = 231;
    exp_47_ram[161] = 216;
    exp_47_ram[162] = 215;
    exp_47_ram[163] = 232;
    exp_47_ram[164] = 8;
    exp_47_ram[165] = 247;
    exp_47_ram[166] = 21;
    exp_47_ram[167] = 8;
    exp_47_ram[168] = 7;
    exp_47_ram[169] = 6;
    exp_47_ram[170] = 21;
    exp_47_ram[171] = 7;
    exp_47_ram[172] = 183;
    exp_47_ram[173] = 167;
    exp_47_ram[174] = 5;
    exp_47_ram[175] = 215;
    exp_47_ram[176] = 7;
    exp_47_ram[177] = 245;
    exp_47_ram[178] = 7;
    exp_47_ram[179] = 215;
    exp_47_ram[180] = 229;
    exp_47_ram[181] = 7;
    exp_47_ram[182] = 215;
    exp_47_ram[183] = 22;
    exp_47_ram[184] = 6;
    exp_47_ram[185] = 6;
    exp_47_ram[186] = 22;
    exp_47_ram[187] = 7;
    exp_47_ram[188] = 215;
    exp_47_ram[189] = 199;
    exp_47_ram[190] = 6;
    exp_47_ram[191] = 167;
    exp_47_ram[192] = 7;
    exp_47_ram[193] = 246;
    exp_47_ram[194] = 7;
    exp_47_ram[195] = 167;
    exp_47_ram[196] = 230;
    exp_47_ram[197] = 7;
    exp_47_ram[198] = 5;
    exp_47_ram[199] = 167;
    exp_47_ram[200] = 229;
    exp_47_ram[201] = 159;
    exp_47_ram[202] = 213;
    exp_47_ram[203] = 1;
    exp_47_ram[204] = 230;
    exp_47_ram[205] = 240;
    exp_47_ram[206] = 215;
    exp_47_ram[207] = 53;
    exp_47_ram[208] = 0;
    exp_47_ram[209] = 182;
    exp_47_ram[210] = 7;
    exp_47_ram[211] = 167;
    exp_47_ram[212] = 7;
    exp_47_ram[213] = 0;
    exp_47_ram[214] = 183;
    exp_47_ram[215] = 229;
    exp_47_ram[216] = 229;
    exp_47_ram[217] = 16;
    exp_47_ram[218] = 246;
    exp_47_ram[219] = 200;
    exp_47_ram[220] = 21;
    exp_47_ram[221] = 31;
    exp_47_ram[222] = 0;
    exp_47_ram[223] = 0;
    exp_47_ram[224] = 230;
    exp_47_ram[225] = 128;
    exp_47_ram[226] = 159;
    exp_47_ram[227] = 230;
    exp_47_ram[228] = 182;
    exp_47_ram[229] = 216;
    exp_47_ram[230] = 231;
    exp_47_ram[231] = 8;
    exp_47_ram[232] = 222;
    exp_47_ram[233] = 183;
    exp_47_ram[234] = 232;
    exp_47_ram[235] = 182;
    exp_47_ram[236] = 247;
    exp_47_ram[237] = 8;
    exp_47_ram[238] = 7;
    exp_47_ram[239] = 6;
    exp_47_ram[240] = 222;
    exp_47_ram[241] = 6;
    exp_47_ram[242] = 230;
    exp_47_ram[243] = 199;
    exp_47_ram[244] = 14;
    exp_47_ram[245] = 231;
    exp_47_ram[246] = 7;
    exp_47_ram[247] = 254;
    exp_47_ram[248] = 7;
    exp_47_ram[249] = 231;
    exp_47_ram[250] = 238;
    exp_47_ram[251] = 7;
    exp_47_ram[252] = 231;
    exp_47_ram[253] = 215;
    exp_47_ram[254] = 215;
    exp_47_ram[255] = 6;
    exp_47_ram[256] = 231;
    exp_47_ram[257] = 6;
    exp_47_ram[258] = 7;
    exp_47_ram[259] = 246;
    exp_47_ram[260] = 7;
    exp_47_ram[261] = 199;
    exp_47_ram[262] = 7;
    exp_47_ram[263] = 247;
    exp_47_ram[264] = 7;
    exp_47_ram[265] = 199;
    exp_47_ram[266] = 231;
    exp_47_ram[267] = 7;
    exp_47_ram[268] = 5;
    exp_47_ram[269] = 1;
    exp_47_ram[270] = 197;
    exp_47_ram[271] = 254;
    exp_47_ram[272] = 213;
    exp_47_ram[273] = 5;
    exp_47_ram[274] = 211;
    exp_47_ram[275] = 3;
    exp_47_ram[276] = 199;
    exp_47_ram[277] = 216;
    exp_47_ram[278] = 214;
    exp_47_ram[279] = 14;
    exp_47_ram[280] = 104;
    exp_47_ram[281] = 216;
    exp_47_ram[282] = 7;
    exp_47_ram[283] = 102;
    exp_47_ram[284] = 215;
    exp_47_ram[285] = 214;
    exp_47_ram[286] = 7;
    exp_47_ram[287] = 198;
    exp_47_ram[288] = 199;
    exp_47_ram[289] = 199;
    exp_47_ram[290] = 1;
    exp_47_ram[291] = 247;
    exp_47_ram[292] = 247;
    exp_47_ram[293] = 7;
    exp_47_ram[294] = 254;
    exp_47_ram[295] = 184;
    exp_47_ram[296] = 199;
    exp_47_ram[297] = 0;
    exp_47_ram[298] = 232;
    exp_47_ram[299] = 245;
    exp_47_ram[300] = 223;
    exp_47_ram[301] = 0;
    exp_47_ram[302] = 0;
    exp_47_ram[303] = 159;
    exp_47_ram[304] = 16;
    exp_47_ram[305] = 247;
    exp_47_ram[306] = 69;
    exp_47_ram[307] = 183;
    exp_47_ram[308] = 5;
    exp_47_ram[309] = 5;
    exp_47_ram[310] = 248;
    exp_47_ram[311] = 245;
    exp_47_ram[312] = 240;
    exp_47_ram[313] = 70;
    exp_47_ram[314] = 215;
    exp_47_ram[315] = 6;
    exp_47_ram[316] = 245;
    exp_47_ram[317] = 246;
    exp_47_ram[318] = 216;
    exp_47_ram[319] = 248;
    exp_47_ram[320] = 14;
    exp_47_ram[321] = 32;
    exp_47_ram[322] = 0;
    exp_47_ram[323] = 213;
    exp_47_ram[324] = 199;
    exp_47_ram[325] = 14;
    exp_47_ram[326] = 8;
    exp_47_ram[327] = 248;
    exp_47_ram[328] = 23;
    exp_47_ram[329] = 5;
    exp_47_ram[330] = 199;
    exp_47_ram[331] = 6;
    exp_47_ram[332] = 7;
    exp_47_ram[333] = 213;
    exp_47_ram[334] = 5;
    exp_47_ram[335] = 5;
    exp_47_ram[336] = 240;
    exp_47_ram[337] = 0;
    exp_47_ram[338] = 240;
    exp_47_ram[339] = 6;
    exp_47_ram[340] = 6;
    exp_47_ram[341] = 0;
    exp_47_ram[342] = 184;
    exp_47_ram[343] = 5;
    exp_47_ram[344] = 0;
    exp_47_ram[345] = 23;
    exp_47_ram[346] = 232;
    exp_47_ram[347] = 110;
    exp_47_ram[348] = 195;
    exp_47_ram[349] = 0;
    exp_47_ram[350] = 0;
    exp_47_ram[351] = 16;
    exp_47_ram[352] = 0;
    exp_47_ram[353] = 7;
    exp_47_ram[354] = 95;
    exp_47_ram[355] = 232;
    exp_47_ram[356] = 95;
    exp_47_ram[357] = 5;
    exp_47_ram[358] = 5;
    exp_47_ram[359] = 0;
    exp_47_ram[360] = 159;
    exp_47_ram[361] = 1;
    exp_47_ram[362] = 129;
    exp_47_ram[363] = 17;
    exp_47_ram[364] = 5;
    exp_47_ram[365] = 5;
    exp_47_ram[366] = 64;
    exp_47_ram[367] = 224;
    exp_47_ram[368] = 160;
    exp_47_ram[369] = 167;
    exp_47_ram[370] = 167;
    exp_47_ram[371] = 176;
    exp_47_ram[372] = 167;
    exp_47_ram[373] = 85;
    exp_47_ram[374] = 244;
    exp_47_ram[375] = 164;
    exp_47_ram[376] = 193;
    exp_47_ram[377] = 4;
    exp_47_ram[378] = 199;
    exp_47_ram[379] = 129;
    exp_47_ram[380] = 71;
    exp_47_ram[381] = 199;
    exp_47_ram[382] = 247;
    exp_47_ram[383] = 6;
    exp_47_ram[384] = 1;
    exp_47_ram[385] = 0;
    exp_47_ram[386] = 85;
    exp_47_ram[387] = 244;
    exp_47_ram[388] = 0;
    exp_47_ram[389] = 223;
    exp_47_ram[390] = 0;
    exp_47_ram[391] = 0;
    exp_47_ram[392] = 31;
    exp_47_ram[393] = 1;
    exp_47_ram[394] = 17;
    exp_47_ram[395] = 129;
    exp_47_ram[396] = 145;
    exp_47_ram[397] = 33;
    exp_47_ram[398] = 49;
    exp_47_ram[399] = 65;
    exp_47_ram[400] = 181;
    exp_47_ram[401] = 7;
    exp_47_ram[402] = 5;
    exp_47_ram[403] = 5;
    exp_47_ram[404] = 5;
    exp_47_ram[405] = 5;
    exp_47_ram[406] = 5;
    exp_47_ram[407] = 0;
    exp_47_ram[408] = 5;
    exp_47_ram[409] = 224;
    exp_47_ram[410] = 58;
    exp_47_ram[411] = 48;
    exp_47_ram[412] = 71;
    exp_47_ram[413] = 176;
    exp_47_ram[414] = 4;
    exp_47_ram[415] = 55;
    exp_47_ram[416] = 160;
    exp_47_ram[417] = 55;
    exp_47_ram[418] = 176;
    exp_47_ram[419] = 89;
    exp_47_ram[420] = 52;
    exp_47_ram[421] = 148;
    exp_47_ram[422] = 233;
    exp_47_ram[423] = 180;
    exp_47_ram[424] = 228;
    exp_47_ram[425] = 193;
    exp_47_ram[426] = 129;
    exp_47_ram[427] = 196;
    exp_47_ram[428] = 74;
    exp_47_ram[429] = 197;
    exp_47_ram[430] = 186;
    exp_47_ram[431] = 65;
    exp_47_ram[432] = 1;
    exp_47_ram[433] = 193;
    exp_47_ram[434] = 129;
    exp_47_ram[435] = 7;
    exp_47_ram[436] = 7;
    exp_47_ram[437] = 1;
    exp_47_ram[438] = 0;
    exp_47_ram[439] = 0;
    exp_47_ram[440] = 5;
    exp_47_ram[441] = 31;
    exp_47_ram[442] = 89;
    exp_47_ram[443] = 180;
    exp_47_ram[444] = 0;
    exp_47_ram[445] = 31;
    exp_47_ram[446] = 96;
    exp_47_ram[447] = 71;
    exp_47_ram[448] = 137;
    exp_47_ram[449] = 4;
    exp_47_ram[450] = 9;
    exp_47_ram[451] = 128;
    exp_47_ram[452] = 181;
    exp_47_ram[453] = 128;
    exp_47_ram[454] = 160;
    exp_47_ram[455] = 9;
    exp_47_ram[456] = 4;
    exp_47_ram[457] = 54;
    exp_47_ram[458] = 64;
    exp_47_ram[459] = 164;
    exp_47_ram[460] = 5;
    exp_47_ram[461] = 128;
    exp_47_ram[462] = 4;
    exp_47_ram[463] = 9;
    exp_47_ram[464] = 55;
    exp_47_ram[465] = 112;
    exp_47_ram[466] = 55;
    exp_47_ram[467] = 137;
    exp_47_ram[468] = 233;
    exp_47_ram[469] = 128;
    exp_47_ram[470] = 57;
    exp_47_ram[471] = 36;
    exp_47_ram[472] = 185;
    exp_47_ram[473] = 228;
    exp_47_ram[474] = 128;
    exp_47_ram[475] = 247;
    exp_47_ram[476] = 229;
    exp_47_ram[477] = 119;
    exp_47_ram[478] = 7;
    exp_47_ram[479] = 247;
    exp_47_ram[480] = 64;
    exp_47_ram[481] = 215;
    exp_47_ram[482] = 71;
    exp_47_ram[483] = 247;
    exp_47_ram[484] = 245;
    exp_47_ram[485] = 7;
    exp_47_ram[486] = 128;
    exp_47_ram[487] = 229;
    exp_47_ram[488] = 7;
    exp_47_ram[489] = 128;
    exp_47_ram[490] = 247;
    exp_47_ram[491] = 240;
    exp_47_ram[492] = 229;
    exp_47_ram[493] = 58;
    exp_47_ram[494] = 55;
    exp_47_ram[495] = 213;
    exp_47_ram[496] = 245;
    exp_47_ram[497] = 53;
    exp_47_ram[498] = 223;
    exp_47_ram[499] = 137;
    exp_47_ram[500] = 180;
    exp_47_ram[501] = 0;
    exp_47_ram[502] = 31;
    exp_47_ram[503] = 0;
    exp_47_ram[504] = 0;
    exp_47_ram[505] = 0;
    exp_47_ram[506] = 223;
    exp_47_ram[507] = 6;
    exp_47_ram[508] = 0;
    exp_47_ram[509] = 199;
    exp_47_ram[510] = 240;
    exp_47_ram[511] = 6;
    exp_47_ram[512] = 0;
    exp_47_ram[513] = 165;
    exp_47_ram[514] = 7;
    exp_47_ram[515] = 0;
    exp_47_ram[516] = 197;
    exp_47_ram[517] = 197;
    exp_47_ram[518] = 245;
    exp_47_ram[519] = 181;
    exp_47_ram[520] = 159;
    exp_47_ram[521] = 6;
    exp_47_ram[522] = 0;
    exp_47_ram[523] = 199;
    exp_47_ram[524] = 240;
    exp_47_ram[525] = 6;
    exp_47_ram[526] = 0;
    exp_47_ram[527] = 181;
    exp_47_ram[528] = 7;
    exp_47_ram[529] = 0;
    exp_47_ram[530] = 197;
    exp_47_ram[531] = 197;
    exp_47_ram[532] = 245;
    exp_47_ram[533] = 165;
    exp_47_ram[534] = 159;
    exp_47_ram[535] = 1;
    exp_47_ram[536] = 245;
    exp_47_ram[537] = 240;
    exp_47_ram[538] = 167;
    exp_47_ram[539] = 55;
    exp_47_ram[540] = 0;
    exp_47_ram[541] = 0;
    exp_47_ram[542] = 246;
    exp_47_ram[543] = 245;
    exp_47_ram[544] = 7;
    exp_47_ram[545] = 167;
    exp_47_ram[546] = 5;
    exp_47_ram[547] = 166;
    exp_47_ram[548] = 0;
    exp_47_ram[549] = 0;
    exp_47_ram[550] = 0;
    exp_47_ram[551] = 229;
    exp_47_ram[552] = 128;
    exp_47_ram[553] = 223;
    exp_47_ram[554] = 110;
    exp_47_ram[555] = 84;
    exp_47_ram[556] = 101;
    exp_47_ram[557] = 117;
    exp_47_ram[558] = 83;
    exp_47_ram[559] = 0;
    exp_47_ram[560] = 110;
    exp_47_ram[561] = 77;
    exp_47_ram[562] = 112;
    exp_47_ram[563] = 121;
    exp_47_ram[564] = 74;
    exp_47_ram[565] = 117;
    exp_47_ram[566] = 112;
    exp_47_ram[567] = 78;
    exp_47_ram[568] = 101;
    exp_47_ram[569] = 0;
    exp_47_ram[570] = 108;
    exp_47_ram[571] = 87;
    exp_47_ram[572] = 100;
    exp_47_ram[573] = 0;
    exp_47_ram[574] = 110;
    exp_47_ram[575] = 103;
    exp_47_ram[576] = 105;
    exp_47_ram[577] = 32;
    exp_47_ram[578] = 101;
    exp_47_ram[579] = 101;
    exp_47_ram[580] = 46;
    exp_47_ram[581] = 0;
    exp_47_ram[582] = 10;
    exp_47_ram[583] = 32;
    exp_47_ram[584] = 98;
    exp_47_ram[585] = 105;
    exp_47_ram[586] = 103;
    exp_47_ram[587] = 109;
    exp_47_ram[588] = 105;
    exp_47_ram[589] = 101;
    exp_47_ram[590] = 110;
    exp_47_ram[591] = 115;
    exp_47_ram[592] = 110;
    exp_47_ram[593] = 0;
    exp_47_ram[594] = 32;
    exp_47_ram[595] = 98;
    exp_47_ram[596] = 105;
    exp_47_ram[597] = 103;
    exp_47_ram[598] = 109;
    exp_47_ram[599] = 105;
    exp_47_ram[600] = 101;
    exp_47_ram[601] = 110;
    exp_47_ram[602] = 115;
    exp_47_ram[603] = 110;
    exp_47_ram[604] = 0;
    exp_47_ram[605] = 32;
    exp_47_ram[606] = 98;
    exp_47_ram[607] = 105;
    exp_47_ram[608] = 103;
    exp_47_ram[609] = 100;
    exp_47_ram[610] = 100;
    exp_47_ram[611] = 105;
    exp_47_ram[612] = 32;
    exp_47_ram[613] = 111;
    exp_47_ram[614] = 0;
    exp_47_ram[615] = 32;
    exp_47_ram[616] = 98;
    exp_47_ram[617] = 105;
    exp_47_ram[618] = 103;
    exp_47_ram[619] = 100;
    exp_47_ram[620] = 100;
    exp_47_ram[621] = 105;
    exp_47_ram[622] = 32;
    exp_47_ram[623] = 111;
    exp_47_ram[624] = 0;
    exp_47_ram[625] = 97;
    exp_47_ram[626] = 0;
    exp_47_ram[627] = 110;
    exp_47_ram[628] = 10;
    exp_47_ram[629] = 121;
    exp_47_ram[630] = 0;
    exp_47_ram[631] = 117;
    exp_47_ram[632] = 0;
    exp_47_ram[633] = 110;
    exp_47_ram[634] = 58;
    exp_47_ram[635] = 0;
    exp_47_ram[636] = 104;
    exp_47_ram[637] = 45;
    exp_47_ram[638] = 101;
    exp_47_ram[639] = 0;
    exp_47_ram[640] = 41;
    exp_47_ram[641] = 108;
    exp_47_ram[642] = 87;
    exp_47_ram[643] = 100;
    exp_47_ram[644] = 0;
    exp_47_ram[645] = 32;
    exp_47_ram[646] = 103;
    exp_47_ram[647] = 82;
    exp_47_ram[648] = 114;
    exp_47_ram[649] = 0;
    exp_47_ram[650] = 32;
    exp_47_ram[651] = 116;
    exp_47_ram[652] = 108;
    exp_47_ram[653] = 108;
    exp_47_ram[654] = 116;
    exp_47_ram[655] = 10;
    exp_47_ram[656] = 32;
    exp_47_ram[657] = 108;
    exp_47_ram[658] = 111;
    exp_47_ram[659] = 0;
    exp_47_ram[660] = 2;
    exp_47_ram[661] = 3;
    exp_47_ram[662] = 4;
    exp_47_ram[663] = 4;
    exp_47_ram[664] = 5;
    exp_47_ram[665] = 5;
    exp_47_ram[666] = 5;
    exp_47_ram[667] = 5;
    exp_47_ram[668] = 6;
    exp_47_ram[669] = 6;
    exp_47_ram[670] = 6;
    exp_47_ram[671] = 6;
    exp_47_ram[672] = 6;
    exp_47_ram[673] = 6;
    exp_47_ram[674] = 6;
    exp_47_ram[675] = 6;
    exp_47_ram[676] = 7;
    exp_47_ram[677] = 7;
    exp_47_ram[678] = 7;
    exp_47_ram[679] = 7;
    exp_47_ram[680] = 7;
    exp_47_ram[681] = 7;
    exp_47_ram[682] = 7;
    exp_47_ram[683] = 7;
    exp_47_ram[684] = 7;
    exp_47_ram[685] = 7;
    exp_47_ram[686] = 7;
    exp_47_ram[687] = 7;
    exp_47_ram[688] = 7;
    exp_47_ram[689] = 7;
    exp_47_ram[690] = 7;
    exp_47_ram[691] = 7;
    exp_47_ram[692] = 8;
    exp_47_ram[693] = 8;
    exp_47_ram[694] = 8;
    exp_47_ram[695] = 8;
    exp_47_ram[696] = 8;
    exp_47_ram[697] = 8;
    exp_47_ram[698] = 8;
    exp_47_ram[699] = 8;
    exp_47_ram[700] = 8;
    exp_47_ram[701] = 8;
    exp_47_ram[702] = 8;
    exp_47_ram[703] = 8;
    exp_47_ram[704] = 8;
    exp_47_ram[705] = 8;
    exp_47_ram[706] = 8;
    exp_47_ram[707] = 8;
    exp_47_ram[708] = 8;
    exp_47_ram[709] = 8;
    exp_47_ram[710] = 8;
    exp_47_ram[711] = 8;
    exp_47_ram[712] = 8;
    exp_47_ram[713] = 8;
    exp_47_ram[714] = 8;
    exp_47_ram[715] = 8;
    exp_47_ram[716] = 8;
    exp_47_ram[717] = 8;
    exp_47_ram[718] = 8;
    exp_47_ram[719] = 8;
    exp_47_ram[720] = 8;
    exp_47_ram[721] = 8;
    exp_47_ram[722] = 8;
    exp_47_ram[723] = 8;
    exp_47_ram[724] = 1;
    exp_47_ram[725] = 129;
    exp_47_ram[726] = 1;
    exp_47_ram[727] = 164;
    exp_47_ram[728] = 196;
    exp_47_ram[729] = 244;
    exp_47_ram[730] = 196;
    exp_47_ram[731] = 7;
    exp_47_ram[732] = 7;
    exp_47_ram[733] = 193;
    exp_47_ram[734] = 1;
    exp_47_ram[735] = 0;
    exp_47_ram[736] = 1;
    exp_47_ram[737] = 129;
    exp_47_ram[738] = 1;
    exp_47_ram[739] = 164;
    exp_47_ram[740] = 180;
    exp_47_ram[741] = 132;
    exp_47_ram[742] = 244;
    exp_47_ram[743] = 196;
    exp_47_ram[744] = 196;
    exp_47_ram[745] = 231;
    exp_47_ram[746] = 196;
    exp_47_ram[747] = 7;
    exp_47_ram[748] = 193;
    exp_47_ram[749] = 1;
    exp_47_ram[750] = 0;
    exp_47_ram[751] = 1;
    exp_47_ram[752] = 17;
    exp_47_ram[753] = 129;
    exp_47_ram[754] = 1;
    exp_47_ram[755] = 0;
    exp_47_ram[756] = 199;
    exp_47_ram[757] = 7;
    exp_47_ram[758] = 159;
    exp_47_ram[759] = 5;
    exp_47_ram[760] = 7;
    exp_47_ram[761] = 193;
    exp_47_ram[762] = 129;
    exp_47_ram[763] = 1;
    exp_47_ram[764] = 0;
    exp_47_ram[765] = 1;
    exp_47_ram[766] = 17;
    exp_47_ram[767] = 129;
    exp_47_ram[768] = 1;
    exp_47_ram[769] = 164;
    exp_47_ram[770] = 180;
    exp_47_ram[771] = 4;
    exp_47_ram[772] = 128;
    exp_47_ram[773] = 196;
    exp_47_ram[774] = 23;
    exp_47_ram[775] = 228;
    exp_47_ram[776] = 196;
    exp_47_ram[777] = 247;
    exp_47_ram[778] = 7;
    exp_47_ram[779] = 132;
    exp_47_ram[780] = 7;
    exp_47_ram[781] = 223;
    exp_47_ram[782] = 196;
    exp_47_ram[783] = 196;
    exp_47_ram[784] = 247;
    exp_47_ram[785] = 7;
    exp_47_ram[786] = 7;
    exp_47_ram[787] = 196;
    exp_47_ram[788] = 7;
    exp_47_ram[789] = 193;
    exp_47_ram[790] = 129;
    exp_47_ram[791] = 1;
    exp_47_ram[792] = 0;
    exp_47_ram[793] = 1;
    exp_47_ram[794] = 17;
    exp_47_ram[795] = 129;
    exp_47_ram[796] = 1;
    exp_47_ram[797] = 164;
    exp_47_ram[798] = 0;
    exp_47_ram[799] = 71;
    exp_47_ram[800] = 7;
    exp_47_ram[801] = 196;
    exp_47_ram[802] = 223;
    exp_47_ram[803] = 0;
    exp_47_ram[804] = 71;
    exp_47_ram[805] = 7;
    exp_47_ram[806] = 160;
    exp_47_ram[807] = 95;
    exp_47_ram[808] = 0;
    exp_47_ram[809] = 7;
    exp_47_ram[810] = 193;
    exp_47_ram[811] = 129;
    exp_47_ram[812] = 1;
    exp_47_ram[813] = 0;
    exp_47_ram[814] = 1;
    exp_47_ram[815] = 129;
    exp_47_ram[816] = 1;
    exp_47_ram[817] = 5;
    exp_47_ram[818] = 180;
    exp_47_ram[819] = 196;
    exp_47_ram[820] = 212;
    exp_47_ram[821] = 244;
    exp_47_ram[822] = 0;
    exp_47_ram[823] = 193;
    exp_47_ram[824] = 1;
    exp_47_ram[825] = 0;
    exp_47_ram[826] = 1;
    exp_47_ram[827] = 17;
    exp_47_ram[828] = 129;
    exp_47_ram[829] = 1;
    exp_47_ram[830] = 5;
    exp_47_ram[831] = 180;
    exp_47_ram[832] = 196;
    exp_47_ram[833] = 212;
    exp_47_ram[834] = 244;
    exp_47_ram[835] = 244;
    exp_47_ram[836] = 7;
    exp_47_ram[837] = 244;
    exp_47_ram[838] = 7;
    exp_47_ram[839] = 192;
    exp_47_ram[840] = 0;
    exp_47_ram[841] = 193;
    exp_47_ram[842] = 129;
    exp_47_ram[843] = 1;
    exp_47_ram[844] = 0;
    exp_47_ram[845] = 1;
    exp_47_ram[846] = 129;
    exp_47_ram[847] = 1;
    exp_47_ram[848] = 164;
    exp_47_ram[849] = 180;
    exp_47_ram[850] = 196;
    exp_47_ram[851] = 244;
    exp_47_ram[852] = 0;
    exp_47_ram[853] = 196;
    exp_47_ram[854] = 23;
    exp_47_ram[855] = 244;
    exp_47_ram[856] = 196;
    exp_47_ram[857] = 7;
    exp_47_ram[858] = 7;
    exp_47_ram[859] = 132;
    exp_47_ram[860] = 247;
    exp_47_ram[861] = 228;
    exp_47_ram[862] = 7;
    exp_47_ram[863] = 196;
    exp_47_ram[864] = 196;
    exp_47_ram[865] = 247;
    exp_47_ram[866] = 7;
    exp_47_ram[867] = 193;
    exp_47_ram[868] = 1;
    exp_47_ram[869] = 0;
    exp_47_ram[870] = 1;
    exp_47_ram[871] = 129;
    exp_47_ram[872] = 1;
    exp_47_ram[873] = 5;
    exp_47_ram[874] = 244;
    exp_47_ram[875] = 244;
    exp_47_ram[876] = 240;
    exp_47_ram[877] = 231;
    exp_47_ram[878] = 244;
    exp_47_ram[879] = 144;
    exp_47_ram[880] = 231;
    exp_47_ram[881] = 16;
    exp_47_ram[882] = 128;
    exp_47_ram[883] = 0;
    exp_47_ram[884] = 23;
    exp_47_ram[885] = 247;
    exp_47_ram[886] = 7;
    exp_47_ram[887] = 193;
    exp_47_ram[888] = 1;
    exp_47_ram[889] = 0;
    exp_47_ram[890] = 1;
    exp_47_ram[891] = 17;
    exp_47_ram[892] = 129;
    exp_47_ram[893] = 1;
    exp_47_ram[894] = 164;
    exp_47_ram[895] = 4;
    exp_47_ram[896] = 0;
    exp_47_ram[897] = 196;
    exp_47_ram[898] = 7;
    exp_47_ram[899] = 39;
    exp_47_ram[900] = 231;
    exp_47_ram[901] = 23;
    exp_47_ram[902] = 7;
    exp_47_ram[903] = 196;
    exp_47_ram[904] = 7;
    exp_47_ram[905] = 23;
    exp_47_ram[906] = 196;
    exp_47_ram[907] = 215;
    exp_47_ram[908] = 7;
    exp_47_ram[909] = 246;
    exp_47_ram[910] = 7;
    exp_47_ram[911] = 244;
    exp_47_ram[912] = 196;
    exp_47_ram[913] = 7;
    exp_47_ram[914] = 7;
    exp_47_ram[915] = 7;
    exp_47_ram[916] = 159;
    exp_47_ram[917] = 5;
    exp_47_ram[918] = 7;
    exp_47_ram[919] = 196;
    exp_47_ram[920] = 7;
    exp_47_ram[921] = 193;
    exp_47_ram[922] = 129;
    exp_47_ram[923] = 1;
    exp_47_ram[924] = 0;
    exp_47_ram[925] = 1;
    exp_47_ram[926] = 17;
    exp_47_ram[927] = 129;
    exp_47_ram[928] = 1;
    exp_47_ram[929] = 164;
    exp_47_ram[930] = 180;
    exp_47_ram[931] = 196;
    exp_47_ram[932] = 212;
    exp_47_ram[933] = 228;
    exp_47_ram[934] = 244;
    exp_47_ram[935] = 4;
    exp_47_ram[936] = 20;
    exp_47_ram[937] = 68;
    exp_47_ram[938] = 244;
    exp_47_ram[939] = 4;
    exp_47_ram[940] = 39;
    exp_47_ram[941] = 7;
    exp_47_ram[942] = 4;
    exp_47_ram[943] = 23;
    exp_47_ram[944] = 7;
    exp_47_ram[945] = 132;
    exp_47_ram[946] = 244;
    exp_47_ram[947] = 64;
    exp_47_ram[948] = 68;
    exp_47_ram[949] = 23;
    exp_47_ram[950] = 228;
    exp_47_ram[951] = 196;
    exp_47_ram[952] = 4;
    exp_47_ram[953] = 7;
    exp_47_ram[954] = 132;
    exp_47_ram[955] = 0;
    exp_47_ram[956] = 7;
    exp_47_ram[957] = 196;
    exp_47_ram[958] = 23;
    exp_47_ram[959] = 244;
    exp_47_ram[960] = 196;
    exp_47_ram[961] = 68;
    exp_47_ram[962] = 247;
    exp_47_ram[963] = 0;
    exp_47_ram[964] = 132;
    exp_47_ram[965] = 247;
    exp_47_ram[966] = 244;
    exp_47_ram[967] = 196;
    exp_47_ram[968] = 132;
    exp_47_ram[969] = 247;
    exp_47_ram[970] = 7;
    exp_47_ram[971] = 68;
    exp_47_ram[972] = 23;
    exp_47_ram[973] = 228;
    exp_47_ram[974] = 196;
    exp_47_ram[975] = 4;
    exp_47_ram[976] = 7;
    exp_47_ram[977] = 132;
    exp_47_ram[978] = 7;
    exp_47_ram[979] = 132;
    exp_47_ram[980] = 7;
    exp_47_ram[981] = 4;
    exp_47_ram[982] = 39;
    exp_47_ram[983] = 7;
    exp_47_ram[984] = 128;
    exp_47_ram[985] = 68;
    exp_47_ram[986] = 23;
    exp_47_ram[987] = 228;
    exp_47_ram[988] = 196;
    exp_47_ram[989] = 4;
    exp_47_ram[990] = 7;
    exp_47_ram[991] = 132;
    exp_47_ram[992] = 0;
    exp_47_ram[993] = 7;
    exp_47_ram[994] = 68;
    exp_47_ram[995] = 132;
    exp_47_ram[996] = 247;
    exp_47_ram[997] = 68;
    exp_47_ram[998] = 231;
    exp_47_ram[999] = 68;
    exp_47_ram[1000] = 7;
    exp_47_ram[1001] = 193;
    exp_47_ram[1002] = 129;
    exp_47_ram[1003] = 1;
    exp_47_ram[1004] = 0;
    exp_47_ram[1005] = 1;
    exp_47_ram[1006] = 17;
    exp_47_ram[1007] = 129;
    exp_47_ram[1008] = 1;
    exp_47_ram[1009] = 164;
    exp_47_ram[1010] = 180;
    exp_47_ram[1011] = 196;
    exp_47_ram[1012] = 212;
    exp_47_ram[1013] = 228;
    exp_47_ram[1014] = 244;
    exp_47_ram[1015] = 8;
    exp_47_ram[1016] = 20;
    exp_47_ram[1017] = 244;
    exp_47_ram[1018] = 132;
    exp_47_ram[1019] = 39;
    exp_47_ram[1020] = 7;
    exp_47_ram[1021] = 68;
    exp_47_ram[1022] = 7;
    exp_47_ram[1023] = 132;
    exp_47_ram[1024] = 23;
    exp_47_ram[1025] = 7;
    exp_47_ram[1026] = 116;
    exp_47_ram[1027] = 7;
    exp_47_ram[1028] = 132;
    exp_47_ram[1029] = 199;
    exp_47_ram[1030] = 7;
    exp_47_ram[1031] = 68;
    exp_47_ram[1032] = 247;
    exp_47_ram[1033] = 244;
    exp_47_ram[1034] = 0;
    exp_47_ram[1035] = 132;
    exp_47_ram[1036] = 23;
    exp_47_ram[1037] = 228;
    exp_47_ram[1038] = 196;
    exp_47_ram[1039] = 247;
    exp_47_ram[1040] = 0;
    exp_47_ram[1041] = 231;
    exp_47_ram[1042] = 132;
    exp_47_ram[1043] = 4;
    exp_47_ram[1044] = 247;
    exp_47_ram[1045] = 132;
    exp_47_ram[1046] = 240;
    exp_47_ram[1047] = 231;
    exp_47_ram[1048] = 0;
    exp_47_ram[1049] = 132;
    exp_47_ram[1050] = 23;
    exp_47_ram[1051] = 228;
    exp_47_ram[1052] = 196;
    exp_47_ram[1053] = 247;
    exp_47_ram[1054] = 0;
    exp_47_ram[1055] = 231;
    exp_47_ram[1056] = 132;
    exp_47_ram[1057] = 23;
    exp_47_ram[1058] = 7;
    exp_47_ram[1059] = 132;
    exp_47_ram[1060] = 68;
    exp_47_ram[1061] = 247;
    exp_47_ram[1062] = 132;
    exp_47_ram[1063] = 240;
    exp_47_ram[1064] = 231;
    exp_47_ram[1065] = 132;
    exp_47_ram[1066] = 7;
    exp_47_ram[1067] = 7;
    exp_47_ram[1068] = 132;
    exp_47_ram[1069] = 7;
    exp_47_ram[1070] = 7;
    exp_47_ram[1071] = 132;
    exp_47_ram[1072] = 7;
    exp_47_ram[1073] = 132;
    exp_47_ram[1074] = 4;
    exp_47_ram[1075] = 247;
    exp_47_ram[1076] = 132;
    exp_47_ram[1077] = 68;
    exp_47_ram[1078] = 247;
    exp_47_ram[1079] = 132;
    exp_47_ram[1080] = 247;
    exp_47_ram[1081] = 244;
    exp_47_ram[1082] = 132;
    exp_47_ram[1083] = 7;
    exp_47_ram[1084] = 4;
    exp_47_ram[1085] = 0;
    exp_47_ram[1086] = 247;
    exp_47_ram[1087] = 132;
    exp_47_ram[1088] = 247;
    exp_47_ram[1089] = 244;
    exp_47_ram[1090] = 4;
    exp_47_ram[1091] = 0;
    exp_47_ram[1092] = 247;
    exp_47_ram[1093] = 132;
    exp_47_ram[1094] = 7;
    exp_47_ram[1095] = 7;
    exp_47_ram[1096] = 132;
    exp_47_ram[1097] = 240;
    exp_47_ram[1098] = 231;
    exp_47_ram[1099] = 132;
    exp_47_ram[1100] = 23;
    exp_47_ram[1101] = 228;
    exp_47_ram[1102] = 196;
    exp_47_ram[1103] = 247;
    exp_47_ram[1104] = 128;
    exp_47_ram[1105] = 231;
    exp_47_ram[1106] = 192;
    exp_47_ram[1107] = 4;
    exp_47_ram[1108] = 0;
    exp_47_ram[1109] = 247;
    exp_47_ram[1110] = 132;
    exp_47_ram[1111] = 7;
    exp_47_ram[1112] = 7;
    exp_47_ram[1113] = 132;
    exp_47_ram[1114] = 240;
    exp_47_ram[1115] = 231;
    exp_47_ram[1116] = 132;
    exp_47_ram[1117] = 23;
    exp_47_ram[1118] = 228;
    exp_47_ram[1119] = 196;
    exp_47_ram[1120] = 247;
    exp_47_ram[1121] = 128;
    exp_47_ram[1122] = 231;
    exp_47_ram[1123] = 128;
    exp_47_ram[1124] = 4;
    exp_47_ram[1125] = 32;
    exp_47_ram[1126] = 247;
    exp_47_ram[1127] = 132;
    exp_47_ram[1128] = 240;
    exp_47_ram[1129] = 231;
    exp_47_ram[1130] = 132;
    exp_47_ram[1131] = 23;
    exp_47_ram[1132] = 228;
    exp_47_ram[1133] = 196;
    exp_47_ram[1134] = 247;
    exp_47_ram[1135] = 32;
    exp_47_ram[1136] = 231;
    exp_47_ram[1137] = 132;
    exp_47_ram[1138] = 240;
    exp_47_ram[1139] = 231;
    exp_47_ram[1140] = 132;
    exp_47_ram[1141] = 23;
    exp_47_ram[1142] = 228;
    exp_47_ram[1143] = 196;
    exp_47_ram[1144] = 247;
    exp_47_ram[1145] = 0;
    exp_47_ram[1146] = 231;
    exp_47_ram[1147] = 132;
    exp_47_ram[1148] = 240;
    exp_47_ram[1149] = 231;
    exp_47_ram[1150] = 116;
    exp_47_ram[1151] = 7;
    exp_47_ram[1152] = 132;
    exp_47_ram[1153] = 23;
    exp_47_ram[1154] = 228;
    exp_47_ram[1155] = 196;
    exp_47_ram[1156] = 247;
    exp_47_ram[1157] = 208;
    exp_47_ram[1158] = 231;
    exp_47_ram[1159] = 128;
    exp_47_ram[1160] = 132;
    exp_47_ram[1161] = 71;
    exp_47_ram[1162] = 7;
    exp_47_ram[1163] = 132;
    exp_47_ram[1164] = 23;
    exp_47_ram[1165] = 228;
    exp_47_ram[1166] = 196;
    exp_47_ram[1167] = 247;
    exp_47_ram[1168] = 176;
    exp_47_ram[1169] = 231;
    exp_47_ram[1170] = 192;
    exp_47_ram[1171] = 132;
    exp_47_ram[1172] = 135;
    exp_47_ram[1173] = 7;
    exp_47_ram[1174] = 132;
    exp_47_ram[1175] = 23;
    exp_47_ram[1176] = 228;
    exp_47_ram[1177] = 196;
    exp_47_ram[1178] = 247;
    exp_47_ram[1179] = 0;
    exp_47_ram[1180] = 231;
    exp_47_ram[1181] = 132;
    exp_47_ram[1182] = 68;
    exp_47_ram[1183] = 132;
    exp_47_ram[1184] = 196;
    exp_47_ram[1185] = 4;
    exp_47_ram[1186] = 68;
    exp_47_ram[1187] = 132;
    exp_47_ram[1188] = 196;
    exp_47_ram[1189] = 31;
    exp_47_ram[1190] = 5;
    exp_47_ram[1191] = 7;
    exp_47_ram[1192] = 193;
    exp_47_ram[1193] = 129;
    exp_47_ram[1194] = 1;
    exp_47_ram[1195] = 0;
    exp_47_ram[1196] = 1;
    exp_47_ram[1197] = 17;
    exp_47_ram[1198] = 129;
    exp_47_ram[1199] = 1;
    exp_47_ram[1200] = 164;
    exp_47_ram[1201] = 180;
    exp_47_ram[1202] = 196;
    exp_47_ram[1203] = 212;
    exp_47_ram[1204] = 228;
    exp_47_ram[1205] = 4;
    exp_47_ram[1206] = 20;
    exp_47_ram[1207] = 244;
    exp_47_ram[1208] = 4;
    exp_47_ram[1209] = 196;
    exp_47_ram[1210] = 7;
    exp_47_ram[1211] = 68;
    exp_47_ram[1212] = 247;
    exp_47_ram[1213] = 244;
    exp_47_ram[1214] = 68;
    exp_47_ram[1215] = 7;
    exp_47_ram[1216] = 7;
    exp_47_ram[1217] = 196;
    exp_47_ram[1218] = 7;
    exp_47_ram[1219] = 196;
    exp_47_ram[1220] = 68;
    exp_47_ram[1221] = 247;
    exp_47_ram[1222] = 244;
    exp_47_ram[1223] = 180;
    exp_47_ram[1224] = 144;
    exp_47_ram[1225] = 231;
    exp_47_ram[1226] = 180;
    exp_47_ram[1227] = 7;
    exp_47_ram[1228] = 247;
    exp_47_ram[1229] = 0;
    exp_47_ram[1230] = 68;
    exp_47_ram[1231] = 7;
    exp_47_ram[1232] = 7;
    exp_47_ram[1233] = 16;
    exp_47_ram[1234] = 128;
    exp_47_ram[1235] = 16;
    exp_47_ram[1236] = 180;
    exp_47_ram[1237] = 231;
    exp_47_ram[1238] = 247;
    exp_47_ram[1239] = 103;
    exp_47_ram[1240] = 247;
    exp_47_ram[1241] = 196;
    exp_47_ram[1242] = 23;
    exp_47_ram[1243] = 212;
    exp_47_ram[1244] = 4;
    exp_47_ram[1245] = 230;
    exp_47_ram[1246] = 247;
    exp_47_ram[1247] = 196;
    exp_47_ram[1248] = 68;
    exp_47_ram[1249] = 247;
    exp_47_ram[1250] = 244;
    exp_47_ram[1251] = 196;
    exp_47_ram[1252] = 7;
    exp_47_ram[1253] = 196;
    exp_47_ram[1254] = 240;
    exp_47_ram[1255] = 231;
    exp_47_ram[1256] = 180;
    exp_47_ram[1257] = 132;
    exp_47_ram[1258] = 68;
    exp_47_ram[1259] = 241;
    exp_47_ram[1260] = 4;
    exp_47_ram[1261] = 241;
    exp_47_ram[1262] = 4;
    exp_47_ram[1263] = 241;
    exp_47_ram[1264] = 68;
    exp_47_ram[1265] = 6;
    exp_47_ram[1266] = 196;
    exp_47_ram[1267] = 4;
    exp_47_ram[1268] = 68;
    exp_47_ram[1269] = 132;
    exp_47_ram[1270] = 196;
    exp_47_ram[1271] = 159;
    exp_47_ram[1272] = 5;
    exp_47_ram[1273] = 7;
    exp_47_ram[1274] = 193;
    exp_47_ram[1275] = 129;
    exp_47_ram[1276] = 1;
    exp_47_ram[1277] = 0;
    exp_47_ram[1278] = 1;
    exp_47_ram[1279] = 17;
    exp_47_ram[1280] = 129;
    exp_47_ram[1281] = 1;
    exp_47_ram[1282] = 164;
    exp_47_ram[1283] = 180;
    exp_47_ram[1284] = 196;
    exp_47_ram[1285] = 212;
    exp_47_ram[1286] = 228;
    exp_47_ram[1287] = 4;
    exp_47_ram[1288] = 132;
    exp_47_ram[1289] = 7;
    exp_47_ram[1290] = 0;
    exp_47_ram[1291] = 135;
    exp_47_ram[1292] = 244;
    exp_47_ram[1293] = 208;
    exp_47_ram[1294] = 4;
    exp_47_ram[1295] = 7;
    exp_47_ram[1296] = 80;
    exp_47_ram[1297] = 247;
    exp_47_ram[1298] = 4;
    exp_47_ram[1299] = 7;
    exp_47_ram[1300] = 196;
    exp_47_ram[1301] = 23;
    exp_47_ram[1302] = 228;
    exp_47_ram[1303] = 196;
    exp_47_ram[1304] = 68;
    exp_47_ram[1305] = 7;
    exp_47_ram[1306] = 132;
    exp_47_ram[1307] = 7;
    exp_47_ram[1308] = 4;
    exp_47_ram[1309] = 23;
    exp_47_ram[1310] = 244;
    exp_47_ram[1311] = 80;
    exp_47_ram[1312] = 4;
    exp_47_ram[1313] = 23;
    exp_47_ram[1314] = 244;
    exp_47_ram[1315] = 4;
    exp_47_ram[1316] = 4;
    exp_47_ram[1317] = 7;
    exp_47_ram[1318] = 7;
    exp_47_ram[1319] = 0;
    exp_47_ram[1320] = 247;
    exp_47_ram[1321] = 39;
    exp_47_ram[1322] = 0;
    exp_47_ram[1323] = 7;
    exp_47_ram[1324] = 247;
    exp_47_ram[1325] = 7;
    exp_47_ram[1326] = 7;
    exp_47_ram[1327] = 196;
    exp_47_ram[1328] = 23;
    exp_47_ram[1329] = 244;
    exp_47_ram[1330] = 4;
    exp_47_ram[1331] = 23;
    exp_47_ram[1332] = 244;
    exp_47_ram[1333] = 16;
    exp_47_ram[1334] = 244;
    exp_47_ram[1335] = 192;
    exp_47_ram[1336] = 196;
    exp_47_ram[1337] = 39;
    exp_47_ram[1338] = 244;
    exp_47_ram[1339] = 4;
    exp_47_ram[1340] = 23;
    exp_47_ram[1341] = 244;
    exp_47_ram[1342] = 16;
    exp_47_ram[1343] = 244;
    exp_47_ram[1344] = 128;
    exp_47_ram[1345] = 196;
    exp_47_ram[1346] = 71;
    exp_47_ram[1347] = 244;
    exp_47_ram[1348] = 4;
    exp_47_ram[1349] = 23;
    exp_47_ram[1350] = 244;
    exp_47_ram[1351] = 16;
    exp_47_ram[1352] = 244;
    exp_47_ram[1353] = 64;
    exp_47_ram[1354] = 196;
    exp_47_ram[1355] = 135;
    exp_47_ram[1356] = 244;
    exp_47_ram[1357] = 4;
    exp_47_ram[1358] = 23;
    exp_47_ram[1359] = 244;
    exp_47_ram[1360] = 16;
    exp_47_ram[1361] = 244;
    exp_47_ram[1362] = 0;
    exp_47_ram[1363] = 196;
    exp_47_ram[1364] = 7;
    exp_47_ram[1365] = 244;
    exp_47_ram[1366] = 4;
    exp_47_ram[1367] = 23;
    exp_47_ram[1368] = 244;
    exp_47_ram[1369] = 16;
    exp_47_ram[1370] = 244;
    exp_47_ram[1371] = 192;
    exp_47_ram[1372] = 4;
    exp_47_ram[1373] = 0;
    exp_47_ram[1374] = 4;
    exp_47_ram[1375] = 7;
    exp_47_ram[1376] = 4;
    exp_47_ram[1377] = 4;
    exp_47_ram[1378] = 7;
    exp_47_ram[1379] = 7;
    exp_47_ram[1380] = 159;
    exp_47_ram[1381] = 5;
    exp_47_ram[1382] = 7;
    exp_47_ram[1383] = 4;
    exp_47_ram[1384] = 7;
    exp_47_ram[1385] = 95;
    exp_47_ram[1386] = 164;
    exp_47_ram[1387] = 0;
    exp_47_ram[1388] = 4;
    exp_47_ram[1389] = 7;
    exp_47_ram[1390] = 160;
    exp_47_ram[1391] = 247;
    exp_47_ram[1392] = 196;
    exp_47_ram[1393] = 71;
    exp_47_ram[1394] = 228;
    exp_47_ram[1395] = 7;
    exp_47_ram[1396] = 244;
    exp_47_ram[1397] = 132;
    exp_47_ram[1398] = 7;
    exp_47_ram[1399] = 196;
    exp_47_ram[1400] = 39;
    exp_47_ram[1401] = 244;
    exp_47_ram[1402] = 132;
    exp_47_ram[1403] = 240;
    exp_47_ram[1404] = 244;
    exp_47_ram[1405] = 192;
    exp_47_ram[1406] = 132;
    exp_47_ram[1407] = 244;
    exp_47_ram[1408] = 4;
    exp_47_ram[1409] = 23;
    exp_47_ram[1410] = 244;
    exp_47_ram[1411] = 4;
    exp_47_ram[1412] = 4;
    exp_47_ram[1413] = 7;
    exp_47_ram[1414] = 224;
    exp_47_ram[1415] = 247;
    exp_47_ram[1416] = 196;
    exp_47_ram[1417] = 7;
    exp_47_ram[1418] = 244;
    exp_47_ram[1419] = 4;
    exp_47_ram[1420] = 23;
    exp_47_ram[1421] = 244;
    exp_47_ram[1422] = 4;
    exp_47_ram[1423] = 7;
    exp_47_ram[1424] = 7;
    exp_47_ram[1425] = 79;
    exp_47_ram[1426] = 5;
    exp_47_ram[1427] = 7;
    exp_47_ram[1428] = 4;
    exp_47_ram[1429] = 7;
    exp_47_ram[1430] = 15;
    exp_47_ram[1431] = 164;
    exp_47_ram[1432] = 64;
    exp_47_ram[1433] = 4;
    exp_47_ram[1434] = 7;
    exp_47_ram[1435] = 160;
    exp_47_ram[1436] = 247;
    exp_47_ram[1437] = 196;
    exp_47_ram[1438] = 71;
    exp_47_ram[1439] = 228;
    exp_47_ram[1440] = 7;
    exp_47_ram[1441] = 244;
    exp_47_ram[1442] = 68;
    exp_47_ram[1443] = 7;
    exp_47_ram[1444] = 0;
    exp_47_ram[1445] = 244;
    exp_47_ram[1446] = 4;
    exp_47_ram[1447] = 23;
    exp_47_ram[1448] = 244;
    exp_47_ram[1449] = 4;
    exp_47_ram[1450] = 7;
    exp_47_ram[1451] = 135;
    exp_47_ram[1452] = 32;
    exp_47_ram[1453] = 247;
    exp_47_ram[1454] = 39;
    exp_47_ram[1455] = 0;
    exp_47_ram[1456] = 71;
    exp_47_ram[1457] = 247;
    exp_47_ram[1458] = 7;
    exp_47_ram[1459] = 7;
    exp_47_ram[1460] = 196;
    exp_47_ram[1461] = 7;
    exp_47_ram[1462] = 244;
    exp_47_ram[1463] = 4;
    exp_47_ram[1464] = 23;
    exp_47_ram[1465] = 244;
    exp_47_ram[1466] = 4;
    exp_47_ram[1467] = 7;
    exp_47_ram[1468] = 192;
    exp_47_ram[1469] = 247;
    exp_47_ram[1470] = 196;
    exp_47_ram[1471] = 7;
    exp_47_ram[1472] = 244;
    exp_47_ram[1473] = 4;
    exp_47_ram[1474] = 23;
    exp_47_ram[1475] = 244;
    exp_47_ram[1476] = 64;
    exp_47_ram[1477] = 196;
    exp_47_ram[1478] = 7;
    exp_47_ram[1479] = 244;
    exp_47_ram[1480] = 4;
    exp_47_ram[1481] = 23;
    exp_47_ram[1482] = 244;
    exp_47_ram[1483] = 4;
    exp_47_ram[1484] = 7;
    exp_47_ram[1485] = 128;
    exp_47_ram[1486] = 247;
    exp_47_ram[1487] = 196;
    exp_47_ram[1488] = 7;
    exp_47_ram[1489] = 244;
    exp_47_ram[1490] = 4;
    exp_47_ram[1491] = 23;
    exp_47_ram[1492] = 244;
    exp_47_ram[1493] = 128;
    exp_47_ram[1494] = 196;
    exp_47_ram[1495] = 7;
    exp_47_ram[1496] = 244;
    exp_47_ram[1497] = 4;
    exp_47_ram[1498] = 23;
    exp_47_ram[1499] = 244;
    exp_47_ram[1500] = 0;
    exp_47_ram[1501] = 196;
    exp_47_ram[1502] = 7;
    exp_47_ram[1503] = 244;
    exp_47_ram[1504] = 4;
    exp_47_ram[1505] = 23;
    exp_47_ram[1506] = 244;
    exp_47_ram[1507] = 64;
    exp_47_ram[1508] = 196;
    exp_47_ram[1509] = 7;
    exp_47_ram[1510] = 244;
    exp_47_ram[1511] = 4;
    exp_47_ram[1512] = 23;
    exp_47_ram[1513] = 244;
    exp_47_ram[1514] = 128;
    exp_47_ram[1515] = 0;
    exp_47_ram[1516] = 0;
    exp_47_ram[1517] = 0;
    exp_47_ram[1518] = 128;
    exp_47_ram[1519] = 0;
    exp_47_ram[1520] = 4;
    exp_47_ram[1521] = 7;
    exp_47_ram[1522] = 183;
    exp_47_ram[1523] = 48;
    exp_47_ram[1524] = 247;
    exp_47_ram[1525] = 39;
    exp_47_ram[1526] = 0;
    exp_47_ram[1527] = 7;
    exp_47_ram[1528] = 247;
    exp_47_ram[1529] = 7;
    exp_47_ram[1530] = 7;
    exp_47_ram[1531] = 4;
    exp_47_ram[1532] = 7;
    exp_47_ram[1533] = 128;
    exp_47_ram[1534] = 247;
    exp_47_ram[1535] = 4;
    exp_47_ram[1536] = 7;
    exp_47_ram[1537] = 128;
    exp_47_ram[1538] = 247;
    exp_47_ram[1539] = 0;
    exp_47_ram[1540] = 244;
    exp_47_ram[1541] = 0;
    exp_47_ram[1542] = 4;
    exp_47_ram[1543] = 7;
    exp_47_ram[1544] = 240;
    exp_47_ram[1545] = 247;
    exp_47_ram[1546] = 128;
    exp_47_ram[1547] = 244;
    exp_47_ram[1548] = 64;
    exp_47_ram[1549] = 4;
    exp_47_ram[1550] = 7;
    exp_47_ram[1551] = 32;
    exp_47_ram[1552] = 247;
    exp_47_ram[1553] = 32;
    exp_47_ram[1554] = 244;
    exp_47_ram[1555] = 128;
    exp_47_ram[1556] = 160;
    exp_47_ram[1557] = 244;
    exp_47_ram[1558] = 196;
    exp_47_ram[1559] = 247;
    exp_47_ram[1560] = 244;
    exp_47_ram[1561] = 4;
    exp_47_ram[1562] = 7;
    exp_47_ram[1563] = 128;
    exp_47_ram[1564] = 247;
    exp_47_ram[1565] = 196;
    exp_47_ram[1566] = 7;
    exp_47_ram[1567] = 244;
    exp_47_ram[1568] = 4;
    exp_47_ram[1569] = 7;
    exp_47_ram[1570] = 144;
    exp_47_ram[1571] = 247;
    exp_47_ram[1572] = 4;
    exp_47_ram[1573] = 7;
    exp_47_ram[1574] = 64;
    exp_47_ram[1575] = 247;
    exp_47_ram[1576] = 196;
    exp_47_ram[1577] = 55;
    exp_47_ram[1578] = 244;
    exp_47_ram[1579] = 196;
    exp_47_ram[1580] = 7;
    exp_47_ram[1581] = 7;
    exp_47_ram[1582] = 196;
    exp_47_ram[1583] = 231;
    exp_47_ram[1584] = 244;
    exp_47_ram[1585] = 4;
    exp_47_ram[1586] = 7;
    exp_47_ram[1587] = 144;
    exp_47_ram[1588] = 247;
    exp_47_ram[1589] = 4;
    exp_47_ram[1590] = 7;
    exp_47_ram[1591] = 64;
    exp_47_ram[1592] = 247;
    exp_47_ram[1593] = 196;
    exp_47_ram[1594] = 7;
    exp_47_ram[1595] = 7;
    exp_47_ram[1596] = 196;
    exp_47_ram[1597] = 7;
    exp_47_ram[1598] = 7;
    exp_47_ram[1599] = 196;
    exp_47_ram[1600] = 71;
    exp_47_ram[1601] = 228;
    exp_47_ram[1602] = 7;
    exp_47_ram[1603] = 244;
    exp_47_ram[1604] = 132;
    exp_47_ram[1605] = 247;
    exp_47_ram[1606] = 132;
    exp_47_ram[1607] = 247;
    exp_47_ram[1608] = 231;
    exp_47_ram[1609] = 7;
    exp_47_ram[1610] = 132;
    exp_47_ram[1611] = 247;
    exp_47_ram[1612] = 247;
    exp_47_ram[1613] = 196;
    exp_47_ram[1614] = 241;
    exp_47_ram[1615] = 132;
    exp_47_ram[1616] = 241;
    exp_47_ram[1617] = 68;
    exp_47_ram[1618] = 132;
    exp_47_ram[1619] = 7;
    exp_47_ram[1620] = 6;
    exp_47_ram[1621] = 68;
    exp_47_ram[1622] = 196;
    exp_47_ram[1623] = 132;
    exp_47_ram[1624] = 196;
    exp_47_ram[1625] = 223;
    exp_47_ram[1626] = 164;
    exp_47_ram[1627] = 192;
    exp_47_ram[1628] = 196;
    exp_47_ram[1629] = 7;
    exp_47_ram[1630] = 7;
    exp_47_ram[1631] = 196;
    exp_47_ram[1632] = 71;
    exp_47_ram[1633] = 228;
    exp_47_ram[1634] = 7;
    exp_47_ram[1635] = 247;
    exp_47_ram[1636] = 192;
    exp_47_ram[1637] = 196;
    exp_47_ram[1638] = 7;
    exp_47_ram[1639] = 7;
    exp_47_ram[1640] = 196;
    exp_47_ram[1641] = 71;
    exp_47_ram[1642] = 228;
    exp_47_ram[1643] = 7;
    exp_47_ram[1644] = 7;
    exp_47_ram[1645] = 7;
    exp_47_ram[1646] = 64;
    exp_47_ram[1647] = 196;
    exp_47_ram[1648] = 71;
    exp_47_ram[1649] = 228;
    exp_47_ram[1650] = 7;
    exp_47_ram[1651] = 244;
    exp_47_ram[1652] = 196;
    exp_47_ram[1653] = 247;
    exp_47_ram[1654] = 196;
    exp_47_ram[1655] = 247;
    exp_47_ram[1656] = 231;
    exp_47_ram[1657] = 7;
    exp_47_ram[1658] = 196;
    exp_47_ram[1659] = 247;
    exp_47_ram[1660] = 247;
    exp_47_ram[1661] = 196;
    exp_47_ram[1662] = 241;
    exp_47_ram[1663] = 132;
    exp_47_ram[1664] = 241;
    exp_47_ram[1665] = 68;
    exp_47_ram[1666] = 132;
    exp_47_ram[1667] = 7;
    exp_47_ram[1668] = 6;
    exp_47_ram[1669] = 68;
    exp_47_ram[1670] = 196;
    exp_47_ram[1671] = 132;
    exp_47_ram[1672] = 196;
    exp_47_ram[1673] = 223;
    exp_47_ram[1674] = 164;
    exp_47_ram[1675] = 192;
    exp_47_ram[1676] = 196;
    exp_47_ram[1677] = 7;
    exp_47_ram[1678] = 7;
    exp_47_ram[1679] = 196;
    exp_47_ram[1680] = 7;
    exp_47_ram[1681] = 7;
    exp_47_ram[1682] = 196;
    exp_47_ram[1683] = 71;
    exp_47_ram[1684] = 228;
    exp_47_ram[1685] = 7;
    exp_47_ram[1686] = 196;
    exp_47_ram[1687] = 241;
    exp_47_ram[1688] = 132;
    exp_47_ram[1689] = 241;
    exp_47_ram[1690] = 68;
    exp_47_ram[1691] = 132;
    exp_47_ram[1692] = 0;
    exp_47_ram[1693] = 68;
    exp_47_ram[1694] = 196;
    exp_47_ram[1695] = 132;
    exp_47_ram[1696] = 196;
    exp_47_ram[1697] = 223;
    exp_47_ram[1698] = 164;
    exp_47_ram[1699] = 192;
    exp_47_ram[1700] = 196;
    exp_47_ram[1701] = 7;
    exp_47_ram[1702] = 7;
    exp_47_ram[1703] = 196;
    exp_47_ram[1704] = 71;
    exp_47_ram[1705] = 228;
    exp_47_ram[1706] = 7;
    exp_47_ram[1707] = 247;
    exp_47_ram[1708] = 192;
    exp_47_ram[1709] = 196;
    exp_47_ram[1710] = 7;
    exp_47_ram[1711] = 7;
    exp_47_ram[1712] = 196;
    exp_47_ram[1713] = 71;
    exp_47_ram[1714] = 228;
    exp_47_ram[1715] = 7;
    exp_47_ram[1716] = 7;
    exp_47_ram[1717] = 7;
    exp_47_ram[1718] = 64;
    exp_47_ram[1719] = 196;
    exp_47_ram[1720] = 71;
    exp_47_ram[1721] = 228;
    exp_47_ram[1722] = 7;
    exp_47_ram[1723] = 244;
    exp_47_ram[1724] = 196;
    exp_47_ram[1725] = 241;
    exp_47_ram[1726] = 132;
    exp_47_ram[1727] = 241;
    exp_47_ram[1728] = 68;
    exp_47_ram[1729] = 132;
    exp_47_ram[1730] = 0;
    exp_47_ram[1731] = 4;
    exp_47_ram[1732] = 68;
    exp_47_ram[1733] = 196;
    exp_47_ram[1734] = 132;
    exp_47_ram[1735] = 196;
    exp_47_ram[1736] = 15;
    exp_47_ram[1737] = 164;
    exp_47_ram[1738] = 4;
    exp_47_ram[1739] = 23;
    exp_47_ram[1740] = 244;
    exp_47_ram[1741] = 192;
    exp_47_ram[1742] = 16;
    exp_47_ram[1743] = 244;
    exp_47_ram[1744] = 196;
    exp_47_ram[1745] = 39;
    exp_47_ram[1746] = 7;
    exp_47_ram[1747] = 128;
    exp_47_ram[1748] = 196;
    exp_47_ram[1749] = 23;
    exp_47_ram[1750] = 228;
    exp_47_ram[1751] = 196;
    exp_47_ram[1752] = 68;
    exp_47_ram[1753] = 7;
    exp_47_ram[1754] = 132;
    exp_47_ram[1755] = 0;
    exp_47_ram[1756] = 7;
    exp_47_ram[1757] = 68;
    exp_47_ram[1758] = 23;
    exp_47_ram[1759] = 228;
    exp_47_ram[1760] = 132;
    exp_47_ram[1761] = 231;
    exp_47_ram[1762] = 196;
    exp_47_ram[1763] = 71;
    exp_47_ram[1764] = 228;
    exp_47_ram[1765] = 7;
    exp_47_ram[1766] = 247;
    exp_47_ram[1767] = 196;
    exp_47_ram[1768] = 23;
    exp_47_ram[1769] = 228;
    exp_47_ram[1770] = 196;
    exp_47_ram[1771] = 68;
    exp_47_ram[1772] = 7;
    exp_47_ram[1773] = 132;
    exp_47_ram[1774] = 7;
    exp_47_ram[1775] = 196;
    exp_47_ram[1776] = 39;
    exp_47_ram[1777] = 7;
    exp_47_ram[1778] = 128;
    exp_47_ram[1779] = 196;
    exp_47_ram[1780] = 23;
    exp_47_ram[1781] = 228;
    exp_47_ram[1782] = 196;
    exp_47_ram[1783] = 68;
    exp_47_ram[1784] = 7;
    exp_47_ram[1785] = 132;
    exp_47_ram[1786] = 0;
    exp_47_ram[1787] = 7;
    exp_47_ram[1788] = 68;
    exp_47_ram[1789] = 23;
    exp_47_ram[1790] = 228;
    exp_47_ram[1791] = 132;
    exp_47_ram[1792] = 231;
    exp_47_ram[1793] = 4;
    exp_47_ram[1794] = 23;
    exp_47_ram[1795] = 244;
    exp_47_ram[1796] = 0;
    exp_47_ram[1797] = 196;
    exp_47_ram[1798] = 71;
    exp_47_ram[1799] = 228;
    exp_47_ram[1800] = 7;
    exp_47_ram[1801] = 244;
    exp_47_ram[1802] = 68;
    exp_47_ram[1803] = 7;
    exp_47_ram[1804] = 68;
    exp_47_ram[1805] = 128;
    exp_47_ram[1806] = 240;
    exp_47_ram[1807] = 7;
    exp_47_ram[1808] = 4;
    exp_47_ram[1809] = 15;
    exp_47_ram[1810] = 164;
    exp_47_ram[1811] = 196;
    exp_47_ram[1812] = 7;
    exp_47_ram[1813] = 7;
    exp_47_ram[1814] = 196;
    exp_47_ram[1815] = 68;
    exp_47_ram[1816] = 247;
    exp_47_ram[1817] = 7;
    exp_47_ram[1818] = 244;
    exp_47_ram[1819] = 196;
    exp_47_ram[1820] = 39;
    exp_47_ram[1821] = 7;
    exp_47_ram[1822] = 128;
    exp_47_ram[1823] = 196;
    exp_47_ram[1824] = 23;
    exp_47_ram[1825] = 228;
    exp_47_ram[1826] = 196;
    exp_47_ram[1827] = 68;
    exp_47_ram[1828] = 7;
    exp_47_ram[1829] = 132;
    exp_47_ram[1830] = 0;
    exp_47_ram[1831] = 7;
    exp_47_ram[1832] = 196;
    exp_47_ram[1833] = 23;
    exp_47_ram[1834] = 228;
    exp_47_ram[1835] = 132;
    exp_47_ram[1836] = 231;
    exp_47_ram[1837] = 64;
    exp_47_ram[1838] = 4;
    exp_47_ram[1839] = 23;
    exp_47_ram[1840] = 228;
    exp_47_ram[1841] = 7;
    exp_47_ram[1842] = 196;
    exp_47_ram[1843] = 23;
    exp_47_ram[1844] = 228;
    exp_47_ram[1845] = 196;
    exp_47_ram[1846] = 68;
    exp_47_ram[1847] = 7;
    exp_47_ram[1848] = 132;
    exp_47_ram[1849] = 7;
    exp_47_ram[1850] = 4;
    exp_47_ram[1851] = 7;
    exp_47_ram[1852] = 7;
    exp_47_ram[1853] = 196;
    exp_47_ram[1854] = 7;
    exp_47_ram[1855] = 7;
    exp_47_ram[1856] = 68;
    exp_47_ram[1857] = 247;
    exp_47_ram[1858] = 228;
    exp_47_ram[1859] = 7;
    exp_47_ram[1860] = 196;
    exp_47_ram[1861] = 39;
    exp_47_ram[1862] = 7;
    exp_47_ram[1863] = 128;
    exp_47_ram[1864] = 196;
    exp_47_ram[1865] = 23;
    exp_47_ram[1866] = 228;
    exp_47_ram[1867] = 196;
    exp_47_ram[1868] = 68;
    exp_47_ram[1869] = 7;
    exp_47_ram[1870] = 132;
    exp_47_ram[1871] = 0;
    exp_47_ram[1872] = 7;
    exp_47_ram[1873] = 196;
    exp_47_ram[1874] = 23;
    exp_47_ram[1875] = 228;
    exp_47_ram[1876] = 132;
    exp_47_ram[1877] = 231;
    exp_47_ram[1878] = 4;
    exp_47_ram[1879] = 23;
    exp_47_ram[1880] = 244;
    exp_47_ram[1881] = 192;
    exp_47_ram[1882] = 128;
    exp_47_ram[1883] = 244;
    exp_47_ram[1884] = 196;
    exp_47_ram[1885] = 23;
    exp_47_ram[1886] = 244;
    exp_47_ram[1887] = 196;
    exp_47_ram[1888] = 71;
    exp_47_ram[1889] = 228;
    exp_47_ram[1890] = 7;
    exp_47_ram[1891] = 7;
    exp_47_ram[1892] = 196;
    exp_47_ram[1893] = 241;
    exp_47_ram[1894] = 132;
    exp_47_ram[1895] = 241;
    exp_47_ram[1896] = 68;
    exp_47_ram[1897] = 0;
    exp_47_ram[1898] = 0;
    exp_47_ram[1899] = 68;
    exp_47_ram[1900] = 196;
    exp_47_ram[1901] = 132;
    exp_47_ram[1902] = 196;
    exp_47_ram[1903] = 79;
    exp_47_ram[1904] = 164;
    exp_47_ram[1905] = 4;
    exp_47_ram[1906] = 23;
    exp_47_ram[1907] = 244;
    exp_47_ram[1908] = 0;
    exp_47_ram[1909] = 196;
    exp_47_ram[1910] = 23;
    exp_47_ram[1911] = 228;
    exp_47_ram[1912] = 196;
    exp_47_ram[1913] = 68;
    exp_47_ram[1914] = 7;
    exp_47_ram[1915] = 132;
    exp_47_ram[1916] = 80;
    exp_47_ram[1917] = 7;
    exp_47_ram[1918] = 4;
    exp_47_ram[1919] = 23;
    exp_47_ram[1920] = 244;
    exp_47_ram[1921] = 192;
    exp_47_ram[1922] = 4;
    exp_47_ram[1923] = 7;
    exp_47_ram[1924] = 196;
    exp_47_ram[1925] = 23;
    exp_47_ram[1926] = 228;
    exp_47_ram[1927] = 196;
    exp_47_ram[1928] = 68;
    exp_47_ram[1929] = 7;
    exp_47_ram[1930] = 132;
    exp_47_ram[1931] = 7;
    exp_47_ram[1932] = 4;
    exp_47_ram[1933] = 23;
    exp_47_ram[1934] = 244;
    exp_47_ram[1935] = 0;
    exp_47_ram[1936] = 4;
    exp_47_ram[1937] = 7;
    exp_47_ram[1938] = 7;
    exp_47_ram[1939] = 196;
    exp_47_ram[1940] = 68;
    exp_47_ram[1941] = 247;
    exp_47_ram[1942] = 68;
    exp_47_ram[1943] = 247;
    exp_47_ram[1944] = 128;
    exp_47_ram[1945] = 196;
    exp_47_ram[1946] = 196;
    exp_47_ram[1947] = 68;
    exp_47_ram[1948] = 7;
    exp_47_ram[1949] = 132;
    exp_47_ram[1950] = 0;
    exp_47_ram[1951] = 7;
    exp_47_ram[1952] = 196;
    exp_47_ram[1953] = 7;
    exp_47_ram[1954] = 193;
    exp_47_ram[1955] = 129;
    exp_47_ram[1956] = 1;
    exp_47_ram[1957] = 0;
    exp_47_ram[1958] = 1;
    exp_47_ram[1959] = 17;
    exp_47_ram[1960] = 129;
    exp_47_ram[1961] = 1;
    exp_47_ram[1962] = 164;
    exp_47_ram[1963] = 180;
    exp_47_ram[1964] = 196;
    exp_47_ram[1965] = 212;
    exp_47_ram[1966] = 228;
    exp_47_ram[1967] = 244;
    exp_47_ram[1968] = 4;
    exp_47_ram[1969] = 20;
    exp_47_ram[1970] = 4;
    exp_47_ram[1971] = 244;
    exp_47_ram[1972] = 132;
    exp_47_ram[1973] = 71;
    exp_47_ram[1974] = 244;
    exp_47_ram[1975] = 132;
    exp_47_ram[1976] = 68;
    exp_47_ram[1977] = 196;
    exp_47_ram[1978] = 240;
    exp_47_ram[1979] = 7;
    exp_47_ram[1980] = 0;
    exp_47_ram[1981] = 135;
    exp_47_ram[1982] = 15;
    exp_47_ram[1983] = 164;
    exp_47_ram[1984] = 196;
    exp_47_ram[1985] = 7;
    exp_47_ram[1986] = 193;
    exp_47_ram[1987] = 129;
    exp_47_ram[1988] = 1;
    exp_47_ram[1989] = 0;
    exp_47_ram[1990] = 1;
    exp_47_ram[1991] = 17;
    exp_47_ram[1992] = 129;
    exp_47_ram[1993] = 1;
    exp_47_ram[1994] = 5;
    exp_47_ram[1995] = 244;
    exp_47_ram[1996] = 244;
    exp_47_ram[1997] = 0;
    exp_47_ram[1998] = 71;
    exp_47_ram[1999] = 7;
    exp_47_ram[2000] = 7;
    exp_47_ram[2001] = 223;
    exp_47_ram[2002] = 0;
    exp_47_ram[2003] = 193;
    exp_47_ram[2004] = 129;
    exp_47_ram[2005] = 1;
    exp_47_ram[2006] = 0;
    exp_47_ram[2007] = 1;
    exp_47_ram[2008] = 17;
    exp_47_ram[2009] = 129;
    exp_47_ram[2010] = 145;
    exp_47_ram[2011] = 1;
    exp_47_ram[2012] = 5;
    exp_47_ram[2013] = 68;
    exp_47_ram[2014] = 244;
    exp_47_ram[2015] = 144;
    exp_47_ram[2016] = 244;
    exp_47_ram[2017] = 240;
    exp_47_ram[2018] = 244;
    exp_47_ram[2019] = 16;
    exp_47_ram[2020] = 244;
    exp_47_ram[2021] = 4;
    exp_47_ram[2022] = 4;
    exp_47_ram[2023] = 4;
    exp_47_ram[2024] = 68;
    exp_47_ram[2025] = 132;
    exp_47_ram[2026] = 196;
    exp_47_ram[2027] = 4;
    exp_47_ram[2028] = 68;
    exp_47_ram[2029] = 132;
    exp_47_ram[2030] = 196;
    exp_47_ram[2031] = 4;
    exp_47_ram[2032] = 68;
    exp_47_ram[2033] = 100;
    exp_47_ram[2034] = 20;
    exp_47_ram[2035] = 4;
    exp_47_ram[2036] = 164;
    exp_47_ram[2037] = 180;
    exp_47_ram[2038] = 196;
    exp_47_ram[2039] = 212;
    exp_47_ram[2040] = 228;
    exp_47_ram[2041] = 244;
    exp_47_ram[2042] = 4;
    exp_47_ram[2043] = 7;
    exp_47_ram[2044] = 64;
    exp_47_ram[2045] = 164;
    exp_47_ram[2046] = 180;
    exp_47_ram[2047] = 68;
    exp_47_ram[2048] = 132;
    exp_47_ram[2049] = 196;
    exp_47_ram[2050] = 7;
    exp_47_ram[2051] = 0;
    exp_47_ram[2052] = 4;
    exp_47_ram[2053] = 196;
    exp_47_ram[2054] = 247;
    exp_47_ram[2055] = 244;
    exp_47_ram[2056] = 68;
    exp_47_ram[2057] = 132;
    exp_47_ram[2058] = 196;
    exp_47_ram[2059] = 4;
    exp_47_ram[2060] = 68;
    exp_47_ram[2061] = 132;
    exp_47_ram[2062] = 196;
    exp_47_ram[2063] = 4;
    exp_47_ram[2064] = 68;
    exp_47_ram[2065] = 100;
    exp_47_ram[2066] = 20;
    exp_47_ram[2067] = 4;
    exp_47_ram[2068] = 164;
    exp_47_ram[2069] = 180;
    exp_47_ram[2070] = 196;
    exp_47_ram[2071] = 212;
    exp_47_ram[2072] = 228;
    exp_47_ram[2073] = 244;
    exp_47_ram[2074] = 4;
    exp_47_ram[2075] = 7;
    exp_47_ram[2076] = 64;
    exp_47_ram[2077] = 164;
    exp_47_ram[2078] = 180;
    exp_47_ram[2079] = 68;
    exp_47_ram[2080] = 244;
    exp_47_ram[2081] = 32;
    exp_47_ram[2082] = 244;
    exp_47_ram[2083] = 240;
    exp_47_ram[2084] = 244;
    exp_47_ram[2085] = 16;
    exp_47_ram[2086] = 244;
    exp_47_ram[2087] = 4;
    exp_47_ram[2088] = 4;
    exp_47_ram[2089] = 4;
    exp_47_ram[2090] = 4;
    exp_47_ram[2091] = 68;
    exp_47_ram[2092] = 132;
    exp_47_ram[2093] = 196;
    exp_47_ram[2094] = 4;
    exp_47_ram[2095] = 68;
    exp_47_ram[2096] = 132;
    exp_47_ram[2097] = 196;
    exp_47_ram[2098] = 4;
    exp_47_ram[2099] = 100;
    exp_47_ram[2100] = 20;
    exp_47_ram[2101] = 4;
    exp_47_ram[2102] = 164;
    exp_47_ram[2103] = 180;
    exp_47_ram[2104] = 196;
    exp_47_ram[2105] = 212;
    exp_47_ram[2106] = 228;
    exp_47_ram[2107] = 244;
    exp_47_ram[2108] = 4;
    exp_47_ram[2109] = 7;
    exp_47_ram[2110] = 192;
    exp_47_ram[2111] = 164;
    exp_47_ram[2112] = 180;
    exp_47_ram[2113] = 4;
    exp_47_ram[2114] = 4;
    exp_47_ram[2115] = 68;
    exp_47_ram[2116] = 7;
    exp_47_ram[2117] = 144;
    exp_47_ram[2118] = 196;
    exp_47_ram[2119] = 132;
    exp_47_ram[2120] = 247;
    exp_47_ram[2121] = 244;
    exp_47_ram[2122] = 4;
    exp_47_ram[2123] = 68;
    exp_47_ram[2124] = 132;
    exp_47_ram[2125] = 196;
    exp_47_ram[2126] = 4;
    exp_47_ram[2127] = 68;
    exp_47_ram[2128] = 132;
    exp_47_ram[2129] = 196;
    exp_47_ram[2130] = 4;
    exp_47_ram[2131] = 100;
    exp_47_ram[2132] = 20;
    exp_47_ram[2133] = 4;
    exp_47_ram[2134] = 164;
    exp_47_ram[2135] = 180;
    exp_47_ram[2136] = 196;
    exp_47_ram[2137] = 212;
    exp_47_ram[2138] = 228;
    exp_47_ram[2139] = 244;
    exp_47_ram[2140] = 4;
    exp_47_ram[2141] = 7;
    exp_47_ram[2142] = 192;
    exp_47_ram[2143] = 164;
    exp_47_ram[2144] = 180;
    exp_47_ram[2145] = 4;
    exp_47_ram[2146] = 68;
    exp_47_ram[2147] = 132;
    exp_47_ram[2148] = 196;
    exp_47_ram[2149] = 4;
    exp_47_ram[2150] = 68;
    exp_47_ram[2151] = 132;
    exp_47_ram[2152] = 196;
    exp_47_ram[2153] = 4;
    exp_47_ram[2154] = 100;
    exp_47_ram[2155] = 20;
    exp_47_ram[2156] = 4;
    exp_47_ram[2157] = 164;
    exp_47_ram[2158] = 180;
    exp_47_ram[2159] = 196;
    exp_47_ram[2160] = 212;
    exp_47_ram[2161] = 228;
    exp_47_ram[2162] = 244;
    exp_47_ram[2163] = 4;
    exp_47_ram[2164] = 7;
    exp_47_ram[2165] = 0;
    exp_47_ram[2166] = 164;
    exp_47_ram[2167] = 180;
    exp_47_ram[2168] = 68;
    exp_47_ram[2169] = 196;
    exp_47_ram[2170] = 231;
    exp_47_ram[2171] = 68;
    exp_47_ram[2172] = 196;
    exp_47_ram[2173] = 247;
    exp_47_ram[2174] = 4;
    exp_47_ram[2175] = 132;
    exp_47_ram[2176] = 231;
    exp_47_ram[2177] = 196;
    exp_47_ram[2178] = 196;
    exp_47_ram[2179] = 231;
    exp_47_ram[2180] = 196;
    exp_47_ram[2181] = 196;
    exp_47_ram[2182] = 247;
    exp_47_ram[2183] = 132;
    exp_47_ram[2184] = 132;
    exp_47_ram[2185] = 231;
    exp_47_ram[2186] = 16;
    exp_47_ram[2187] = 128;
    exp_47_ram[2188] = 0;
    exp_47_ram[2189] = 7;
    exp_47_ram[2190] = 193;
    exp_47_ram[2191] = 129;
    exp_47_ram[2192] = 65;
    exp_47_ram[2193] = 1;
    exp_47_ram[2194] = 0;
    exp_47_ram[2195] = 1;
    exp_47_ram[2196] = 17;
    exp_47_ram[2197] = 129;
    exp_47_ram[2198] = 1;
    exp_47_ram[2199] = 164;
    exp_47_ram[2200] = 180;
    exp_47_ram[2201] = 196;
    exp_47_ram[2202] = 132;
    exp_47_ram[2203] = 196;
    exp_47_ram[2204] = 7;
    exp_47_ram[2205] = 144;
    exp_47_ram[2206] = 196;
    exp_47_ram[2207] = 4;
    exp_47_ram[2208] = 68;
    exp_47_ram[2209] = 132;
    exp_47_ram[2210] = 196;
    exp_47_ram[2211] = 4;
    exp_47_ram[2212] = 68;
    exp_47_ram[2213] = 132;
    exp_47_ram[2214] = 196;
    exp_47_ram[2215] = 100;
    exp_47_ram[2216] = 20;
    exp_47_ram[2217] = 4;
    exp_47_ram[2218] = 164;
    exp_47_ram[2219] = 180;
    exp_47_ram[2220] = 196;
    exp_47_ram[2221] = 212;
    exp_47_ram[2222] = 228;
    exp_47_ram[2223] = 244;
    exp_47_ram[2224] = 4;
    exp_47_ram[2225] = 7;
    exp_47_ram[2226] = 95;
    exp_47_ram[2227] = 5;
    exp_47_ram[2228] = 7;
    exp_47_ram[2229] = 193;
    exp_47_ram[2230] = 129;
    exp_47_ram[2231] = 1;
    exp_47_ram[2232] = 0;
    exp_47_ram[2233] = 1;
    exp_47_ram[2234] = 129;
    exp_47_ram[2235] = 1;
    exp_47_ram[2236] = 0;
    exp_47_ram[2237] = 212;
    exp_47_ram[2238] = 0;
    exp_47_ram[2239] = 70;
    exp_47_ram[2240] = 212;
    exp_47_ram[2241] = 196;
    exp_47_ram[2242] = 6;
    exp_47_ram[2243] = 70;
    exp_47_ram[2244] = 132;
    exp_47_ram[2245] = 72;
    exp_47_ram[2246] = 8;
    exp_47_ram[2247] = 8;
    exp_47_ram[2248] = 0;
    exp_47_ram[2249] = 230;
    exp_47_ram[2250] = 246;
    exp_47_ram[2251] = 5;
    exp_47_ram[2252] = 5;
    exp_47_ram[2253] = 7;
    exp_47_ram[2254] = 7;
    exp_47_ram[2255] = 193;
    exp_47_ram[2256] = 1;
    exp_47_ram[2257] = 0;
    exp_47_ram[2258] = 1;
    exp_47_ram[2259] = 17;
    exp_47_ram[2260] = 129;
    exp_47_ram[2261] = 1;
    exp_47_ram[2262] = 164;
    exp_47_ram[2263] = 180;
    exp_47_ram[2264] = 196;
    exp_47_ram[2265] = 212;
    exp_47_ram[2266] = 132;
    exp_47_ram[2267] = 196;
    exp_47_ram[2268] = 4;
    exp_47_ram[2269] = 68;
    exp_47_ram[2270] = 167;
    exp_47_ram[2271] = 6;
    exp_47_ram[2272] = 7;
    exp_47_ram[2273] = 183;
    exp_47_ram[2274] = 6;
    exp_47_ram[2275] = 7;
    exp_47_ram[2276] = 6;
    exp_47_ram[2277] = 6;
    exp_47_ram[2278] = 7;
    exp_47_ram[2279] = 7;
    exp_47_ram[2280] = 79;
    exp_47_ram[2281] = 5;
    exp_47_ram[2282] = 5;
    exp_47_ram[2283] = 7;
    exp_47_ram[2284] = 7;
    exp_47_ram[2285] = 193;
    exp_47_ram[2286] = 129;
    exp_47_ram[2287] = 1;
    exp_47_ram[2288] = 0;
    exp_47_ram[2289] = 1;
    exp_47_ram[2290] = 129;
    exp_47_ram[2291] = 1;
    exp_47_ram[2292] = 164;
    exp_47_ram[2293] = 196;
    exp_47_ram[2294] = 55;
    exp_47_ram[2295] = 7;
    exp_47_ram[2296] = 196;
    exp_47_ram[2297] = 64;
    exp_47_ram[2298] = 247;
    exp_47_ram[2299] = 7;
    exp_47_ram[2300] = 196;
    exp_47_ram[2301] = 0;
    exp_47_ram[2302] = 247;
    exp_47_ram[2303] = 7;
    exp_47_ram[2304] = 16;
    exp_47_ram[2305] = 128;
    exp_47_ram[2306] = 0;
    exp_47_ram[2307] = 7;
    exp_47_ram[2308] = 193;
    exp_47_ram[2309] = 1;
    exp_47_ram[2310] = 0;
    exp_47_ram[2311] = 1;
    exp_47_ram[2312] = 17;
    exp_47_ram[2313] = 129;
    exp_47_ram[2314] = 1;
    exp_47_ram[2315] = 164;
    exp_47_ram[2316] = 196;
    exp_47_ram[2317] = 31;
    exp_47_ram[2318] = 5;
    exp_47_ram[2319] = 7;
    exp_47_ram[2320] = 224;
    exp_47_ram[2321] = 128;
    exp_47_ram[2322] = 208;
    exp_47_ram[2323] = 7;
    exp_47_ram[2324] = 193;
    exp_47_ram[2325] = 129;
    exp_47_ram[2326] = 1;
    exp_47_ram[2327] = 0;
    exp_47_ram[2328] = 1;
    exp_47_ram[2329] = 17;
    exp_47_ram[2330] = 129;
    exp_47_ram[2331] = 1;
    exp_47_ram[2332] = 164;
    exp_47_ram[2333] = 180;
    exp_47_ram[2334] = 132;
    exp_47_ram[2335] = 48;
    exp_47_ram[2336] = 247;
    exp_47_ram[2337] = 132;
    exp_47_ram[2338] = 128;
    exp_47_ram[2339] = 247;
    exp_47_ram[2340] = 132;
    exp_47_ram[2341] = 80;
    exp_47_ram[2342] = 247;
    exp_47_ram[2343] = 132;
    exp_47_ram[2344] = 160;
    exp_47_ram[2345] = 247;
    exp_47_ram[2346] = 224;
    exp_47_ram[2347] = 64;
    exp_47_ram[2348] = 132;
    exp_47_ram[2349] = 16;
    exp_47_ram[2350] = 247;
    exp_47_ram[2351] = 196;
    exp_47_ram[2352] = 95;
    exp_47_ram[2353] = 5;
    exp_47_ram[2354] = 7;
    exp_47_ram[2355] = 208;
    exp_47_ram[2356] = 0;
    exp_47_ram[2357] = 192;
    exp_47_ram[2358] = 128;
    exp_47_ram[2359] = 240;
    exp_47_ram[2360] = 7;
    exp_47_ram[2361] = 193;
    exp_47_ram[2362] = 129;
    exp_47_ram[2363] = 1;
    exp_47_ram[2364] = 0;
    exp_47_ram[2365] = 1;
    exp_47_ram[2366] = 17;
    exp_47_ram[2367] = 129;
    exp_47_ram[2368] = 145;
    exp_47_ram[2369] = 33;
    exp_47_ram[2370] = 49;
    exp_47_ram[2371] = 65;
    exp_47_ram[2372] = 81;
    exp_47_ram[2373] = 97;
    exp_47_ram[2374] = 113;
    exp_47_ram[2375] = 129;
    exp_47_ram[2376] = 145;
    exp_47_ram[2377] = 161;
    exp_47_ram[2378] = 177;
    exp_47_ram[2379] = 1;
    exp_47_ram[2380] = 5;
    exp_47_ram[2381] = 0;
    exp_47_ram[2382] = 0;
    exp_47_ram[2383] = 244;
    exp_47_ram[2384] = 4;
    exp_47_ram[2385] = 32;
    exp_47_ram[2386] = 244;
    exp_47_ram[2387] = 68;
    exp_47_ram[2388] = 244;
    exp_47_ram[2389] = 196;
    exp_47_ram[2390] = 199;
    exp_47_ram[2391] = 68;
    exp_47_ram[2392] = 247;
    exp_47_ram[2393] = 68;
    exp_47_ram[2394] = 95;
    exp_47_ram[2395] = 5;
    exp_47_ram[2396] = 1;
    exp_47_ram[2397] = 7;
    exp_47_ram[2398] = 247;
    exp_47_ram[2399] = 244;
    exp_47_ram[2400] = 4;
    exp_47_ram[2401] = 132;
    exp_47_ram[2402] = 196;
    exp_47_ram[2403] = 132;
    exp_47_ram[2404] = 196;
    exp_47_ram[2405] = 8;
    exp_47_ram[2406] = 182;
    exp_47_ram[2407] = 7;
    exp_47_ram[2408] = 197;
    exp_47_ram[2409] = 8;
    exp_47_ram[2410] = 166;
    exp_47_ram[2411] = 245;
    exp_47_ram[2412] = 6;
    exp_47_ram[2413] = 228;
    exp_47_ram[2414] = 244;
    exp_47_ram[2415] = 68;
    exp_47_ram[2416] = 23;
    exp_47_ram[2417] = 244;
    exp_47_ram[2418] = 223;
    exp_47_ram[2419] = 0;
    exp_47_ram[2420] = 4;
    exp_47_ram[2421] = 4;
    exp_47_ram[2422] = 7;
    exp_47_ram[2423] = 4;
    exp_47_ram[2424] = 231;
    exp_47_ram[2425] = 4;
    exp_47_ram[2426] = 68;
    exp_47_ram[2427] = 95;
    exp_47_ram[2428] = 5;
    exp_47_ram[2429] = 1;
    exp_47_ram[2430] = 7;
    exp_47_ram[2431] = 247;
    exp_47_ram[2432] = 7;
    exp_47_ram[2433] = 0;
    exp_47_ram[2434] = 132;
    exp_47_ram[2435] = 196;
    exp_47_ram[2436] = 166;
    exp_47_ram[2437] = 7;
    exp_47_ram[2438] = 197;
    exp_47_ram[2439] = 182;
    exp_47_ram[2440] = 245;
    exp_47_ram[2441] = 6;
    exp_47_ram[2442] = 228;
    exp_47_ram[2443] = 244;
    exp_47_ram[2444] = 4;
    exp_47_ram[2445] = 23;
    exp_47_ram[2446] = 244;
    exp_47_ram[2447] = 159;
    exp_47_ram[2448] = 0;
    exp_47_ram[2449] = 196;
    exp_47_ram[2450] = 247;
    exp_47_ram[2451] = 1;
    exp_47_ram[2452] = 7;
    exp_47_ram[2453] = 247;
    exp_47_ram[2454] = 7;
    exp_47_ram[2455] = 247;
    exp_47_ram[2456] = 7;
    exp_47_ram[2457] = 132;
    exp_47_ram[2458] = 196;
    exp_47_ram[2459] = 134;
    exp_47_ram[2460] = 7;
    exp_47_ram[2461] = 197;
    exp_47_ram[2462] = 150;
    exp_47_ram[2463] = 245;
    exp_47_ram[2464] = 6;
    exp_47_ram[2465] = 228;
    exp_47_ram[2466] = 244;
    exp_47_ram[2467] = 132;
    exp_47_ram[2468] = 0;
    exp_47_ram[2469] = 7;
    exp_47_ram[2470] = 247;
    exp_47_ram[2471] = 7;
    exp_47_ram[2472] = 247;
    exp_47_ram[2473] = 7;
    exp_47_ram[2474] = 132;
    exp_47_ram[2475] = 196;
    exp_47_ram[2476] = 102;
    exp_47_ram[2477] = 7;
    exp_47_ram[2478] = 197;
    exp_47_ram[2479] = 118;
    exp_47_ram[2480] = 245;
    exp_47_ram[2481] = 6;
    exp_47_ram[2482] = 228;
    exp_47_ram[2483] = 244;
    exp_47_ram[2484] = 68;
    exp_47_ram[2485] = 7;
    exp_47_ram[2486] = 71;
    exp_47_ram[2487] = 231;
    exp_47_ram[2488] = 39;
    exp_47_ram[2489] = 7;
    exp_47_ram[2490] = 247;
    exp_47_ram[2491] = 7;
    exp_47_ram[2492] = 132;
    exp_47_ram[2493] = 196;
    exp_47_ram[2494] = 70;
    exp_47_ram[2495] = 7;
    exp_47_ram[2496] = 197;
    exp_47_ram[2497] = 86;
    exp_47_ram[2498] = 245;
    exp_47_ram[2499] = 6;
    exp_47_ram[2500] = 228;
    exp_47_ram[2501] = 244;
    exp_47_ram[2502] = 4;
    exp_47_ram[2503] = 7;
    exp_47_ram[2504] = 247;
    exp_47_ram[2505] = 7;
    exp_47_ram[2506] = 132;
    exp_47_ram[2507] = 196;
    exp_47_ram[2508] = 38;
    exp_47_ram[2509] = 7;
    exp_47_ram[2510] = 197;
    exp_47_ram[2511] = 54;
    exp_47_ram[2512] = 245;
    exp_47_ram[2513] = 6;
    exp_47_ram[2514] = 228;
    exp_47_ram[2515] = 244;
    exp_47_ram[2516] = 132;
    exp_47_ram[2517] = 196;
    exp_47_ram[2518] = 7;
    exp_47_ram[2519] = 7;
    exp_47_ram[2520] = 193;
    exp_47_ram[2521] = 129;
    exp_47_ram[2522] = 65;
    exp_47_ram[2523] = 1;
    exp_47_ram[2524] = 193;
    exp_47_ram[2525] = 129;
    exp_47_ram[2526] = 65;
    exp_47_ram[2527] = 1;
    exp_47_ram[2528] = 193;
    exp_47_ram[2529] = 129;
    exp_47_ram[2530] = 65;
    exp_47_ram[2531] = 1;
    exp_47_ram[2532] = 193;
    exp_47_ram[2533] = 1;
    exp_47_ram[2534] = 0;
    exp_47_ram[2535] = 1;
    exp_47_ram[2536] = 17;
    exp_47_ram[2537] = 129;
    exp_47_ram[2538] = 145;
    exp_47_ram[2539] = 33;
    exp_47_ram[2540] = 49;
    exp_47_ram[2541] = 1;
    exp_47_ram[2542] = 164;
    exp_47_ram[2543] = 196;
    exp_47_ram[2544] = 7;
    exp_47_ram[2545] = 71;
    exp_47_ram[2546] = 135;
    exp_47_ram[2547] = 199;
    exp_47_ram[2548] = 7;
    exp_47_ram[2549] = 71;
    exp_47_ram[2550] = 135;
    exp_47_ram[2551] = 199;
    exp_47_ram[2552] = 7;
    exp_47_ram[2553] = 100;
    exp_47_ram[2554] = 20;
    exp_47_ram[2555] = 4;
    exp_47_ram[2556] = 164;
    exp_47_ram[2557] = 180;
    exp_47_ram[2558] = 196;
    exp_47_ram[2559] = 212;
    exp_47_ram[2560] = 228;
    exp_47_ram[2561] = 244;
    exp_47_ram[2562] = 196;
    exp_47_ram[2563] = 4;
    exp_47_ram[2564] = 68;
    exp_47_ram[2565] = 132;
    exp_47_ram[2566] = 196;
    exp_47_ram[2567] = 4;
    exp_47_ram[2568] = 68;
    exp_47_ram[2569] = 132;
    exp_47_ram[2570] = 196;
    exp_47_ram[2571] = 100;
    exp_47_ram[2572] = 20;
    exp_47_ram[2573] = 4;
    exp_47_ram[2574] = 164;
    exp_47_ram[2575] = 180;
    exp_47_ram[2576] = 196;
    exp_47_ram[2577] = 212;
    exp_47_ram[2578] = 228;
    exp_47_ram[2579] = 244;
    exp_47_ram[2580] = 4;
    exp_47_ram[2581] = 7;
    exp_47_ram[2582] = 223;
    exp_47_ram[2583] = 164;
    exp_47_ram[2584] = 180;
    exp_47_ram[2585] = 196;
    exp_47_ram[2586] = 240;
    exp_47_ram[2587] = 4;
    exp_47_ram[2588] = 68;
    exp_47_ram[2589] = 255;
    exp_47_ram[2590] = 5;
    exp_47_ram[2591] = 240;
    exp_47_ram[2592] = 166;
    exp_47_ram[2593] = 7;
    exp_47_ram[2594] = 200;
    exp_47_ram[2595] = 182;
    exp_47_ram[2596] = 248;
    exp_47_ram[2597] = 6;
    exp_47_ram[2598] = 228;
    exp_47_ram[2599] = 244;
    exp_47_ram[2600] = 192;
    exp_47_ram[2601] = 196;
    exp_47_ram[2602] = 7;
    exp_47_ram[2603] = 196;
    exp_47_ram[2604] = 4;
    exp_47_ram[2605] = 68;
    exp_47_ram[2606] = 132;
    exp_47_ram[2607] = 196;
    exp_47_ram[2608] = 4;
    exp_47_ram[2609] = 68;
    exp_47_ram[2610] = 132;
    exp_47_ram[2611] = 196;
    exp_47_ram[2612] = 100;
    exp_47_ram[2613] = 20;
    exp_47_ram[2614] = 4;
    exp_47_ram[2615] = 164;
    exp_47_ram[2616] = 180;
    exp_47_ram[2617] = 196;
    exp_47_ram[2618] = 212;
    exp_47_ram[2619] = 228;
    exp_47_ram[2620] = 244;
    exp_47_ram[2621] = 4;
    exp_47_ram[2622] = 7;
    exp_47_ram[2623] = 15;
    exp_47_ram[2624] = 5;
    exp_47_ram[2625] = 7;
    exp_47_ram[2626] = 0;
    exp_47_ram[2627] = 6;
    exp_47_ram[2628] = 0;
    exp_47_ram[2629] = 192;
    exp_47_ram[2630] = 0;
    exp_47_ram[2631] = 0;
    exp_47_ram[2632] = 4;
    exp_47_ram[2633] = 68;
    exp_47_ram[2634] = 197;
    exp_47_ram[2635] = 7;
    exp_47_ram[2636] = 5;
    exp_47_ram[2637] = 213;
    exp_47_ram[2638] = 7;
    exp_47_ram[2639] = 6;
    exp_47_ram[2640] = 228;
    exp_47_ram[2641] = 244;
    exp_47_ram[2642] = 64;
    exp_47_ram[2643] = 4;
    exp_47_ram[2644] = 68;
    exp_47_ram[2645] = 228;
    exp_47_ram[2646] = 244;
    exp_47_ram[2647] = 0;
    exp_47_ram[2648] = 7;
    exp_47_ram[2649] = 7;
    exp_47_ram[2650] = 247;
    exp_47_ram[2651] = 7;
    exp_47_ram[2652] = 132;
    exp_47_ram[2653] = 196;
    exp_47_ram[2654] = 38;
    exp_47_ram[2655] = 7;
    exp_47_ram[2656] = 182;
    exp_47_ram[2657] = 54;
    exp_47_ram[2658] = 183;
    exp_47_ram[2659] = 6;
    exp_47_ram[2660] = 228;
    exp_47_ram[2661] = 244;
    exp_47_ram[2662] = 196;
    exp_47_ram[2663] = 4;
    exp_47_ram[2664] = 132;
    exp_47_ram[2665] = 196;
    exp_47_ram[2666] = 7;
    exp_47_ram[2667] = 0;
    exp_47_ram[2668] = 4;
    exp_47_ram[2669] = 68;
    exp_47_ram[2670] = 132;
    exp_47_ram[2671] = 196;
    exp_47_ram[2672] = 4;
    exp_47_ram[2673] = 68;
    exp_47_ram[2674] = 132;
    exp_47_ram[2675] = 196;
    exp_47_ram[2676] = 4;
    exp_47_ram[2677] = 100;
    exp_47_ram[2678] = 20;
    exp_47_ram[2679] = 4;
    exp_47_ram[2680] = 164;
    exp_47_ram[2681] = 180;
    exp_47_ram[2682] = 196;
    exp_47_ram[2683] = 212;
    exp_47_ram[2684] = 228;
    exp_47_ram[2685] = 244;
    exp_47_ram[2686] = 196;
    exp_47_ram[2687] = 240;
    exp_47_ram[2688] = 196;
    exp_47_ram[2689] = 16;
    exp_47_ram[2690] = 231;
    exp_47_ram[2691] = 128;
    exp_47_ram[2692] = 196;
    exp_47_ram[2693] = 7;
    exp_47_ram[2694] = 196;
    exp_47_ram[2695] = 4;
    exp_47_ram[2696] = 68;
    exp_47_ram[2697] = 132;
    exp_47_ram[2698] = 196;
    exp_47_ram[2699] = 4;
    exp_47_ram[2700] = 68;
    exp_47_ram[2701] = 132;
    exp_47_ram[2702] = 196;
    exp_47_ram[2703] = 100;
    exp_47_ram[2704] = 20;
    exp_47_ram[2705] = 4;
    exp_47_ram[2706] = 164;
    exp_47_ram[2707] = 180;
    exp_47_ram[2708] = 196;
    exp_47_ram[2709] = 212;
    exp_47_ram[2710] = 228;
    exp_47_ram[2711] = 244;
    exp_47_ram[2712] = 4;
    exp_47_ram[2713] = 7;
    exp_47_ram[2714] = 79;
    exp_47_ram[2715] = 5;
    exp_47_ram[2716] = 196;
    exp_47_ram[2717] = 231;
    exp_47_ram[2718] = 192;
    exp_47_ram[2719] = 196;
    exp_47_ram[2720] = 7;
    exp_47_ram[2721] = 132;
    exp_47_ram[2722] = 196;
    exp_47_ram[2723] = 7;
    exp_47_ram[2724] = 7;
    exp_47_ram[2725] = 193;
    exp_47_ram[2726] = 129;
    exp_47_ram[2727] = 65;
    exp_47_ram[2728] = 1;
    exp_47_ram[2729] = 193;
    exp_47_ram[2730] = 1;
    exp_47_ram[2731] = 0;
    exp_47_ram[2732] = 1;
    exp_47_ram[2733] = 17;
    exp_47_ram[2734] = 129;
    exp_47_ram[2735] = 33;
    exp_47_ram[2736] = 49;
    exp_47_ram[2737] = 65;
    exp_47_ram[2738] = 81;
    exp_47_ram[2739] = 97;
    exp_47_ram[2740] = 113;
    exp_47_ram[2741] = 1;
    exp_47_ram[2742] = 164;
    exp_47_ram[2743] = 159;
    exp_47_ram[2744] = 5;
    exp_47_ram[2745] = 5;
    exp_47_ram[2746] = 0;
    exp_47_ram[2747] = 6;
    exp_47_ram[2748] = 6;
    exp_47_ram[2749] = 0;
    exp_47_ram[2750] = 10;
    exp_47_ram[2751] = 10;
    exp_47_ram[2752] = 7;
    exp_47_ram[2753] = 7;
    exp_47_ram[2754] = 79;
    exp_47_ram[2755] = 5;
    exp_47_ram[2756] = 5;
    exp_47_ram[2757] = 228;
    exp_47_ram[2758] = 0;
    exp_47_ram[2759] = 135;
    exp_47_ram[2760] = 199;
    exp_47_ram[2761] = 196;
    exp_47_ram[2762] = 231;
    exp_47_ram[2763] = 244;
    exp_47_ram[2764] = 196;
    exp_47_ram[2765] = 7;
    exp_47_ram[2766] = 196;
    exp_47_ram[2767] = 7;
    exp_47_ram[2768] = 0;
    exp_47_ram[2769] = 196;
    exp_47_ram[2770] = 39;
    exp_47_ram[2771] = 55;
    exp_47_ram[2772] = 196;
    exp_47_ram[2773] = 7;
    exp_47_ram[2774] = 0;
    exp_47_ram[2775] = 11;
    exp_47_ram[2776] = 11;
    exp_47_ram[2777] = 7;
    exp_47_ram[2778] = 7;
    exp_47_ram[2779] = 193;
    exp_47_ram[2780] = 129;
    exp_47_ram[2781] = 65;
    exp_47_ram[2782] = 1;
    exp_47_ram[2783] = 193;
    exp_47_ram[2784] = 129;
    exp_47_ram[2785] = 65;
    exp_47_ram[2786] = 1;
    exp_47_ram[2787] = 1;
    exp_47_ram[2788] = 0;
    exp_47_ram[2789] = 1;
    exp_47_ram[2790] = 17;
    exp_47_ram[2791] = 129;
    exp_47_ram[2792] = 33;
    exp_47_ram[2793] = 49;
    exp_47_ram[2794] = 1;
    exp_47_ram[2795] = 164;
    exp_47_ram[2796] = 180;
    exp_47_ram[2797] = 15;
    exp_47_ram[2798] = 5;
    exp_47_ram[2799] = 5;
    exp_47_ram[2800] = 0;
    exp_47_ram[2801] = 6;
    exp_47_ram[2802] = 6;
    exp_47_ram[2803] = 0;
    exp_47_ram[2804] = 9;
    exp_47_ram[2805] = 9;
    exp_47_ram[2806] = 7;
    exp_47_ram[2807] = 7;
    exp_47_ram[2808] = 207;
    exp_47_ram[2809] = 5;
    exp_47_ram[2810] = 5;
    exp_47_ram[2811] = 228;
    exp_47_ram[2812] = 244;
    exp_47_ram[2813] = 132;
    exp_47_ram[2814] = 196;
    exp_47_ram[2815] = 132;
    exp_47_ram[2816] = 196;
    exp_47_ram[2817] = 167;
    exp_47_ram[2818] = 6;
    exp_47_ram[2819] = 7;
    exp_47_ram[2820] = 183;
    exp_47_ram[2821] = 6;
    exp_47_ram[2822] = 7;
    exp_47_ram[2823] = 6;
    exp_47_ram[2824] = 6;
    exp_47_ram[2825] = 0;
    exp_47_ram[2826] = 230;
    exp_47_ram[2827] = 246;
    exp_47_ram[2828] = 0;
    exp_47_ram[2829] = 193;
    exp_47_ram[2830] = 129;
    exp_47_ram[2831] = 65;
    exp_47_ram[2832] = 1;
    exp_47_ram[2833] = 1;
    exp_47_ram[2834] = 0;
    exp_47_ram[2835] = 1;
    exp_47_ram[2836] = 17;
    exp_47_ram[2837] = 129;
    exp_47_ram[2838] = 1;
    exp_47_ram[2839] = 164;
    exp_47_ram[2840] = 0;
    exp_47_ram[2841] = 135;
    exp_47_ram[2842] = 7;
    exp_47_ram[2843] = 71;
    exp_47_ram[2844] = 135;
    exp_47_ram[2845] = 199;
    exp_47_ram[2846] = 7;
    exp_47_ram[2847] = 164;
    exp_47_ram[2848] = 180;
    exp_47_ram[2849] = 196;
    exp_47_ram[2850] = 212;
    exp_47_ram[2851] = 228;
    exp_47_ram[2852] = 71;
    exp_47_ram[2853] = 244;
    exp_47_ram[2854] = 0;
    exp_47_ram[2855] = 7;
    exp_47_ram[2856] = 7;
    exp_47_ram[2857] = 71;
    exp_47_ram[2858] = 135;
    exp_47_ram[2859] = 199;
    exp_47_ram[2860] = 7;
    exp_47_ram[2861] = 71;
    exp_47_ram[2862] = 135;
    exp_47_ram[2863] = 199;
    exp_47_ram[2864] = 7;
    exp_47_ram[2865] = 196;
    exp_47_ram[2866] = 100;
    exp_47_ram[2867] = 20;
    exp_47_ram[2868] = 4;
    exp_47_ram[2869] = 164;
    exp_47_ram[2870] = 180;
    exp_47_ram[2871] = 196;
    exp_47_ram[2872] = 212;
    exp_47_ram[2873] = 228;
    exp_47_ram[2874] = 71;
    exp_47_ram[2875] = 244;
    exp_47_ram[2876] = 4;
    exp_47_ram[2877] = 192;
    exp_47_ram[2878] = 196;
    exp_47_ram[2879] = 135;
    exp_47_ram[2880] = 7;
    exp_47_ram[2881] = 23;
    exp_47_ram[2882] = 231;
    exp_47_ram[2883] = 196;
    exp_47_ram[2884] = 247;
    exp_47_ram[2885] = 4;
    exp_47_ram[2886] = 247;
    exp_47_ram[2887] = 71;
    exp_47_ram[2888] = 0;
    exp_47_ram[2889] = 7;
    exp_47_ram[2890] = 196;
    exp_47_ram[2891] = 246;
    exp_47_ram[2892] = 231;
    exp_47_ram[2893] = 196;
    exp_47_ram[2894] = 23;
    exp_47_ram[2895] = 244;
    exp_47_ram[2896] = 196;
    exp_47_ram[2897] = 32;
    exp_47_ram[2898] = 231;
    exp_47_ram[2899] = 0;
    exp_47_ram[2900] = 7;
    exp_47_ram[2901] = 0;
    exp_47_ram[2902] = 231;
    exp_47_ram[2903] = 4;
    exp_47_ram[2904] = 0;
    exp_47_ram[2905] = 196;
    exp_47_ram[2906] = 7;
    exp_47_ram[2907] = 7;
    exp_47_ram[2908] = 23;
    exp_47_ram[2909] = 231;
    exp_47_ram[2910] = 196;
    exp_47_ram[2911] = 247;
    exp_47_ram[2912] = 196;
    exp_47_ram[2913] = 71;
    exp_47_ram[2914] = 4;
    exp_47_ram[2915] = 230;
    exp_47_ram[2916] = 199;
    exp_47_ram[2917] = 0;
    exp_47_ram[2918] = 6;
    exp_47_ram[2919] = 246;
    exp_47_ram[2920] = 231;
    exp_47_ram[2921] = 196;
    exp_47_ram[2922] = 23;
    exp_47_ram[2923] = 244;
    exp_47_ram[2924] = 196;
    exp_47_ram[2925] = 32;
    exp_47_ram[2926] = 231;
    exp_47_ram[2927] = 0;
    exp_47_ram[2928] = 7;
    exp_47_ram[2929] = 0;
    exp_47_ram[2930] = 231;
    exp_47_ram[2931] = 196;
    exp_47_ram[2932] = 199;
    exp_47_ram[2933] = 160;
    exp_47_ram[2934] = 7;
    exp_47_ram[2935] = 128;
    exp_47_ram[2936] = 5;
    exp_47_ram[2937] = 5;
    exp_47_ram[2938] = 228;
    exp_47_ram[2939] = 244;
    exp_47_ram[2940] = 68;
    exp_47_ram[2941] = 247;
    exp_47_ram[2942] = 7;
    exp_47_ram[2943] = 247;
    exp_47_ram[2944] = 0;
    exp_47_ram[2945] = 7;
    exp_47_ram[2946] = 231;
    exp_47_ram[2947] = 132;
    exp_47_ram[2948] = 247;
    exp_47_ram[2949] = 7;
    exp_47_ram[2950] = 247;
    exp_47_ram[2951] = 0;
    exp_47_ram[2952] = 7;
    exp_47_ram[2953] = 231;
    exp_47_ram[2954] = 0;
    exp_47_ram[2955] = 7;
    exp_47_ram[2956] = 0;
    exp_47_ram[2957] = 231;
    exp_47_ram[2958] = 196;
    exp_47_ram[2959] = 135;
    exp_47_ram[2960] = 160;
    exp_47_ram[2961] = 7;
    exp_47_ram[2962] = 192;
    exp_47_ram[2963] = 5;
    exp_47_ram[2964] = 5;
    exp_47_ram[2965] = 228;
    exp_47_ram[2966] = 244;
    exp_47_ram[2967] = 68;
    exp_47_ram[2968] = 247;
    exp_47_ram[2969] = 7;
    exp_47_ram[2970] = 247;
    exp_47_ram[2971] = 0;
    exp_47_ram[2972] = 7;
    exp_47_ram[2973] = 231;
    exp_47_ram[2974] = 132;
    exp_47_ram[2975] = 247;
    exp_47_ram[2976] = 7;
    exp_47_ram[2977] = 247;
    exp_47_ram[2978] = 0;
    exp_47_ram[2979] = 7;
    exp_47_ram[2980] = 231;
    exp_47_ram[2981] = 0;
    exp_47_ram[2982] = 7;
    exp_47_ram[2983] = 160;
    exp_47_ram[2984] = 231;
    exp_47_ram[2985] = 196;
    exp_47_ram[2986] = 71;
    exp_47_ram[2987] = 160;
    exp_47_ram[2988] = 7;
    exp_47_ram[2989] = 0;
    exp_47_ram[2990] = 5;
    exp_47_ram[2991] = 5;
    exp_47_ram[2992] = 228;
    exp_47_ram[2993] = 244;
    exp_47_ram[2994] = 68;
    exp_47_ram[2995] = 247;
    exp_47_ram[2996] = 7;
    exp_47_ram[2997] = 247;
    exp_47_ram[2998] = 0;
    exp_47_ram[2999] = 7;
    exp_47_ram[3000] = 231;
    exp_47_ram[3001] = 132;
    exp_47_ram[3002] = 247;
    exp_47_ram[3003] = 7;
    exp_47_ram[3004] = 247;
    exp_47_ram[3005] = 0;
    exp_47_ram[3006] = 7;
    exp_47_ram[3007] = 231;
    exp_47_ram[3008] = 0;
    exp_47_ram[3009] = 7;
    exp_47_ram[3010] = 160;
    exp_47_ram[3011] = 231;
    exp_47_ram[3012] = 196;
    exp_47_ram[3013] = 7;
    exp_47_ram[3014] = 160;
    exp_47_ram[3015] = 7;
    exp_47_ram[3016] = 64;
    exp_47_ram[3017] = 5;
    exp_47_ram[3018] = 5;
    exp_47_ram[3019] = 228;
    exp_47_ram[3020] = 244;
    exp_47_ram[3021] = 68;
    exp_47_ram[3022] = 247;
    exp_47_ram[3023] = 7;
    exp_47_ram[3024] = 247;
    exp_47_ram[3025] = 0;
    exp_47_ram[3026] = 7;
    exp_47_ram[3027] = 231;
    exp_47_ram[3028] = 132;
    exp_47_ram[3029] = 247;
    exp_47_ram[3030] = 7;
    exp_47_ram[3031] = 247;
    exp_47_ram[3032] = 0;
    exp_47_ram[3033] = 7;
    exp_47_ram[3034] = 231;
    exp_47_ram[3035] = 0;
    exp_47_ram[3036] = 7;
    exp_47_ram[3037] = 0;
    exp_47_ram[3038] = 231;
    exp_47_ram[3039] = 196;
    exp_47_ram[3040] = 71;
    exp_47_ram[3041] = 199;
    exp_47_ram[3042] = 128;
    exp_47_ram[3043] = 7;
    exp_47_ram[3044] = 64;
    exp_47_ram[3045] = 5;
    exp_47_ram[3046] = 5;
    exp_47_ram[3047] = 228;
    exp_47_ram[3048] = 244;
    exp_47_ram[3049] = 68;
    exp_47_ram[3050] = 247;
    exp_47_ram[3051] = 7;
    exp_47_ram[3052] = 247;
    exp_47_ram[3053] = 0;
    exp_47_ram[3054] = 7;
    exp_47_ram[3055] = 231;
    exp_47_ram[3056] = 132;
    exp_47_ram[3057] = 64;
    exp_47_ram[3058] = 7;
    exp_47_ram[3059] = 128;
    exp_47_ram[3060] = 5;
    exp_47_ram[3061] = 5;
    exp_47_ram[3062] = 228;
    exp_47_ram[3063] = 244;
    exp_47_ram[3064] = 68;
    exp_47_ram[3065] = 247;
    exp_47_ram[3066] = 7;
    exp_47_ram[3067] = 247;
    exp_47_ram[3068] = 0;
    exp_47_ram[3069] = 7;
    exp_47_ram[3070] = 231;
    exp_47_ram[3071] = 132;
    exp_47_ram[3072] = 160;
    exp_47_ram[3073] = 7;
    exp_47_ram[3074] = 192;
    exp_47_ram[3075] = 5;
    exp_47_ram[3076] = 5;
    exp_47_ram[3077] = 228;
    exp_47_ram[3078] = 244;
    exp_47_ram[3079] = 68;
    exp_47_ram[3080] = 247;
    exp_47_ram[3081] = 7;
    exp_47_ram[3082] = 247;
    exp_47_ram[3083] = 0;
    exp_47_ram[3084] = 7;
    exp_47_ram[3085] = 231;
    exp_47_ram[3086] = 132;
    exp_47_ram[3087] = 247;
    exp_47_ram[3088] = 7;
    exp_47_ram[3089] = 247;
    exp_47_ram[3090] = 0;
    exp_47_ram[3091] = 7;
    exp_47_ram[3092] = 231;
    exp_47_ram[3093] = 0;
    exp_47_ram[3094] = 7;
    exp_47_ram[3095] = 160;
    exp_47_ram[3096] = 231;
    exp_47_ram[3097] = 0;
    exp_47_ram[3098] = 7;
    exp_47_ram[3099] = 7;
    exp_47_ram[3100] = 0;
    exp_47_ram[3101] = 7;
    exp_47_ram[3102] = 7;
    exp_47_ram[3103] = 193;
    exp_47_ram[3104] = 129;
    exp_47_ram[3105] = 1;
    exp_47_ram[3106] = 0;
    exp_47_ram[3107] = 1;
    exp_47_ram[3108] = 17;
    exp_47_ram[3109] = 129;
    exp_47_ram[3110] = 1;
    exp_47_ram[3111] = 164;
    exp_47_ram[3112] = 196;
    exp_47_ram[3113] = 64;
    exp_47_ram[3114] = 5;
    exp_47_ram[3115] = 7;
    exp_47_ram[3116] = 223;
    exp_47_ram[3117] = 5;
    exp_47_ram[3118] = 7;
    exp_47_ram[3119] = 193;
    exp_47_ram[3120] = 129;
    exp_47_ram[3121] = 1;
    exp_47_ram[3122] = 0;
    exp_47_ram[3123] = 1;
    exp_47_ram[3124] = 17;
    exp_47_ram[3125] = 129;
    exp_47_ram[3126] = 33;
    exp_47_ram[3127] = 49;
    exp_47_ram[3128] = 65;
    exp_47_ram[3129] = 81;
    exp_47_ram[3130] = 97;
    exp_47_ram[3131] = 113;
    exp_47_ram[3132] = 129;
    exp_47_ram[3133] = 145;
    exp_47_ram[3134] = 1;
    exp_47_ram[3135] = 164;
    exp_47_ram[3136] = 180;
    exp_47_ram[3137] = 196;
    exp_47_ram[3138] = 32;
    exp_47_ram[3139] = 244;
    exp_47_ram[3140] = 64;
    exp_47_ram[3141] = 244;
    exp_47_ram[3142] = 132;
    exp_47_ram[3143] = 7;
    exp_47_ram[3144] = 207;
    exp_47_ram[3145] = 164;
    exp_47_ram[3146] = 196;
    exp_47_ram[3147] = 1;
    exp_47_ram[3148] = 7;
    exp_47_ram[3149] = 247;
    exp_47_ram[3150] = 244;
    exp_47_ram[3151] = 132;
    exp_47_ram[3152] = 7;
    exp_47_ram[3153] = 0;
    exp_47_ram[3154] = 68;
    exp_47_ram[3155] = 12;
    exp_47_ram[3156] = 231;
    exp_47_ram[3157] = 68;
    exp_47_ram[3158] = 12;
    exp_47_ram[3159] = 231;
    exp_47_ram[3160] = 4;
    exp_47_ram[3161] = 12;
    exp_47_ram[3162] = 231;
    exp_47_ram[3163] = 132;
    exp_47_ram[3164] = 23;
    exp_47_ram[3165] = 244;
    exp_47_ram[3166] = 196;
    exp_47_ram[3167] = 7;
    exp_47_ram[3168] = 196;
    exp_47_ram[3169] = 247;
    exp_47_ram[3170] = 244;
    exp_47_ram[3171] = 132;
    exp_47_ram[3172] = 7;
    exp_47_ram[3173] = 0;
    exp_47_ram[3174] = 4;
    exp_47_ram[3175] = 68;
    exp_47_ram[3176] = 70;
    exp_47_ram[3177] = 7;
    exp_47_ram[3178] = 182;
    exp_47_ram[3179] = 86;
    exp_47_ram[3180] = 183;
    exp_47_ram[3181] = 6;
    exp_47_ram[3182] = 228;
    exp_47_ram[3183] = 244;
    exp_47_ram[3184] = 159;
    exp_47_ram[3185] = 0;
    exp_47_ram[3186] = 4;
    exp_47_ram[3187] = 4;
    exp_47_ram[3188] = 132;
    exp_47_ram[3189] = 7;
    exp_47_ram[3190] = 68;
    exp_47_ram[3191] = 7;
    exp_47_ram[3192] = 7;
    exp_47_ram[3193] = 207;
    exp_47_ram[3194] = 164;
    exp_47_ram[3195] = 196;
    exp_47_ram[3196] = 1;
    exp_47_ram[3197] = 7;
    exp_47_ram[3198] = 247;
    exp_47_ram[3199] = 244;
    exp_47_ram[3200] = 132;
    exp_47_ram[3201] = 7;
    exp_47_ram[3202] = 0;
    exp_47_ram[3203] = 68;
    exp_47_ram[3204] = 11;
    exp_47_ram[3205] = 231;
    exp_47_ram[3206] = 68;
    exp_47_ram[3207] = 11;
    exp_47_ram[3208] = 231;
    exp_47_ram[3209] = 4;
    exp_47_ram[3210] = 11;
    exp_47_ram[3211] = 231;
    exp_47_ram[3212] = 68;
    exp_47_ram[3213] = 23;
    exp_47_ram[3214] = 244;
    exp_47_ram[3215] = 196;
    exp_47_ram[3216] = 7;
    exp_47_ram[3217] = 196;
    exp_47_ram[3218] = 247;
    exp_47_ram[3219] = 244;
    exp_47_ram[3220] = 4;
    exp_47_ram[3221] = 7;
    exp_47_ram[3222] = 196;
    exp_47_ram[3223] = 247;
    exp_47_ram[3224] = 244;
    exp_47_ram[3225] = 132;
    exp_47_ram[3226] = 7;
    exp_47_ram[3227] = 0;
    exp_47_ram[3228] = 4;
    exp_47_ram[3229] = 68;
    exp_47_ram[3230] = 38;
    exp_47_ram[3231] = 7;
    exp_47_ram[3232] = 182;
    exp_47_ram[3233] = 54;
    exp_47_ram[3234] = 183;
    exp_47_ram[3235] = 6;
    exp_47_ram[3236] = 228;
    exp_47_ram[3237] = 244;
    exp_47_ram[3238] = 159;
    exp_47_ram[3239] = 0;
    exp_47_ram[3240] = 132;
    exp_47_ram[3241] = 71;
    exp_47_ram[3242] = 244;
    exp_47_ram[3243] = 4;
    exp_47_ram[3244] = 1;
    exp_47_ram[3245] = 7;
    exp_47_ram[3246] = 7;
    exp_47_ram[3247] = 144;
    exp_47_ram[3248] = 5;
    exp_47_ram[3249] = 5;
    exp_47_ram[3250] = 228;
    exp_47_ram[3251] = 244;
    exp_47_ram[3252] = 196;
    exp_47_ram[3253] = 23;
    exp_47_ram[3254] = 244;
    exp_47_ram[3255] = 196;
    exp_47_ram[3256] = 196;
    exp_47_ram[3257] = 247;
    exp_47_ram[3258] = 244;
    exp_47_ram[3259] = 196;
    exp_47_ram[3260] = 112;
    exp_47_ram[3261] = 247;
    exp_47_ram[3262] = 244;
    exp_47_ram[3263] = 4;
    exp_47_ram[3264] = 196;
    exp_47_ram[3265] = 247;
    exp_47_ram[3266] = 244;
    exp_47_ram[3267] = 4;
    exp_47_ram[3268] = 244;
    exp_47_ram[3269] = 247;
    exp_47_ram[3270] = 244;
    exp_47_ram[3271] = 4;
    exp_47_ram[3272] = 0;
    exp_47_ram[3273] = 7;
    exp_47_ram[3274] = 7;
    exp_47_ram[3275] = 144;
    exp_47_ram[3276] = 5;
    exp_47_ram[3277] = 5;
    exp_47_ram[3278] = 228;
    exp_47_ram[3279] = 244;
    exp_47_ram[3280] = 196;
    exp_47_ram[3281] = 244;
    exp_47_ram[3282] = 4;
    exp_47_ram[3283] = 244;
    exp_47_ram[3284] = 247;
    exp_47_ram[3285] = 244;
    exp_47_ram[3286] = 4;
    exp_47_ram[3287] = 192;
    exp_47_ram[3288] = 7;
    exp_47_ram[3289] = 16;
    exp_47_ram[3290] = 5;
    exp_47_ram[3291] = 5;
    exp_47_ram[3292] = 228;
    exp_47_ram[3293] = 244;
    exp_47_ram[3294] = 196;
    exp_47_ram[3295] = 244;
    exp_47_ram[3296] = 4;
    exp_47_ram[3297] = 244;
    exp_47_ram[3298] = 247;
    exp_47_ram[3299] = 244;
    exp_47_ram[3300] = 4;
    exp_47_ram[3301] = 244;
    exp_47_ram[3302] = 196;
    exp_47_ram[3303] = 68;
    exp_47_ram[3304] = 132;
    exp_47_ram[3305] = 196;
    exp_47_ram[3306] = 4;
    exp_47_ram[3307] = 68;
    exp_47_ram[3308] = 132;
    exp_47_ram[3309] = 196;
    exp_47_ram[3310] = 4;
    exp_47_ram[3311] = 68;
    exp_47_ram[3312] = 199;
    exp_47_ram[3313] = 103;
    exp_47_ram[3314] = 23;
    exp_47_ram[3315] = 7;
    exp_47_ram[3316] = 167;
    exp_47_ram[3317] = 183;
    exp_47_ram[3318] = 199;
    exp_47_ram[3319] = 215;
    exp_47_ram[3320] = 231;
    exp_47_ram[3321] = 196;
    exp_47_ram[3322] = 193;
    exp_47_ram[3323] = 129;
    exp_47_ram[3324] = 65;
    exp_47_ram[3325] = 1;
    exp_47_ram[3326] = 193;
    exp_47_ram[3327] = 129;
    exp_47_ram[3328] = 65;
    exp_47_ram[3329] = 1;
    exp_47_ram[3330] = 193;
    exp_47_ram[3331] = 129;
    exp_47_ram[3332] = 1;
    exp_47_ram[3333] = 0;
    exp_47_ram[3334] = 1;
    exp_47_ram[3335] = 17;
    exp_47_ram[3336] = 129;
    exp_47_ram[3337] = 145;
    exp_47_ram[3338] = 33;
    exp_47_ram[3339] = 49;
    exp_47_ram[3340] = 1;
    exp_47_ram[3341] = 164;
    exp_47_ram[3342] = 0;
    exp_47_ram[3343] = 0;
    exp_47_ram[3344] = 244;
    exp_47_ram[3345] = 4;
    exp_47_ram[3346] = 196;
    exp_47_ram[3347] = 7;
    exp_47_ram[3348] = 71;
    exp_47_ram[3349] = 228;
    exp_47_ram[3350] = 244;
    exp_47_ram[3351] = 4;
    exp_47_ram[3352] = 68;
    exp_47_ram[3353] = 159;
    exp_47_ram[3354] = 5;
    exp_47_ram[3355] = 7;
    exp_47_ram[3356] = 0;
    exp_47_ram[3357] = 7;
    exp_47_ram[3358] = 0;
    exp_47_ram[3359] = 228;
    exp_47_ram[3360] = 244;
    exp_47_ram[3361] = 0;
    exp_47_ram[3362] = 7;
    exp_47_ram[3363] = 7;
    exp_47_ram[3364] = 247;
    exp_47_ram[3365] = 7;
    exp_47_ram[3366] = 4;
    exp_47_ram[3367] = 68;
    exp_47_ram[3368] = 201;
    exp_47_ram[3369] = 7;
    exp_47_ram[3370] = 37;
    exp_47_ram[3371] = 217;
    exp_47_ram[3372] = 245;
    exp_47_ram[3373] = 6;
    exp_47_ram[3374] = 7;
    exp_47_ram[3375] = 7;
    exp_47_ram[3376] = 132;
    exp_47_ram[3377] = 196;
    exp_47_ram[3378] = 166;
    exp_47_ram[3379] = 7;
    exp_47_ram[3380] = 200;
    exp_47_ram[3381] = 182;
    exp_47_ram[3382] = 248;
    exp_47_ram[3383] = 6;
    exp_47_ram[3384] = 228;
    exp_47_ram[3385] = 244;
    exp_47_ram[3386] = 0;
    exp_47_ram[3387] = 199;
    exp_47_ram[3388] = 4;
    exp_47_ram[3389] = 132;
    exp_47_ram[3390] = 196;
    exp_47_ram[3391] = 7;
    exp_47_ram[3392] = 223;
    exp_47_ram[3393] = 4;
    exp_47_ram[3394] = 68;
    exp_47_ram[3395] = 132;
    exp_47_ram[3396] = 196;
    exp_47_ram[3397] = 4;
    exp_47_ram[3398] = 68;
    exp_47_ram[3399] = 132;
    exp_47_ram[3400] = 196;
    exp_47_ram[3401] = 4;
    exp_47_ram[3402] = 100;
    exp_47_ram[3403] = 20;
    exp_47_ram[3404] = 4;
    exp_47_ram[3405] = 164;
    exp_47_ram[3406] = 180;
    exp_47_ram[3407] = 196;
    exp_47_ram[3408] = 212;
    exp_47_ram[3409] = 228;
    exp_47_ram[3410] = 244;
    exp_47_ram[3411] = 4;
    exp_47_ram[3412] = 68;
    exp_47_ram[3413] = 159;
    exp_47_ram[3414] = 5;
    exp_47_ram[3415] = 0;
    exp_47_ram[3416] = 199;
    exp_47_ram[3417] = 231;
    exp_47_ram[3418] = 0;
    exp_47_ram[3419] = 199;
    exp_47_ram[3420] = 7;
    exp_47_ram[3421] = 193;
    exp_47_ram[3422] = 129;
    exp_47_ram[3423] = 65;
    exp_47_ram[3424] = 1;
    exp_47_ram[3425] = 193;
    exp_47_ram[3426] = 1;
    exp_47_ram[3427] = 0;
    exp_47_ram[3428] = 1;
    exp_47_ram[3429] = 17;
    exp_47_ram[3430] = 129;
    exp_47_ram[3431] = 1;
    exp_47_ram[3432] = 164;
    exp_47_ram[3433] = 4;
    exp_47_ram[3434] = 196;
    exp_47_ram[3435] = 79;
    exp_47_ram[3436] = 5;
    exp_47_ram[3437] = 244;
    exp_47_ram[3438] = 180;
    exp_47_ram[3439] = 7;
    exp_47_ram[3440] = 144;
    exp_47_ram[3441] = 231;
    exp_47_ram[3442] = 196;
    exp_47_ram[3443] = 7;
    exp_47_ram[3444] = 39;
    exp_47_ram[3445] = 231;
    exp_47_ram[3446] = 23;
    exp_47_ram[3447] = 244;
    exp_47_ram[3448] = 180;
    exp_47_ram[3449] = 196;
    exp_47_ram[3450] = 247;
    exp_47_ram[3451] = 7;
    exp_47_ram[3452] = 244;
    exp_47_ram[3453] = 95;
    exp_47_ram[3454] = 0;
    exp_47_ram[3455] = 196;
    exp_47_ram[3456] = 7;
    exp_47_ram[3457] = 193;
    exp_47_ram[3458] = 129;
    exp_47_ram[3459] = 1;
    exp_47_ram[3460] = 0;
    exp_47_ram[3461] = 1;
    exp_47_ram[3462] = 17;
    exp_47_ram[3463] = 129;
    exp_47_ram[3464] = 1;
    exp_47_ram[3465] = 0;
    exp_47_ram[3466] = 199;
    exp_47_ram[3467] = 7;
    exp_47_ram[3468] = 31;
    exp_47_ram[3469] = 5;
    exp_47_ram[3470] = 7;
    exp_47_ram[3471] = 193;
    exp_47_ram[3472] = 129;
    exp_47_ram[3473] = 1;
    exp_47_ram[3474] = 0;
    exp_47_ram[3475] = 1;
    exp_47_ram[3476] = 17;
    exp_47_ram[3477] = 129;
    exp_47_ram[3478] = 33;
    exp_47_ram[3479] = 49;
    exp_47_ram[3480] = 1;
    exp_47_ram[3481] = 164;
    exp_47_ram[3482] = 223;
    exp_47_ram[3483] = 164;
    exp_47_ram[3484] = 180;
    exp_47_ram[3485] = 0;
    exp_47_ram[3486] = 223;
    exp_47_ram[3487] = 5;
    exp_47_ram[3488] = 5;
    exp_47_ram[3489] = 132;
    exp_47_ram[3490] = 196;
    exp_47_ram[3491] = 166;
    exp_47_ram[3492] = 7;
    exp_47_ram[3493] = 6;
    exp_47_ram[3494] = 182;
    exp_47_ram[3495] = 7;
    exp_47_ram[3496] = 6;
    exp_47_ram[3497] = 196;
    exp_47_ram[3498] = 6;
    exp_47_ram[3499] = 0;
    exp_47_ram[3500] = 9;
    exp_47_ram[3501] = 7;
    exp_47_ram[3502] = 198;
    exp_47_ram[3503] = 9;
    exp_47_ram[3504] = 7;
    exp_47_ram[3505] = 214;
    exp_47_ram[3506] = 9;
    exp_47_ram[3507] = 7;
    exp_47_ram[3508] = 215;
    exp_47_ram[3509] = 0;
    exp_47_ram[3510] = 7;
    exp_47_ram[3511] = 193;
    exp_47_ram[3512] = 129;
    exp_47_ram[3513] = 65;
    exp_47_ram[3514] = 1;
    exp_47_ram[3515] = 1;
    exp_47_ram[3516] = 0;
    exp_47_ram[3517] = 1;
    exp_47_ram[3518] = 17;
    exp_47_ram[3519] = 129;
    exp_47_ram[3520] = 1;
    exp_47_ram[3521] = 0;
    exp_47_ram[3522] = 135;
    exp_47_ram[3523] = 207;
    exp_47_ram[3524] = 0;
    exp_47_ram[3525] = 193;
    exp_47_ram[3526] = 129;
    exp_47_ram[3527] = 1;
    exp_47_ram[3528] = 0;
    exp_47_ram[3529] = 1;
    exp_47_ram[3530] = 17;
    exp_47_ram[3531] = 129;
    exp_47_ram[3532] = 1;
    exp_47_ram[3533] = 0;
    exp_47_ram[3534] = 135;
    exp_47_ram[3535] = 207;
    exp_47_ram[3536] = 16;
    exp_47_ram[3537] = 244;
    exp_47_ram[3538] = 4;
    exp_47_ram[3539] = 0;
    exp_47_ram[3540] = 132;
    exp_47_ram[3541] = 0;
    exp_47_ram[3542] = 135;
    exp_47_ram[3543] = 207;
    exp_47_ram[3544] = 192;
    exp_47_ram[3545] = 196;
    exp_47_ram[3546] = 23;
    exp_47_ram[3547] = 244;
    exp_47_ram[3548] = 0;
    exp_47_ram[3549] = 135;
    exp_47_ram[3550] = 7;
    exp_47_ram[3551] = 196;
    exp_47_ram[3552] = 15;
    exp_47_ram[3553] = 0;
    exp_47_ram[3554] = 7;
    exp_47_ram[3555] = 160;
    exp_47_ram[3556] = 247;
    exp_47_ram[3557] = 7;
    exp_47_ram[3558] = 95;
    exp_47_ram[3559] = 196;
    exp_47_ram[3560] = 240;
    exp_47_ram[3561] = 231;
    exp_47_ram[3562] = 192;
    exp_47_ram[3563] = 196;
    exp_47_ram[3564] = 23;
    exp_47_ram[3565] = 244;
    exp_47_ram[3566] = 0;
    exp_47_ram[3567] = 135;
    exp_47_ram[3568] = 7;
    exp_47_ram[3569] = 196;
    exp_47_ram[3570] = 143;
    exp_47_ram[3571] = 0;
    exp_47_ram[3572] = 7;
    exp_47_ram[3573] = 160;
    exp_47_ram[3574] = 247;
    exp_47_ram[3575] = 7;
    exp_47_ram[3576] = 223;
    exp_47_ram[3577] = 196;
    exp_47_ram[3578] = 16;
    exp_47_ram[3579] = 231;
    exp_47_ram[3580] = 132;
    exp_47_ram[3581] = 23;
    exp_47_ram[3582] = 244;
    exp_47_ram[3583] = 132;
    exp_47_ram[3584] = 144;
    exp_47_ram[3585] = 231;
    exp_47_ram[3586] = 0;
    exp_47_ram[3587] = 135;
    exp_47_ram[3588] = 7;
    exp_47_ram[3589] = 0;
    exp_47_ram[3590] = 143;
    exp_47_ram[3591] = 0;
    exp_47_ram[3592] = 193;
    exp_47_ram[3593] = 129;
    exp_47_ram[3594] = 1;
    exp_47_ram[3595] = 0;
    exp_47_ram[3596] = 1;
    exp_47_ram[3597] = 17;
    exp_47_ram[3598] = 129;
    exp_47_ram[3599] = 33;
    exp_47_ram[3600] = 49;
    exp_47_ram[3601] = 65;
    exp_47_ram[3602] = 81;
    exp_47_ram[3603] = 97;
    exp_47_ram[3604] = 113;
    exp_47_ram[3605] = 129;
    exp_47_ram[3606] = 145;
    exp_47_ram[3607] = 161;
    exp_47_ram[3608] = 177;
    exp_47_ram[3609] = 1;
    exp_47_ram[3610] = 16;
    exp_47_ram[3611] = 244;
    exp_47_ram[3612] = 16;
    exp_47_ram[3613] = 0;
    exp_47_ram[3614] = 228;
    exp_47_ram[3615] = 244;
    exp_47_ram[3616] = 95;
    exp_47_ram[3617] = 164;
    exp_47_ram[3618] = 180;
    exp_47_ram[3619] = 4;
    exp_47_ram[3620] = 0;
    exp_47_ram[3621] = 196;
    exp_47_ram[3622] = 52;
    exp_47_ram[3623] = 135;
    exp_47_ram[3624] = 247;
    exp_47_ram[3625] = 244;
    exp_47_ram[3626] = 196;
    exp_47_ram[3627] = 52;
    exp_47_ram[3628] = 135;
    exp_47_ram[3629] = 247;
    exp_47_ram[3630] = 244;
    exp_47_ram[3631] = 196;
    exp_47_ram[3632] = 52;
    exp_47_ram[3633] = 135;
    exp_47_ram[3634] = 247;
    exp_47_ram[3635] = 244;
    exp_47_ram[3636] = 196;
    exp_47_ram[3637] = 52;
    exp_47_ram[3638] = 135;
    exp_47_ram[3639] = 247;
    exp_47_ram[3640] = 244;
    exp_47_ram[3641] = 196;
    exp_47_ram[3642] = 71;
    exp_47_ram[3643] = 244;
    exp_47_ram[3644] = 95;
    exp_47_ram[3645] = 5;
    exp_47_ram[3646] = 5;
    exp_47_ram[3647] = 4;
    exp_47_ram[3648] = 68;
    exp_47_ram[3649] = 166;
    exp_47_ram[3650] = 7;
    exp_47_ram[3651] = 6;
    exp_47_ram[3652] = 182;
    exp_47_ram[3653] = 7;
    exp_47_ram[3654] = 6;
    exp_47_ram[3655] = 0;
    exp_47_ram[3656] = 6;
    exp_47_ram[3657] = 212;
    exp_47_ram[3658] = 4;
    exp_47_ram[3659] = 132;
    exp_47_ram[3660] = 196;
    exp_47_ram[3661] = 5;
    exp_47_ram[3662] = 7;
    exp_47_ram[3663] = 198;
    exp_47_ram[3664] = 5;
    exp_47_ram[3665] = 7;
    exp_47_ram[3666] = 214;
    exp_47_ram[3667] = 5;
    exp_47_ram[3668] = 7;
    exp_47_ram[3669] = 215;
    exp_47_ram[3670] = 196;
    exp_47_ram[3671] = 0;
    exp_47_ram[3672] = 199;
    exp_47_ram[3673] = 79;
    exp_47_ram[3674] = 223;
    exp_47_ram[3675] = 164;
    exp_47_ram[3676] = 180;
    exp_47_ram[3677] = 4;
    exp_47_ram[3678] = 0;
    exp_47_ram[3679] = 4;
    exp_47_ram[3680] = 68;
    exp_47_ram[3681] = 52;
    exp_47_ram[3682] = 134;
    exp_47_ram[3683] = 215;
    exp_47_ram[3684] = 0;
    exp_47_ram[3685] = 215;
    exp_47_ram[3686] = 214;
    exp_47_ram[3687] = 52;
    exp_47_ram[3688] = 134;
    exp_47_ram[3689] = 215;
    exp_47_ram[3690] = 215;
    exp_47_ram[3691] = 5;
    exp_47_ram[3692] = 54;
    exp_47_ram[3693] = 7;
    exp_47_ram[3694] = 36;
    exp_47_ram[3695] = 52;
    exp_47_ram[3696] = 4;
    exp_47_ram[3697] = 68;
    exp_47_ram[3698] = 52;
    exp_47_ram[3699] = 134;
    exp_47_ram[3700] = 215;
    exp_47_ram[3701] = 0;
    exp_47_ram[3702] = 215;
    exp_47_ram[3703] = 214;
    exp_47_ram[3704] = 52;
    exp_47_ram[3705] = 134;
    exp_47_ram[3706] = 215;
    exp_47_ram[3707] = 215;
    exp_47_ram[3708] = 5;
    exp_47_ram[3709] = 86;
    exp_47_ram[3710] = 7;
    exp_47_ram[3711] = 68;
    exp_47_ram[3712] = 84;
    exp_47_ram[3713] = 4;
    exp_47_ram[3714] = 68;
    exp_47_ram[3715] = 52;
    exp_47_ram[3716] = 134;
    exp_47_ram[3717] = 215;
    exp_47_ram[3718] = 0;
    exp_47_ram[3719] = 215;
    exp_47_ram[3720] = 214;
    exp_47_ram[3721] = 52;
    exp_47_ram[3722] = 134;
    exp_47_ram[3723] = 215;
    exp_47_ram[3724] = 215;
    exp_47_ram[3725] = 5;
    exp_47_ram[3726] = 118;
    exp_47_ram[3727] = 7;
    exp_47_ram[3728] = 100;
    exp_47_ram[3729] = 116;
    exp_47_ram[3730] = 4;
    exp_47_ram[3731] = 68;
    exp_47_ram[3732] = 52;
    exp_47_ram[3733] = 134;
    exp_47_ram[3734] = 215;
    exp_47_ram[3735] = 0;
    exp_47_ram[3736] = 215;
    exp_47_ram[3737] = 214;
    exp_47_ram[3738] = 52;
    exp_47_ram[3739] = 134;
    exp_47_ram[3740] = 215;
    exp_47_ram[3741] = 215;
    exp_47_ram[3742] = 5;
    exp_47_ram[3743] = 150;
    exp_47_ram[3744] = 7;
    exp_47_ram[3745] = 132;
    exp_47_ram[3746] = 148;
    exp_47_ram[3747] = 196;
    exp_47_ram[3748] = 71;
    exp_47_ram[3749] = 244;
    exp_47_ram[3750] = 223;
    exp_47_ram[3751] = 5;
    exp_47_ram[3752] = 5;
    exp_47_ram[3753] = 4;
    exp_47_ram[3754] = 68;
    exp_47_ram[3755] = 166;
    exp_47_ram[3756] = 7;
    exp_47_ram[3757] = 6;
    exp_47_ram[3758] = 182;
    exp_47_ram[3759] = 7;
    exp_47_ram[3760] = 6;
    exp_47_ram[3761] = 0;
    exp_47_ram[3762] = 6;
    exp_47_ram[3763] = 212;
    exp_47_ram[3764] = 4;
    exp_47_ram[3765] = 4;
    exp_47_ram[3766] = 68;
    exp_47_ram[3767] = 5;
    exp_47_ram[3768] = 7;
    exp_47_ram[3769] = 198;
    exp_47_ram[3770] = 5;
    exp_47_ram[3771] = 7;
    exp_47_ram[3772] = 214;
    exp_47_ram[3773] = 5;
    exp_47_ram[3774] = 7;
    exp_47_ram[3775] = 215;
    exp_47_ram[3776] = 196;
    exp_47_ram[3777] = 0;
    exp_47_ram[3778] = 135;
    exp_47_ram[3779] = 207;
    exp_47_ram[3780] = 79;
    exp_47_ram[3781] = 164;
    exp_47_ram[3782] = 180;
    exp_47_ram[3783] = 4;
    exp_47_ram[3784] = 0;
    exp_47_ram[3785] = 196;
    exp_47_ram[3786] = 52;
    exp_47_ram[3787] = 135;
    exp_47_ram[3788] = 247;
    exp_47_ram[3789] = 244;
    exp_47_ram[3790] = 196;
    exp_47_ram[3791] = 52;
    exp_47_ram[3792] = 135;
    exp_47_ram[3793] = 247;
    exp_47_ram[3794] = 244;
    exp_47_ram[3795] = 196;
    exp_47_ram[3796] = 52;
    exp_47_ram[3797] = 135;
    exp_47_ram[3798] = 247;
    exp_47_ram[3799] = 244;
    exp_47_ram[3800] = 196;
    exp_47_ram[3801] = 52;
    exp_47_ram[3802] = 135;
    exp_47_ram[3803] = 247;
    exp_47_ram[3804] = 244;
    exp_47_ram[3805] = 196;
    exp_47_ram[3806] = 71;
    exp_47_ram[3807] = 244;
    exp_47_ram[3808] = 79;
    exp_47_ram[3809] = 5;
    exp_47_ram[3810] = 5;
    exp_47_ram[3811] = 4;
    exp_47_ram[3812] = 68;
    exp_47_ram[3813] = 166;
    exp_47_ram[3814] = 7;
    exp_47_ram[3815] = 6;
    exp_47_ram[3816] = 182;
    exp_47_ram[3817] = 7;
    exp_47_ram[3818] = 6;
    exp_47_ram[3819] = 0;
    exp_47_ram[3820] = 6;
    exp_47_ram[3821] = 212;
    exp_47_ram[3822] = 4;
    exp_47_ram[3823] = 132;
    exp_47_ram[3824] = 196;
    exp_47_ram[3825] = 5;
    exp_47_ram[3826] = 7;
    exp_47_ram[3827] = 198;
    exp_47_ram[3828] = 5;
    exp_47_ram[3829] = 7;
    exp_47_ram[3830] = 214;
    exp_47_ram[3831] = 5;
    exp_47_ram[3832] = 7;
    exp_47_ram[3833] = 215;
    exp_47_ram[3834] = 196;
    exp_47_ram[3835] = 0;
    exp_47_ram[3836] = 71;
    exp_47_ram[3837] = 79;
    exp_47_ram[3838] = 207;
    exp_47_ram[3839] = 164;
    exp_47_ram[3840] = 180;
    exp_47_ram[3841] = 4;
    exp_47_ram[3842] = 0;
    exp_47_ram[3843] = 4;
    exp_47_ram[3844] = 68;
    exp_47_ram[3845] = 52;
    exp_47_ram[3846] = 134;
    exp_47_ram[3847] = 0;
    exp_47_ram[3848] = 7;
    exp_47_ram[3849] = 7;
    exp_47_ram[3850] = 79;
    exp_47_ram[3851] = 5;
    exp_47_ram[3852] = 5;
    exp_47_ram[3853] = 228;
    exp_47_ram[3854] = 244;
    exp_47_ram[3855] = 4;
    exp_47_ram[3856] = 68;
    exp_47_ram[3857] = 52;
    exp_47_ram[3858] = 134;
    exp_47_ram[3859] = 0;
    exp_47_ram[3860] = 7;
    exp_47_ram[3861] = 7;
    exp_47_ram[3862] = 79;
    exp_47_ram[3863] = 5;
    exp_47_ram[3864] = 5;
    exp_47_ram[3865] = 228;
    exp_47_ram[3866] = 244;
    exp_47_ram[3867] = 4;
    exp_47_ram[3868] = 68;
    exp_47_ram[3869] = 52;
    exp_47_ram[3870] = 134;
    exp_47_ram[3871] = 0;
    exp_47_ram[3872] = 7;
    exp_47_ram[3873] = 7;
    exp_47_ram[3874] = 79;
    exp_47_ram[3875] = 5;
    exp_47_ram[3876] = 5;
    exp_47_ram[3877] = 228;
    exp_47_ram[3878] = 244;
    exp_47_ram[3879] = 4;
    exp_47_ram[3880] = 68;
    exp_47_ram[3881] = 52;
    exp_47_ram[3882] = 134;
    exp_47_ram[3883] = 0;
    exp_47_ram[3884] = 7;
    exp_47_ram[3885] = 7;
    exp_47_ram[3886] = 79;
    exp_47_ram[3887] = 5;
    exp_47_ram[3888] = 5;
    exp_47_ram[3889] = 228;
    exp_47_ram[3890] = 244;
    exp_47_ram[3891] = 196;
    exp_47_ram[3892] = 71;
    exp_47_ram[3893] = 244;
    exp_47_ram[3894] = 207;
    exp_47_ram[3895] = 5;
    exp_47_ram[3896] = 5;
    exp_47_ram[3897] = 4;
    exp_47_ram[3898] = 68;
    exp_47_ram[3899] = 166;
    exp_47_ram[3900] = 7;
    exp_47_ram[3901] = 6;
    exp_47_ram[3902] = 182;
    exp_47_ram[3903] = 7;
    exp_47_ram[3904] = 6;
    exp_47_ram[3905] = 0;
    exp_47_ram[3906] = 6;
    exp_47_ram[3907] = 6;
    exp_47_ram[3908] = 0;
    exp_47_ram[3909] = 13;
    exp_47_ram[3910] = 7;
    exp_47_ram[3911] = 198;
    exp_47_ram[3912] = 13;
    exp_47_ram[3913] = 7;
    exp_47_ram[3914] = 214;
    exp_47_ram[3915] = 13;
    exp_47_ram[3916] = 7;
    exp_47_ram[3917] = 215;
    exp_47_ram[3918] = 196;
    exp_47_ram[3919] = 0;
    exp_47_ram[3920] = 199;
    exp_47_ram[3921] = 79;
    exp_47_ram[3922] = 0;
    exp_47_ram[3923] = 193;
    exp_47_ram[3924] = 129;
    exp_47_ram[3925] = 65;
    exp_47_ram[3926] = 1;
    exp_47_ram[3927] = 193;
    exp_47_ram[3928] = 129;
    exp_47_ram[3929] = 65;
    exp_47_ram[3930] = 1;
    exp_47_ram[3931] = 193;
    exp_47_ram[3932] = 129;
    exp_47_ram[3933] = 65;
    exp_47_ram[3934] = 1;
    exp_47_ram[3935] = 1;
    exp_47_ram[3936] = 0;
    exp_47_ram[3937] = 1;
    exp_47_ram[3938] = 17;
    exp_47_ram[3939] = 129;
    exp_47_ram[3940] = 33;
    exp_47_ram[3941] = 49;
    exp_47_ram[3942] = 65;
    exp_47_ram[3943] = 81;
    exp_47_ram[3944] = 1;
    exp_47_ram[3945] = 0;
    exp_47_ram[3946] = 71;
    exp_47_ram[3947] = 207;
    exp_47_ram[3948] = 95;
    exp_47_ram[3949] = 5;
    exp_47_ram[3950] = 71;
    exp_47_ram[3951] = 244;
    exp_47_ram[3952] = 0;
    exp_47_ram[3953] = 199;
    exp_47_ram[3954] = 15;
    exp_47_ram[3955] = 159;
    exp_47_ram[3956] = 5;
    exp_47_ram[3957] = 247;
    exp_47_ram[3958] = 244;
    exp_47_ram[3959] = 0;
    exp_47_ram[3960] = 71;
    exp_47_ram[3961] = 79;
    exp_47_ram[3962] = 223;
    exp_47_ram[3963] = 5;
    exp_47_ram[3964] = 244;
    exp_47_ram[3965] = 0;
    exp_47_ram[3966] = 199;
    exp_47_ram[3967] = 207;
    exp_47_ram[3968] = 95;
    exp_47_ram[3969] = 5;
    exp_47_ram[3970] = 244;
    exp_47_ram[3971] = 0;
    exp_47_ram[3972] = 71;
    exp_47_ram[3973] = 79;
    exp_47_ram[3974] = 207;
    exp_47_ram[3975] = 5;
    exp_47_ram[3976] = 244;
    exp_47_ram[3977] = 112;
    exp_47_ram[3978] = 244;
    exp_47_ram[3979] = 16;
    exp_47_ram[3980] = 244;
    exp_47_ram[3981] = 4;
    exp_47_ram[3982] = 7;
    exp_47_ram[3983] = 31;
    exp_47_ram[3984] = 5;
    exp_47_ram[3985] = 5;
    exp_47_ram[3986] = 228;
    exp_47_ram[3987] = 244;
    exp_47_ram[3988] = 4;
    exp_47_ram[3989] = 7;
    exp_47_ram[3990] = 95;
    exp_47_ram[3991] = 5;
    exp_47_ram[3992] = 7;
    exp_47_ram[3993] = 31;
    exp_47_ram[3994] = 132;
    exp_47_ram[3995] = 7;
    exp_47_ram[3996] = 207;
    exp_47_ram[3997] = 5;
    exp_47_ram[3998] = 7;
    exp_47_ram[3999] = 159;
    exp_47_ram[4000] = 132;
    exp_47_ram[4001] = 196;
    exp_47_ram[4002] = 7;
    exp_47_ram[4003] = 7;
    exp_47_ram[4004] = 95;
    exp_47_ram[4005] = 0;
    exp_47_ram[4006] = 159;
    exp_47_ram[4007] = 5;
    exp_47_ram[4008] = 5;
    exp_47_ram[4009] = 228;
    exp_47_ram[4010] = 244;
    exp_47_ram[4011] = 132;
    exp_47_ram[4012] = 7;
    exp_47_ram[4013] = 143;
    exp_47_ram[4014] = 5;
    exp_47_ram[4015] = 7;
    exp_47_ram[4016] = 95;
    exp_47_ram[4017] = 15;
    exp_47_ram[4018] = 164;
    exp_47_ram[4019] = 180;
    exp_47_ram[4020] = 4;
    exp_47_ram[4021] = 128;
    exp_47_ram[4022] = 0;
    exp_47_ram[4023] = 143;
    exp_47_ram[4024] = 5;
    exp_47_ram[4025] = 5;
    exp_47_ram[4026] = 132;
    exp_47_ram[4027] = 196;
    exp_47_ram[4028] = 7;
    exp_47_ram[4029] = 7;
    exp_47_ram[4030] = 15;
    exp_47_ram[4031] = 5;
    exp_47_ram[4032] = 5;
    exp_47_ram[4033] = 0;
    exp_47_ram[4034] = 7;
    exp_47_ram[4035] = 7;
    exp_47_ram[4036] = 79;
    exp_47_ram[4037] = 5;
    exp_47_ram[4038] = 5;
    exp_47_ram[4039] = 7;
    exp_47_ram[4040] = 7;
    exp_47_ram[4041] = 10;
    exp_47_ram[4042] = 10;
    exp_47_ram[4043] = 79;
    exp_47_ram[4044] = 5;
    exp_47_ram[4045] = 7;
    exp_47_ram[4046] = 0;
    exp_47_ram[4047] = 7;
    exp_47_ram[4048] = 7;
    exp_47_ram[4049] = 0;
    exp_47_ram[4050] = 132;
    exp_47_ram[4051] = 196;
    exp_47_ram[4052] = 38;
    exp_47_ram[4053] = 7;
    exp_47_ram[4054] = 197;
    exp_47_ram[4055] = 54;
    exp_47_ram[4056] = 245;
    exp_47_ram[4057] = 6;
    exp_47_ram[4058] = 228;
    exp_47_ram[4059] = 244;
    exp_47_ram[4060] = 0;
    exp_47_ram[4061] = 223;
    exp_47_ram[4062] = 5;
    exp_47_ram[4063] = 5;
    exp_47_ram[4064] = 228;
    exp_47_ram[4065] = 244;
    exp_47_ram[4066] = 132;
    exp_47_ram[4067] = 7;
    exp_47_ram[4068] = 207;
    exp_47_ram[4069] = 5;
    exp_47_ram[4070] = 7;
    exp_47_ram[4071] = 159;
    exp_47_ram[4072] = 68;
    exp_47_ram[4073] = 23;
    exp_47_ram[4074] = 244;
    exp_47_ram[4075] = 68;
    exp_47_ram[4076] = 48;
    exp_47_ram[4077] = 231;
    exp_47_ram[4078] = 0;
    exp_47_ram[4079] = 0;
    exp_47_ram[4080] = 193;
    exp_47_ram[4081] = 129;
    exp_47_ram[4082] = 65;
    exp_47_ram[4083] = 1;
    exp_47_ram[4084] = 193;
    exp_47_ram[4085] = 129;
    exp_47_ram[4086] = 1;
    exp_47_ram[4087] = 0;
    exp_47_ram[4088] = 1;
    exp_47_ram[4089] = 17;
    exp_47_ram[4090] = 129;
    exp_47_ram[4091] = 1;
    exp_47_ram[4092] = 0;
    exp_47_ram[4093] = 7;
    exp_47_ram[4094] = 31;
    exp_47_ram[4095] = 0;
    exp_47_ram[4096] = 7;
    exp_47_ram[4097] = 95;
    exp_47_ram[4098] = 0;
    exp_47_ram[4099] = 71;
    exp_47_ram[4100] = 159;
    exp_47_ram[4101] = 0;
    exp_47_ram[4102] = 135;
    exp_47_ram[4103] = 223;
    exp_47_ram[4104] = 0;
    exp_47_ram[4105] = 7;
    exp_47_ram[4106] = 31;
    exp_47_ram[4107] = 31;
    exp_47_ram[4108] = 5;
    exp_47_ram[4109] = 244;
    exp_47_ram[4110] = 244;
    exp_47_ram[4111] = 64;
    exp_47_ram[4112] = 231;
    exp_47_ram[4113] = 64;
    exp_47_ram[4114] = 247;
    exp_47_ram[4115] = 48;
    exp_47_ram[4116] = 231;
    exp_47_ram[4117] = 48;
    exp_47_ram[4118] = 247;
    exp_47_ram[4119] = 16;
    exp_47_ram[4120] = 231;
    exp_47_ram[4121] = 32;
    exp_47_ram[4122] = 231;
    exp_47_ram[4123] = 64;
    exp_47_ram[4124] = 79;
    exp_47_ram[4125] = 192;
    exp_47_ram[4126] = 207;
    exp_47_ram[4127] = 64;
    exp_47_ram[4128] = 15;
    exp_47_ram[4129] = 192;
    exp_47_ram[4130] = 223;
    exp_47_ram[4131] = 0;
    exp_47_ram[4132] = 31;
    exp_47_ram[4133] = 5;
    exp_47_ram[4134] = 5;
    exp_47_ram[4135] = 181;
    exp_47_ram[4136] = 1;
    exp_47_ram[4137] = 183;
    exp_47_ram[4138] = 7;
    exp_47_ram[4139] = 5;
    exp_47_ram[4140] = 21;
    exp_47_ram[4141] = 245;
    exp_47_ram[4142] = 1;
    exp_47_ram[4143] = 0;
    exp_47_ram[4144] = 176;
    exp_47_ram[4145] = 245;
    exp_47_ram[4146] = 245;
    exp_47_ram[4147] = 223;
    exp_47_ram[4148] = 250;
    exp_47_ram[4149] = 0;
    exp_47_ram[4150] = 0;
    exp_47_ram[4151] = 0;
    exp_47_ram[4152] = 0;
    exp_47_ram[4153] = 0;
    exp_47_ram[4154] = 0;
    exp_47_ram[4155] = 0;
    exp_47_ram[4156] = 0;
    exp_47_ram[4157] = 0;
    exp_47_ram[4158] = 0;
    exp_47_ram[4159] = 0;
    exp_47_ram[4160] = 0;
    exp_47_ram[4161] = 0;
    exp_47_ram[4162] = 0;
    exp_47_ram[4163] = 0;
    exp_47_ram[4164] = 0;
    exp_47_ram[4165] = 0;
    exp_47_ram[4166] = 0;
    exp_47_ram[4167] = 0;
    exp_47_ram[4168] = 0;
    exp_47_ram[4169] = 0;
    exp_47_ram[4170] = 0;
    exp_47_ram[4171] = 0;
    exp_47_ram[4172] = 0;
    exp_47_ram[4173] = 0;
    exp_47_ram[4174] = 0;
    exp_47_ram[4175] = 0;
    exp_47_ram[4176] = 0;
    exp_47_ram[4177] = 0;
    exp_47_ram[4178] = 0;
    exp_47_ram[4179] = 0;
    exp_47_ram[4180] = 0;
    exp_47_ram[4181] = 0;
    exp_47_ram[4182] = 0;
    exp_47_ram[4183] = 0;
    exp_47_ram[4184] = 0;
    exp_47_ram[4185] = 0;
    exp_47_ram[4186] = 0;
    exp_47_ram[4187] = 0;
    exp_47_ram[4188] = 0;
    exp_47_ram[4189] = 0;
    exp_47_ram[4190] = 0;
    exp_47_ram[4191] = 0;
    exp_47_ram[4192] = 0;
    exp_47_ram[4193] = 0;
    exp_47_ram[4194] = 0;
    exp_47_ram[4195] = 0;
    exp_47_ram[4196] = 0;
    exp_47_ram[4197] = 0;
    exp_47_ram[4198] = 0;
    exp_47_ram[4199] = 0;
    exp_47_ram[4200] = 0;
    exp_47_ram[4201] = 0;
    exp_47_ram[4202] = 0;
    exp_47_ram[4203] = 0;
    exp_47_ram[4204] = 0;
    exp_47_ram[4205] = 0;
    exp_47_ram[4206] = 0;
    exp_47_ram[4207] = 0;
    exp_47_ram[4208] = 0;
    exp_47_ram[4209] = 0;
    exp_47_ram[4210] = 0;
    exp_47_ram[4211] = 0;
    exp_47_ram[4212] = 0;
    exp_47_ram[4213] = 0;
    exp_47_ram[4214] = 0;
    exp_47_ram[4215] = 0;
    exp_47_ram[4216] = 0;
    exp_47_ram[4217] = 0;
    exp_47_ram[4218] = 0;
    exp_47_ram[4219] = 0;
    exp_47_ram[4220] = 0;
    exp_47_ram[4221] = 0;
    exp_47_ram[4222] = 0;
    exp_47_ram[4223] = 0;
    exp_47_ram[4224] = 0;
    exp_47_ram[4225] = 0;
    exp_47_ram[4226] = 0;
    exp_47_ram[4227] = 0;
    exp_47_ram[4228] = 0;
    exp_47_ram[4229] = 0;
    exp_47_ram[4230] = 0;
    exp_47_ram[4231] = 0;
    exp_47_ram[4232] = 0;
    exp_47_ram[4233] = 0;
    exp_47_ram[4234] = 0;
    exp_47_ram[4235] = 0;
    exp_47_ram[4236] = 0;
    exp_47_ram[4237] = 0;
    exp_47_ram[4238] = 0;
    exp_47_ram[4239] = 0;
    exp_47_ram[4240] = 0;
    exp_47_ram[4241] = 0;
    exp_47_ram[4242] = 0;
    exp_47_ram[4243] = 0;
    exp_47_ram[4244] = 0;
    exp_47_ram[4245] = 0;
    exp_47_ram[4246] = 0;
    exp_47_ram[4247] = 0;
    exp_47_ram[4248] = 0;
    exp_47_ram[4249] = 0;
    exp_47_ram[4250] = 0;
    exp_47_ram[4251] = 0;
    exp_47_ram[4252] = 0;
    exp_47_ram[4253] = 0;
    exp_47_ram[4254] = 0;
    exp_47_ram[4255] = 0;
    exp_47_ram[4256] = 0;
    exp_47_ram[4257] = 0;
    exp_47_ram[4258] = 0;
    exp_47_ram[4259] = 0;
    exp_47_ram[4260] = 0;
    exp_47_ram[4261] = 0;
    exp_47_ram[4262] = 0;
    exp_47_ram[4263] = 0;
    exp_47_ram[4264] = 0;
    exp_47_ram[4265] = 0;
    exp_47_ram[4266] = 0;
    exp_47_ram[4267] = 0;
    exp_47_ram[4268] = 0;
    exp_47_ram[4269] = 0;
    exp_47_ram[4270] = 0;
    exp_47_ram[4271] = 0;
    exp_47_ram[4272] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 81;
    exp_40_ram[32] = 1;
    exp_40_ram[33] = 48;
    exp_40_ram[34] = 0;
    exp_40_ram[35] = 8;
    exp_40_ram[36] = 135;
    exp_40_ram[37] = 8;
    exp_40_ram[38] = 133;
    exp_40_ram[39] = 131;
    exp_40_ram[40] = 148;
    exp_40_ram[41] = 22;
    exp_40_ram[42] = 134;
    exp_40_ram[43] = 246;
    exp_40_ram[44] = 7;
    exp_40_ram[45] = 120;
    exp_40_ram[46] = 7;
    exp_40_ram[47] = 55;
    exp_40_ram[48] = 23;
    exp_40_ram[49] = 85;
    exp_40_ram[50] = 134;
    exp_40_ram[51] = 198;
    exp_40_ram[52] = 5;
    exp_40_ram[53] = 135;
    exp_40_ram[54] = 6;
    exp_40_ram[55] = 12;
    exp_40_ram[56] = 149;
    exp_40_ram[57] = 215;
    exp_40_ram[58] = 24;
    exp_40_ram[59] = 101;
    exp_40_ram[60] = 147;
    exp_40_ram[61] = 88;
    exp_40_ram[62] = 214;
    exp_40_ram[63] = 22;
    exp_40_ram[64] = 86;
    exp_40_ram[65] = 87;
    exp_40_ram[66] = 247;
    exp_40_ram[67] = 133;
    exp_40_ram[68] = 5;
    exp_40_ram[69] = 23;
    exp_40_ram[70] = 103;
    exp_40_ram[71] = 254;
    exp_40_ram[72] = 135;
    exp_40_ram[73] = 133;
    exp_40_ram[74] = 232;
    exp_40_ram[75] = 246;
    exp_40_ram[76] = 133;
    exp_40_ram[77] = 135;
    exp_40_ram[78] = 135;
    exp_40_ram[79] = 247;
    exp_40_ram[80] = 19;
    exp_40_ram[81] = 83;
    exp_40_ram[82] = 215;
    exp_40_ram[83] = 23;
    exp_40_ram[84] = 99;
    exp_40_ram[85] = 6;
    exp_40_ram[86] = 134;
    exp_40_ram[87] = 124;
    exp_40_ram[88] = 3;
    exp_40_ram[89] = 134;
    exp_40_ram[90] = 102;
    exp_40_ram[91] = 116;
    exp_40_ram[92] = 134;
    exp_40_ram[93] = 21;
    exp_40_ram[94] = 101;
    exp_40_ram[95] = 5;
    exp_40_ram[96] = 0;
    exp_40_ram[97] = 5;
    exp_40_ram[98] = 7;
    exp_40_ram[99] = 108;
    exp_40_ram[100] = 7;
    exp_40_ram[101] = 240;
    exp_40_ram[102] = 22;
    exp_40_ram[103] = 7;
    exp_40_ram[104] = 88;
    exp_40_ram[105] = 7;
    exp_40_ram[106] = 112;
    exp_40_ram[107] = 7;
    exp_40_ram[108] = 116;
    exp_40_ram[109] = 5;
    exp_40_ram[110] = 87;
    exp_40_ram[111] = 134;
    exp_40_ram[112] = 199;
    exp_40_ram[113] = 6;
    exp_40_ram[114] = 7;
    exp_40_ram[115] = 6;
    exp_40_ram[116] = 22;
    exp_40_ram[117] = 135;
    exp_40_ram[118] = 5;
    exp_40_ram[119] = 88;
    exp_40_ram[120] = 22;
    exp_40_ram[121] = 86;
    exp_40_ram[122] = 87;
    exp_40_ram[123] = 246;
    exp_40_ram[124] = 215;
    exp_40_ram[125] = 150;
    exp_40_ram[126] = 231;
    exp_40_ram[127] = 14;
    exp_40_ram[128] = 133;
    exp_40_ram[129] = 126;
    exp_40_ram[130] = 7;
    exp_40_ram[131] = 133;
    exp_40_ram[132] = 104;
    exp_40_ram[133] = 118;
    exp_40_ram[134] = 133;
    exp_40_ram[135] = 7;
    exp_40_ram[136] = 7;
    exp_40_ram[137] = 119;
    exp_40_ram[138] = 19;
    exp_40_ram[139] = 83;
    exp_40_ram[140] = 87;
    exp_40_ram[141] = 151;
    exp_40_ram[142] = 227;
    exp_40_ram[143] = 6;
    exp_40_ram[144] = 6;
    exp_40_ram[145] = 124;
    exp_40_ram[146] = 3;
    exp_40_ram[147] = 6;
    exp_40_ram[148] = 102;
    exp_40_ram[149] = 116;
    exp_40_ram[150] = 6;
    exp_40_ram[151] = 21;
    exp_40_ram[152] = 101;
    exp_40_ram[153] = 128;
    exp_40_ram[154] = 7;
    exp_40_ram[155] = 5;
    exp_40_ram[156] = 100;
    exp_40_ram[157] = 5;
    exp_40_ram[158] = 240;
    exp_40_ram[159] = 24;
    exp_40_ram[160] = 213;
    exp_40_ram[161] = 147;
    exp_40_ram[162] = 151;
    exp_40_ram[163] = 215;
    exp_40_ram[164] = 88;
    exp_40_ram[165] = 102;
    exp_40_ram[166] = 119;
    exp_40_ram[167] = 23;
    exp_40_ram[168] = 215;
    exp_40_ram[169] = 85;
    exp_40_ram[170] = 85;
    exp_40_ram[171] = 23;
    exp_40_ram[172] = 103;
    exp_40_ram[173] = 134;
    exp_40_ram[174] = 5;
    exp_40_ram[175] = 126;
    exp_40_ram[176] = 7;
    exp_40_ram[177] = 5;
    exp_40_ram[178] = 104;
    exp_40_ram[179] = 118;
    exp_40_ram[180] = 5;
    exp_40_ram[181] = 7;
    exp_40_ram[182] = 6;
    exp_40_ram[183] = 247;
    exp_40_ram[184] = 22;
    exp_40_ram[185] = 86;
    exp_40_ram[186] = 214;
    exp_40_ram[187] = 23;
    exp_40_ram[188] = 133;
    exp_40_ram[189] = 103;
    exp_40_ram[190] = 135;
    exp_40_ram[191] = 254;
    exp_40_ram[192] = 135;
    exp_40_ram[193] = 135;
    exp_40_ram[194] = 232;
    exp_40_ram[195] = 246;
    exp_40_ram[196] = 135;
    exp_40_ram[197] = 135;
    exp_40_ram[198] = 149;
    exp_40_ram[199] = 135;
    exp_40_ram[200] = 229;
    exp_40_ram[201] = 240;
    exp_40_ram[202] = 230;
    exp_40_ram[203] = 7;
    exp_40_ram[204] = 244;
    exp_40_ram[205] = 7;
    exp_40_ram[206] = 53;
    exp_40_ram[207] = 149;
    exp_40_ram[208] = 23;
    exp_40_ram[209] = 213;
    exp_40_ram[210] = 7;
    exp_40_ram[211] = 7;
    exp_40_ram[212] = 71;
    exp_40_ram[213] = 5;
    exp_40_ram[214] = 7;
    exp_40_ram[215] = 5;
    exp_40_ram[216] = 22;
    exp_40_ram[217] = 5;
    exp_40_ram[218] = 238;
    exp_40_ram[219] = 181;
    exp_40_ram[220] = 69;
    exp_40_ram[221] = 240;
    exp_40_ram[222] = 7;
    exp_40_ram[223] = 5;
    exp_40_ram[224] = 224;
    exp_40_ram[225] = 5;
    exp_40_ram[226] = 240;
    exp_40_ram[227] = 88;
    exp_40_ram[228] = 150;
    exp_40_ram[229] = 104;
    exp_40_ram[230] = 222;
    exp_40_ram[231] = 94;
    exp_40_ram[232] = 118;
    exp_40_ram[233] = 151;
    exp_40_ram[234] = 215;
    exp_40_ram[235] = 19;
    exp_40_ram[236] = 102;
    exp_40_ram[237] = 23;
    exp_40_ram[238] = 215;
    exp_40_ram[239] = 87;
    exp_40_ram[240] = 94;
    exp_40_ram[241] = 150;
    exp_40_ram[242] = 231;
    exp_40_ram[243] = 143;
    exp_40_ram[244] = 5;
    exp_40_ram[245] = 126;
    exp_40_ram[246] = 7;
    exp_40_ram[247] = 5;
    exp_40_ram[248] = 104;
    exp_40_ram[249] = 118;
    exp_40_ram[250] = 5;
    exp_40_ram[251] = 7;
    exp_40_ram[252] = 7;
    exp_40_ram[253] = 118;
    exp_40_ram[254] = 87;
    exp_40_ram[255] = 150;
    exp_40_ram[256] = 142;
    exp_40_ram[257] = 23;
    exp_40_ram[258] = 215;
    exp_40_ram[259] = 231;
    exp_40_ram[260] = 6;
    exp_40_ram[261] = 254;
    exp_40_ram[262] = 135;
    exp_40_ram[263] = 6;
    exp_40_ram[264] = 232;
    exp_40_ram[265] = 246;
    exp_40_ram[266] = 6;
    exp_40_ram[267] = 135;
    exp_40_ram[268] = 21;
    exp_40_ram[269] = 14;
    exp_40_ram[270] = 101;
    exp_40_ram[271] = 134;
    exp_40_ram[272] = 120;
    exp_40_ram[273] = 86;
    exp_40_ram[274] = 118;
    exp_40_ram[275] = 83;
    exp_40_ram[276] = 135;
    exp_40_ram[277] = 14;
    exp_40_ram[278] = 6;
    exp_40_ram[279] = 87;
    exp_40_ram[280] = 8;
    exp_40_ram[281] = 8;
    exp_40_ram[282] = 7;
    exp_40_ram[283] = 6;
    exp_40_ram[284] = 116;
    exp_40_ram[285] = 6;
    exp_40_ram[286] = 86;
    exp_40_ram[287] = 134;
    exp_40_ram[288] = 230;
    exp_40_ram[289] = 156;
    exp_40_ram[290] = 7;
    exp_40_ram[291] = 135;
    exp_40_ram[292] = 119;
    exp_40_ram[293] = 23;
    exp_40_ram[294] = 126;
    exp_40_ram[295] = 152;
    exp_40_ram[296] = 7;
    exp_40_ram[297] = 5;
    exp_40_ram[298] = 254;
    exp_40_ram[299] = 5;
    exp_40_ram[300] = 240;
    exp_40_ram[301] = 5;
    exp_40_ram[302] = 5;
    exp_40_ram[303] = 240;
    exp_40_ram[304] = 7;
    exp_40_ram[305] = 7;
    exp_40_ram[306] = 216;
    exp_40_ram[307] = 120;
    exp_40_ram[308] = 7;
    exp_40_ram[309] = 3;
    exp_40_ram[310] = 120;
    exp_40_ram[311] = 213;
    exp_40_ram[312] = 14;
    exp_40_ram[313] = 213;
    exp_40_ram[314] = 119;
    exp_40_ram[315] = 14;
    exp_40_ram[316] = 245;
    exp_40_ram[317] = 214;
    exp_40_ram[318] = 26;
    exp_40_ram[319] = 238;
    exp_40_ram[320] = 138;
    exp_40_ram[321] = 5;
    exp_40_ram[322] = 128;
    exp_40_ram[323] = 150;
    exp_40_ram[324] = 110;
    exp_40_ram[325] = 152;
    exp_40_ram[326] = 16;
    exp_40_ram[327] = 231;
    exp_40_ram[328] = 183;
    exp_40_ram[329] = 150;
    exp_40_ram[330] = 102;
    exp_40_ram[331] = 12;
    exp_40_ram[332] = 156;
    exp_40_ram[333] = 20;
    exp_40_ram[334] = 208;
    exp_40_ram[335] = 0;
    exp_40_ram[336] = 5;
    exp_40_ram[337] = 128;
    exp_40_ram[338] = 5;
    exp_40_ram[339] = 138;
    exp_40_ram[340] = 133;
    exp_40_ram[341] = 128;
    exp_40_ram[342] = 86;
    exp_40_ram[343] = 2;
    exp_40_ram[344] = 128;
    exp_40_ram[345] = 108;
    exp_40_ram[346] = 146;
    exp_40_ram[347] = 104;
    exp_40_ram[348] = 102;
    exp_40_ram[349] = 5;
    exp_40_ram[350] = 128;
    exp_40_ram[351] = 5;
    exp_40_ram[352] = 128;
    exp_40_ram[353] = 152;
    exp_40_ram[354] = 240;
    exp_40_ram[355] = 232;
    exp_40_ram[356] = 240;
    exp_40_ram[357] = 142;
    exp_40_ram[358] = 158;
    exp_40_ram[359] = 7;
    exp_40_ram[360] = 240;
    exp_40_ram[361] = 1;
    exp_40_ram[362] = 36;
    exp_40_ram[363] = 38;
    exp_40_ram[364] = 4;
    exp_40_ram[365] = 2;
    exp_40_ram[366] = 0;
    exp_40_ram[367] = 7;
    exp_40_ram[368] = 7;
    exp_40_ram[369] = 7;
    exp_40_ram[370] = 192;
    exp_40_ram[371] = 7;
    exp_40_ram[372] = 135;
    exp_40_ram[373] = 5;
    exp_40_ram[374] = 87;
    exp_40_ram[375] = 20;
    exp_40_ram[376] = 32;
    exp_40_ram[377] = 5;
    exp_40_ram[378] = 151;
    exp_40_ram[379] = 36;
    exp_40_ram[380] = 23;
    exp_40_ram[381] = 215;
    exp_40_ram[382] = 102;
    exp_40_ram[383] = 133;
    exp_40_ram[384] = 1;
    exp_40_ram[385] = 128;
    exp_40_ram[386] = 7;
    exp_40_ram[387] = 23;
    exp_40_ram[388] = 4;
    exp_40_ram[389] = 240;
    exp_40_ram[390] = 7;
    exp_40_ram[391] = 7;
    exp_40_ram[392] = 240;
    exp_40_ram[393] = 1;
    exp_40_ram[394] = 46;
    exp_40_ram[395] = 44;
    exp_40_ram[396] = 42;
    exp_40_ram[397] = 40;
    exp_40_ram[398] = 38;
    exp_40_ram[399] = 36;
    exp_40_ram[400] = 103;
    exp_40_ram[401] = 140;
    exp_40_ram[402] = 4;
    exp_40_ram[403] = 137;
    exp_40_ram[404] = 132;
    exp_40_ram[405] = 132;
    exp_40_ram[406] = 133;
    exp_40_ram[407] = 0;
    exp_40_ram[408] = 9;
    exp_40_ram[409] = 10;
    exp_40_ram[410] = 10;
    exp_40_ram[411] = 7;
    exp_40_ram[412] = 196;
    exp_40_ram[413] = 7;
    exp_40_ram[414] = 7;
    exp_40_ram[415] = 84;
    exp_40_ram[416] = 7;
    exp_40_ram[417] = 66;
    exp_40_ram[418] = 4;
    exp_40_ram[419] = 135;
    exp_40_ram[420] = 132;
    exp_40_ram[421] = 84;
    exp_40_ram[422] = 21;
    exp_40_ram[423] = 228;
    exp_40_ram[424] = 23;
    exp_40_ram[425] = 32;
    exp_40_ram[426] = 36;
    exp_40_ram[427] = 149;
    exp_40_ram[428] = 26;
    exp_40_ram[429] = 213;
    exp_40_ram[430] = 103;
    exp_40_ram[431] = 36;
    exp_40_ram[432] = 41;
    exp_40_ram[433] = 41;
    exp_40_ram[434] = 42;
    exp_40_ram[435] = 133;
    exp_40_ram[436] = 5;
    exp_40_ram[437] = 1;
    exp_40_ram[438] = 128;
    exp_40_ram[439] = 0;
    exp_40_ram[440] = 9;
    exp_40_ram[441] = 240;
    exp_40_ram[442] = 133;
    exp_40_ram[443] = 20;
    exp_40_ram[444] = 7;
    exp_40_ram[445] = 240;
    exp_40_ram[446] = 7;
    exp_40_ram[447] = 220;
    exp_40_ram[448] = 134;
    exp_40_ram[449] = 5;
    exp_40_ram[450] = 5;
    exp_40_ram[451] = 0;
    exp_40_ram[452] = 101;
    exp_40_ram[453] = 6;
    exp_40_ram[454] = 52;
    exp_40_ram[455] = 5;
    exp_40_ram[456] = 5;
    exp_40_ram[457] = 6;
    exp_40_ram[458] = 0;
    exp_40_ram[459] = 228;
    exp_40_ram[460] = 137;
    exp_40_ram[461] = 7;
    exp_40_ram[462] = 7;
    exp_40_ram[463] = 5;
    exp_40_ram[464] = 84;
    exp_40_ram[465] = 7;
    exp_40_ram[466] = 66;
    exp_40_ram[467] = 135;
    exp_40_ram[468] = 21;
    exp_40_ram[469] = 9;
    exp_40_ram[470] = 9;
    exp_40_ram[471] = 89;
    exp_40_ram[472] = 101;
    exp_40_ram[473] = 23;
    exp_40_ram[474] = 7;
    exp_40_ram[475] = 7;
    exp_40_ram[476] = 245;
    exp_40_ram[477] = 247;
    exp_40_ram[478] = 0;
    exp_40_ram[479] = 247;
    exp_40_ram[480] = 6;
    exp_40_ram[481] = 10;
    exp_40_ram[482] = 135;
    exp_40_ram[483] = 55;
    exp_40_ram[484] = 133;
    exp_40_ram[485] = 7;
    exp_40_ram[486] = 7;
    exp_40_ram[487] = 247;
    exp_40_ram[488] = 12;
    exp_40_ram[489] = 7;
    exp_40_ram[490] = 7;
    exp_40_ram[491] = 10;
    exp_40_ram[492] = 245;
    exp_40_ram[493] = 10;
    exp_40_ram[494] = 215;
    exp_40_ram[495] = 149;
    exp_40_ram[496] = 103;
    exp_40_ram[497] = 212;
    exp_40_ram[498] = 240;
    exp_40_ram[499] = 133;
    exp_40_ram[500] = 21;
    exp_40_ram[501] = 7;
    exp_40_ram[502] = 240;
    exp_40_ram[503] = 4;
    exp_40_ram[504] = 7;
    exp_40_ram[505] = 10;
    exp_40_ram[506] = 240;
    exp_40_ram[507] = 0;
    exp_40_ram[508] = 7;
    exp_40_ram[509] = 135;
    exp_40_ram[510] = 76;
    exp_40_ram[511] = 5;
    exp_40_ram[512] = 7;
    exp_40_ram[513] = 213;
    exp_40_ram[514] = 5;
    exp_40_ram[515] = 128;
    exp_40_ram[516] = 215;
    exp_40_ram[517] = 85;
    exp_40_ram[518] = 149;
    exp_40_ram[519] = 101;
    exp_40_ram[520] = 240;
    exp_40_ram[521] = 0;
    exp_40_ram[522] = 7;
    exp_40_ram[523] = 135;
    exp_40_ram[524] = 76;
    exp_40_ram[525] = 5;
    exp_40_ram[526] = 7;
    exp_40_ram[527] = 21;
    exp_40_ram[528] = 5;
    exp_40_ram[529] = 128;
    exp_40_ram[530] = 23;
    exp_40_ram[531] = 149;
    exp_40_ram[532] = 85;
    exp_40_ram[533] = 229;
    exp_40_ram[534] = 240;
    exp_40_ram[535] = 7;
    exp_40_ram[536] = 122;
    exp_40_ram[537] = 7;
    exp_40_ram[538] = 183;
    exp_40_ram[539] = 151;
    exp_40_ram[540] = 23;
    exp_40_ram[541] = 6;
    exp_40_ram[542] = 134;
    exp_40_ram[543] = 85;
    exp_40_ram[544] = 7;
    exp_40_ram[545] = 133;
    exp_40_ram[546] = 69;
    exp_40_ram[547] = 133;
    exp_40_ram[548] = 128;
    exp_40_ram[549] = 7;
    exp_40_ram[550] = 7;
    exp_40_ram[551] = 106;
    exp_40_ram[552] = 7;
    exp_40_ram[553] = 240;
    exp_40_ram[554] = 117;
    exp_40_ram[555] = 110;
    exp_40_ram[556] = 87;
    exp_40_ram[557] = 104;
    exp_40_ram[558] = 105;
    exp_40_ram[559] = 0;
    exp_40_ram[560] = 97;
    exp_40_ram[561] = 98;
    exp_40_ram[562] = 65;
    exp_40_ram[563] = 97;
    exp_40_ram[564] = 110;
    exp_40_ram[565] = 65;
    exp_40_ram[566] = 101;
    exp_40_ram[567] = 116;
    exp_40_ram[568] = 68;
    exp_40_ram[569] = 0;
    exp_40_ram[570] = 101;
    exp_40_ram[571] = 32;
    exp_40_ram[572] = 108;
    exp_40_ram[573] = 0;
    exp_40_ram[574] = 117;
    exp_40_ram[575] = 110;
    exp_40_ram[576] = 110;
    exp_40_ram[577] = 116;
    exp_40_ram[578] = 100;
    exp_40_ram[579] = 100;
    exp_40_ram[580] = 46;
    exp_40_ram[581] = 0;
    exp_40_ram[582] = 117;
    exp_40_ram[583] = 117;
    exp_40_ram[584] = 45;
    exp_40_ram[585] = 32;
    exp_40_ram[586] = 101;
    exp_40_ram[587] = 32;
    exp_40_ram[588] = 116;
    exp_40_ram[589] = 105;
    exp_40_ram[590] = 105;
    exp_40_ram[591] = 32;
    exp_40_ram[592] = 111;
    exp_40_ram[593] = 0;
    exp_40_ram[594] = 117;
    exp_40_ram[595] = 45;
    exp_40_ram[596] = 32;
    exp_40_ram[597] = 101;
    exp_40_ram[598] = 32;
    exp_40_ram[599] = 116;
    exp_40_ram[600] = 105;
    exp_40_ram[601] = 105;
    exp_40_ram[602] = 32;
    exp_40_ram[603] = 111;
    exp_40_ram[604] = 0;
    exp_40_ram[605] = 117;
    exp_40_ram[606] = 45;
    exp_40_ram[607] = 32;
    exp_40_ram[608] = 101;
    exp_40_ram[609] = 32;
    exp_40_ram[610] = 105;
    exp_40_ram[611] = 32;
    exp_40_ram[612] = 49;
    exp_40_ram[613] = 99;
    exp_40_ram[614] = 10;
    exp_40_ram[615] = 117;
    exp_40_ram[616] = 45;
    exp_40_ram[617] = 32;
    exp_40_ram[618] = 101;
    exp_40_ram[619] = 32;
    exp_40_ram[620] = 105;
    exp_40_ram[621] = 32;
    exp_40_ram[622] = 49;
    exp_40_ram[623] = 99;
    exp_40_ram[624] = 10;
    exp_40_ram[625] = 101;
    exp_40_ram[626] = 10;
    exp_40_ram[627] = 111;
    exp_40_ram[628] = 58;
    exp_40_ram[629] = 97;
    exp_40_ram[630] = 0;
    exp_40_ram[631] = 111;
    exp_40_ram[632] = 10;
    exp_40_ram[633] = 105;
    exp_40_ram[634] = 101;
    exp_40_ram[635] = 0;
    exp_40_ram[636] = 67;
    exp_40_ram[637] = 115;
    exp_40_ram[638] = 68;
    exp_40_ram[639] = 10;
    exp_40_ram[640] = 97;
    exp_40_ram[641] = 101;
    exp_40_ram[642] = 32;
    exp_40_ram[643] = 108;
    exp_40_ram[644] = 0;
    exp_40_ram[645] = 41;
    exp_40_ram[646] = 105;
    exp_40_ram[647] = 32;
    exp_40_ram[648] = 101;
    exp_40_ram[649] = 0;
    exp_40_ram[650] = 41;
    exp_40_ram[651] = 115;
    exp_40_ram[652] = 117;
    exp_40_ram[653] = 112;
    exp_40_ram[654] = 97;
    exp_40_ram[655] = 110;
    exp_40_ram[656] = 41;
    exp_40_ram[657] = 108;
    exp_40_ram[658] = 108;
    exp_40_ram[659] = 10;
    exp_40_ram[660] = 1;
    exp_40_ram[661] = 3;
    exp_40_ram[662] = 4;
    exp_40_ram[663] = 4;
    exp_40_ram[664] = 5;
    exp_40_ram[665] = 5;
    exp_40_ram[666] = 5;
    exp_40_ram[667] = 5;
    exp_40_ram[668] = 6;
    exp_40_ram[669] = 6;
    exp_40_ram[670] = 6;
    exp_40_ram[671] = 6;
    exp_40_ram[672] = 6;
    exp_40_ram[673] = 6;
    exp_40_ram[674] = 6;
    exp_40_ram[675] = 6;
    exp_40_ram[676] = 7;
    exp_40_ram[677] = 7;
    exp_40_ram[678] = 7;
    exp_40_ram[679] = 7;
    exp_40_ram[680] = 7;
    exp_40_ram[681] = 7;
    exp_40_ram[682] = 7;
    exp_40_ram[683] = 7;
    exp_40_ram[684] = 7;
    exp_40_ram[685] = 7;
    exp_40_ram[686] = 7;
    exp_40_ram[687] = 7;
    exp_40_ram[688] = 7;
    exp_40_ram[689] = 7;
    exp_40_ram[690] = 7;
    exp_40_ram[691] = 7;
    exp_40_ram[692] = 8;
    exp_40_ram[693] = 8;
    exp_40_ram[694] = 8;
    exp_40_ram[695] = 8;
    exp_40_ram[696] = 8;
    exp_40_ram[697] = 8;
    exp_40_ram[698] = 8;
    exp_40_ram[699] = 8;
    exp_40_ram[700] = 8;
    exp_40_ram[701] = 8;
    exp_40_ram[702] = 8;
    exp_40_ram[703] = 8;
    exp_40_ram[704] = 8;
    exp_40_ram[705] = 8;
    exp_40_ram[706] = 8;
    exp_40_ram[707] = 8;
    exp_40_ram[708] = 8;
    exp_40_ram[709] = 8;
    exp_40_ram[710] = 8;
    exp_40_ram[711] = 8;
    exp_40_ram[712] = 8;
    exp_40_ram[713] = 8;
    exp_40_ram[714] = 8;
    exp_40_ram[715] = 8;
    exp_40_ram[716] = 8;
    exp_40_ram[717] = 8;
    exp_40_ram[718] = 8;
    exp_40_ram[719] = 8;
    exp_40_ram[720] = 8;
    exp_40_ram[721] = 8;
    exp_40_ram[722] = 8;
    exp_40_ram[723] = 8;
    exp_40_ram[724] = 1;
    exp_40_ram[725] = 38;
    exp_40_ram[726] = 4;
    exp_40_ram[727] = 46;
    exp_40_ram[728] = 39;
    exp_40_ram[729] = 38;
    exp_40_ram[730] = 39;
    exp_40_ram[731] = 167;
    exp_40_ram[732] = 133;
    exp_40_ram[733] = 36;
    exp_40_ram[734] = 1;
    exp_40_ram[735] = 128;
    exp_40_ram[736] = 1;
    exp_40_ram[737] = 38;
    exp_40_ram[738] = 4;
    exp_40_ram[739] = 46;
    exp_40_ram[740] = 44;
    exp_40_ram[741] = 39;
    exp_40_ram[742] = 38;
    exp_40_ram[743] = 39;
    exp_40_ram[744] = 39;
    exp_40_ram[745] = 160;
    exp_40_ram[746] = 39;
    exp_40_ram[747] = 133;
    exp_40_ram[748] = 36;
    exp_40_ram[749] = 1;
    exp_40_ram[750] = 128;
    exp_40_ram[751] = 1;
    exp_40_ram[752] = 38;
    exp_40_ram[753] = 36;
    exp_40_ram[754] = 4;
    exp_40_ram[755] = 71;
    exp_40_ram[756] = 167;
    exp_40_ram[757] = 133;
    exp_40_ram[758] = 240;
    exp_40_ram[759] = 7;
    exp_40_ram[760] = 133;
    exp_40_ram[761] = 32;
    exp_40_ram[762] = 36;
    exp_40_ram[763] = 1;
    exp_40_ram[764] = 128;
    exp_40_ram[765] = 1;
    exp_40_ram[766] = 38;
    exp_40_ram[767] = 36;
    exp_40_ram[768] = 4;
    exp_40_ram[769] = 46;
    exp_40_ram[770] = 44;
    exp_40_ram[771] = 38;
    exp_40_ram[772] = 0;
    exp_40_ram[773] = 39;
    exp_40_ram[774] = 135;
    exp_40_ram[775] = 38;
    exp_40_ram[776] = 39;
    exp_40_ram[777] = 7;
    exp_40_ram[778] = 199;
    exp_40_ram[779] = 37;
    exp_40_ram[780] = 133;
    exp_40_ram[781] = 240;
    exp_40_ram[782] = 39;
    exp_40_ram[783] = 39;
    exp_40_ram[784] = 7;
    exp_40_ram[785] = 199;
    exp_40_ram[786] = 150;
    exp_40_ram[787] = 39;
    exp_40_ram[788] = 133;
    exp_40_ram[789] = 32;
    exp_40_ram[790] = 36;
    exp_40_ram[791] = 1;
    exp_40_ram[792] = 128;
    exp_40_ram[793] = 1;
    exp_40_ram[794] = 46;
    exp_40_ram[795] = 44;
    exp_40_ram[796] = 4;
    exp_40_ram[797] = 38;
    exp_40_ram[798] = 71;
    exp_40_ram[799] = 167;
    exp_40_ram[800] = 133;
    exp_40_ram[801] = 37;
    exp_40_ram[802] = 240;
    exp_40_ram[803] = 71;
    exp_40_ram[804] = 167;
    exp_40_ram[805] = 133;
    exp_40_ram[806] = 5;
    exp_40_ram[807] = 240;
    exp_40_ram[808] = 7;
    exp_40_ram[809] = 133;
    exp_40_ram[810] = 32;
    exp_40_ram[811] = 36;
    exp_40_ram[812] = 1;
    exp_40_ram[813] = 128;
    exp_40_ram[814] = 1;
    exp_40_ram[815] = 46;
    exp_40_ram[816] = 4;
    exp_40_ram[817] = 7;
    exp_40_ram[818] = 36;
    exp_40_ram[819] = 34;
    exp_40_ram[820] = 32;
    exp_40_ram[821] = 7;
    exp_40_ram[822] = 0;
    exp_40_ram[823] = 36;
    exp_40_ram[824] = 1;
    exp_40_ram[825] = 128;
    exp_40_ram[826] = 1;
    exp_40_ram[827] = 46;
    exp_40_ram[828] = 44;
    exp_40_ram[829] = 4;
    exp_40_ram[830] = 7;
    exp_40_ram[831] = 36;
    exp_40_ram[832] = 34;
    exp_40_ram[833] = 32;
    exp_40_ram[834] = 7;
    exp_40_ram[835] = 71;
    exp_40_ram[836] = 136;
    exp_40_ram[837] = 71;
    exp_40_ram[838] = 133;
    exp_40_ram[839] = 16;
    exp_40_ram[840] = 0;
    exp_40_ram[841] = 32;
    exp_40_ram[842] = 36;
    exp_40_ram[843] = 1;
    exp_40_ram[844] = 128;
    exp_40_ram[845] = 1;
    exp_40_ram[846] = 38;
    exp_40_ram[847] = 4;
    exp_40_ram[848] = 46;
    exp_40_ram[849] = 44;
    exp_40_ram[850] = 39;
    exp_40_ram[851] = 38;
    exp_40_ram[852] = 0;
    exp_40_ram[853] = 39;
    exp_40_ram[854] = 135;
    exp_40_ram[855] = 38;
    exp_40_ram[856] = 39;
    exp_40_ram[857] = 199;
    exp_40_ram[858] = 138;
    exp_40_ram[859] = 39;
    exp_40_ram[860] = 135;
    exp_40_ram[861] = 44;
    exp_40_ram[862] = 158;
    exp_40_ram[863] = 39;
    exp_40_ram[864] = 39;
    exp_40_ram[865] = 7;
    exp_40_ram[866] = 133;
    exp_40_ram[867] = 36;
    exp_40_ram[868] = 1;
    exp_40_ram[869] = 128;
    exp_40_ram[870] = 1;
    exp_40_ram[871] = 46;
    exp_40_ram[872] = 4;
    exp_40_ram[873] = 7;
    exp_40_ram[874] = 7;
    exp_40_ram[875] = 71;
    exp_40_ram[876] = 7;
    exp_40_ram[877] = 252;
    exp_40_ram[878] = 71;
    exp_40_ram[879] = 7;
    exp_40_ram[880] = 230;
    exp_40_ram[881] = 7;
    exp_40_ram[882] = 0;
    exp_40_ram[883] = 7;
    exp_40_ram[884] = 247;
    exp_40_ram[885] = 247;
    exp_40_ram[886] = 133;
    exp_40_ram[887] = 36;
    exp_40_ram[888] = 1;
    exp_40_ram[889] = 128;
    exp_40_ram[890] = 1;
    exp_40_ram[891] = 38;
    exp_40_ram[892] = 36;
    exp_40_ram[893] = 4;
    exp_40_ram[894] = 46;
    exp_40_ram[895] = 38;
    exp_40_ram[896] = 0;
    exp_40_ram[897] = 39;
    exp_40_ram[898] = 7;
    exp_40_ram[899] = 151;
    exp_40_ram[900] = 135;
    exp_40_ram[901] = 151;
    exp_40_ram[902] = 134;
    exp_40_ram[903] = 39;
    exp_40_ram[904] = 167;
    exp_40_ram[905] = 134;
    exp_40_ram[906] = 39;
    exp_40_ram[907] = 32;
    exp_40_ram[908] = 199;
    exp_40_ram[909] = 7;
    exp_40_ram[910] = 135;
    exp_40_ram[911] = 38;
    exp_40_ram[912] = 39;
    exp_40_ram[913] = 167;
    exp_40_ram[914] = 199;
    exp_40_ram[915] = 133;
    exp_40_ram[916] = 240;
    exp_40_ram[917] = 7;
    exp_40_ram[918] = 150;
    exp_40_ram[919] = 39;
    exp_40_ram[920] = 133;
    exp_40_ram[921] = 32;
    exp_40_ram[922] = 36;
    exp_40_ram[923] = 1;
    exp_40_ram[924] = 128;
    exp_40_ram[925] = 1;
    exp_40_ram[926] = 46;
    exp_40_ram[927] = 44;
    exp_40_ram[928] = 4;
    exp_40_ram[929] = 46;
    exp_40_ram[930] = 44;
    exp_40_ram[931] = 42;
    exp_40_ram[932] = 40;
    exp_40_ram[933] = 38;
    exp_40_ram[934] = 36;
    exp_40_ram[935] = 34;
    exp_40_ram[936] = 32;
    exp_40_ram[937] = 39;
    exp_40_ram[938] = 36;
    exp_40_ram[939] = 39;
    exp_40_ram[940] = 247;
    exp_40_ram[941] = 156;
    exp_40_ram[942] = 39;
    exp_40_ram[943] = 247;
    exp_40_ram[944] = 150;
    exp_40_ram[945] = 39;
    exp_40_ram[946] = 38;
    exp_40_ram[947] = 0;
    exp_40_ram[948] = 39;
    exp_40_ram[949] = 135;
    exp_40_ram[950] = 42;
    exp_40_ram[951] = 39;
    exp_40_ram[952] = 38;
    exp_40_ram[953] = 134;
    exp_40_ram[954] = 37;
    exp_40_ram[955] = 5;
    exp_40_ram[956] = 0;
    exp_40_ram[957] = 39;
    exp_40_ram[958] = 135;
    exp_40_ram[959] = 38;
    exp_40_ram[960] = 39;
    exp_40_ram[961] = 39;
    exp_40_ram[962] = 100;
    exp_40_ram[963] = 0;
    exp_40_ram[964] = 39;
    exp_40_ram[965] = 135;
    exp_40_ram[966] = 36;
    exp_40_ram[967] = 39;
    exp_40_ram[968] = 39;
    exp_40_ram[969] = 7;
    exp_40_ram[970] = 197;
    exp_40_ram[971] = 39;
    exp_40_ram[972] = 135;
    exp_40_ram[973] = 42;
    exp_40_ram[974] = 39;
    exp_40_ram[975] = 38;
    exp_40_ram[976] = 134;
    exp_40_ram[977] = 37;
    exp_40_ram[978] = 0;
    exp_40_ram[979] = 39;
    exp_40_ram[980] = 144;
    exp_40_ram[981] = 39;
    exp_40_ram[982] = 247;
    exp_40_ram[983] = 128;
    exp_40_ram[984] = 0;
    exp_40_ram[985] = 39;
    exp_40_ram[986] = 135;
    exp_40_ram[987] = 42;
    exp_40_ram[988] = 39;
    exp_40_ram[989] = 38;
    exp_40_ram[990] = 134;
    exp_40_ram[991] = 37;
    exp_40_ram[992] = 5;
    exp_40_ram[993] = 0;
    exp_40_ram[994] = 39;
    exp_40_ram[995] = 39;
    exp_40_ram[996] = 7;
    exp_40_ram[997] = 39;
    exp_40_ram[998] = 230;
    exp_40_ram[999] = 39;
    exp_40_ram[1000] = 133;
    exp_40_ram[1001] = 32;
    exp_40_ram[1002] = 36;
    exp_40_ram[1003] = 1;
    exp_40_ram[1004] = 128;
    exp_40_ram[1005] = 1;
    exp_40_ram[1006] = 38;
    exp_40_ram[1007] = 36;
    exp_40_ram[1008] = 4;
    exp_40_ram[1009] = 38;
    exp_40_ram[1010] = 36;
    exp_40_ram[1011] = 34;
    exp_40_ram[1012] = 32;
    exp_40_ram[1013] = 46;
    exp_40_ram[1014] = 44;
    exp_40_ram[1015] = 7;
    exp_40_ram[1016] = 40;
    exp_40_ram[1017] = 11;
    exp_40_ram[1018] = 39;
    exp_40_ram[1019] = 247;
    exp_40_ram[1020] = 154;
    exp_40_ram[1021] = 39;
    exp_40_ram[1022] = 136;
    exp_40_ram[1023] = 39;
    exp_40_ram[1024] = 247;
    exp_40_ram[1025] = 130;
    exp_40_ram[1026] = 71;
    exp_40_ram[1027] = 152;
    exp_40_ram[1028] = 39;
    exp_40_ram[1029] = 247;
    exp_40_ram[1030] = 136;
    exp_40_ram[1031] = 39;
    exp_40_ram[1032] = 135;
    exp_40_ram[1033] = 34;
    exp_40_ram[1034] = 0;
    exp_40_ram[1035] = 39;
    exp_40_ram[1036] = 135;
    exp_40_ram[1037] = 44;
    exp_40_ram[1038] = 39;
    exp_40_ram[1039] = 7;
    exp_40_ram[1040] = 7;
    exp_40_ram[1041] = 128;
    exp_40_ram[1042] = 39;
    exp_40_ram[1043] = 39;
    exp_40_ram[1044] = 120;
    exp_40_ram[1045] = 39;
    exp_40_ram[1046] = 7;
    exp_40_ram[1047] = 248;
    exp_40_ram[1048] = 0;
    exp_40_ram[1049] = 39;
    exp_40_ram[1050] = 135;
    exp_40_ram[1051] = 44;
    exp_40_ram[1052] = 39;
    exp_40_ram[1053] = 7;
    exp_40_ram[1054] = 7;
    exp_40_ram[1055] = 128;
    exp_40_ram[1056] = 39;
    exp_40_ram[1057] = 247;
    exp_40_ram[1058] = 142;
    exp_40_ram[1059] = 39;
    exp_40_ram[1060] = 39;
    exp_40_ram[1061] = 120;
    exp_40_ram[1062] = 39;
    exp_40_ram[1063] = 7;
    exp_40_ram[1064] = 242;
    exp_40_ram[1065] = 39;
    exp_40_ram[1066] = 247;
    exp_40_ram[1067] = 128;
    exp_40_ram[1068] = 39;
    exp_40_ram[1069] = 247;
    exp_40_ram[1070] = 152;
    exp_40_ram[1071] = 39;
    exp_40_ram[1072] = 132;
    exp_40_ram[1073] = 39;
    exp_40_ram[1074] = 39;
    exp_40_ram[1075] = 8;
    exp_40_ram[1076] = 39;
    exp_40_ram[1077] = 39;
    exp_40_ram[1078] = 24;
    exp_40_ram[1079] = 39;
    exp_40_ram[1080] = 135;
    exp_40_ram[1081] = 44;
    exp_40_ram[1082] = 39;
    exp_40_ram[1083] = 142;
    exp_40_ram[1084] = 39;
    exp_40_ram[1085] = 7;
    exp_40_ram[1086] = 24;
    exp_40_ram[1087] = 39;
    exp_40_ram[1088] = 135;
    exp_40_ram[1089] = 44;
    exp_40_ram[1090] = 39;
    exp_40_ram[1091] = 7;
    exp_40_ram[1092] = 30;
    exp_40_ram[1093] = 39;
    exp_40_ram[1094] = 247;
    exp_40_ram[1095] = 152;
    exp_40_ram[1096] = 39;
    exp_40_ram[1097] = 7;
    exp_40_ram[1098] = 226;
    exp_40_ram[1099] = 39;
    exp_40_ram[1100] = 135;
    exp_40_ram[1101] = 44;
    exp_40_ram[1102] = 39;
    exp_40_ram[1103] = 7;
    exp_40_ram[1104] = 7;
    exp_40_ram[1105] = 128;
    exp_40_ram[1106] = 0;
    exp_40_ram[1107] = 39;
    exp_40_ram[1108] = 7;
    exp_40_ram[1109] = 30;
    exp_40_ram[1110] = 39;
    exp_40_ram[1111] = 247;
    exp_40_ram[1112] = 136;
    exp_40_ram[1113] = 39;
    exp_40_ram[1114] = 7;
    exp_40_ram[1115] = 226;
    exp_40_ram[1116] = 39;
    exp_40_ram[1117] = 135;
    exp_40_ram[1118] = 44;
    exp_40_ram[1119] = 39;
    exp_40_ram[1120] = 7;
    exp_40_ram[1121] = 7;
    exp_40_ram[1122] = 128;
    exp_40_ram[1123] = 0;
    exp_40_ram[1124] = 39;
    exp_40_ram[1125] = 7;
    exp_40_ram[1126] = 22;
    exp_40_ram[1127] = 39;
    exp_40_ram[1128] = 7;
    exp_40_ram[1129] = 224;
    exp_40_ram[1130] = 39;
    exp_40_ram[1131] = 135;
    exp_40_ram[1132] = 44;
    exp_40_ram[1133] = 39;
    exp_40_ram[1134] = 7;
    exp_40_ram[1135] = 7;
    exp_40_ram[1136] = 128;
    exp_40_ram[1137] = 39;
    exp_40_ram[1138] = 7;
    exp_40_ram[1139] = 224;
    exp_40_ram[1140] = 39;
    exp_40_ram[1141] = 135;
    exp_40_ram[1142] = 44;
    exp_40_ram[1143] = 39;
    exp_40_ram[1144] = 7;
    exp_40_ram[1145] = 7;
    exp_40_ram[1146] = 128;
    exp_40_ram[1147] = 39;
    exp_40_ram[1148] = 7;
    exp_40_ram[1149] = 224;
    exp_40_ram[1150] = 71;
    exp_40_ram[1151] = 130;
    exp_40_ram[1152] = 39;
    exp_40_ram[1153] = 135;
    exp_40_ram[1154] = 44;
    exp_40_ram[1155] = 39;
    exp_40_ram[1156] = 7;
    exp_40_ram[1157] = 7;
    exp_40_ram[1158] = 128;
    exp_40_ram[1159] = 0;
    exp_40_ram[1160] = 39;
    exp_40_ram[1161] = 247;
    exp_40_ram[1162] = 130;
    exp_40_ram[1163] = 39;
    exp_40_ram[1164] = 135;
    exp_40_ram[1165] = 44;
    exp_40_ram[1166] = 39;
    exp_40_ram[1167] = 7;
    exp_40_ram[1168] = 7;
    exp_40_ram[1169] = 128;
    exp_40_ram[1170] = 0;
    exp_40_ram[1171] = 39;
    exp_40_ram[1172] = 247;
    exp_40_ram[1173] = 128;
    exp_40_ram[1174] = 39;
    exp_40_ram[1175] = 135;
    exp_40_ram[1176] = 44;
    exp_40_ram[1177] = 39;
    exp_40_ram[1178] = 7;
    exp_40_ram[1179] = 7;
    exp_40_ram[1180] = 128;
    exp_40_ram[1181] = 40;
    exp_40_ram[1182] = 40;
    exp_40_ram[1183] = 39;
    exp_40_ram[1184] = 39;
    exp_40_ram[1185] = 38;
    exp_40_ram[1186] = 38;
    exp_40_ram[1187] = 37;
    exp_40_ram[1188] = 37;
    exp_40_ram[1189] = 240;
    exp_40_ram[1190] = 7;
    exp_40_ram[1191] = 133;
    exp_40_ram[1192] = 32;
    exp_40_ram[1193] = 36;
    exp_40_ram[1194] = 1;
    exp_40_ram[1195] = 128;
    exp_40_ram[1196] = 1;
    exp_40_ram[1197] = 38;
    exp_40_ram[1198] = 36;
    exp_40_ram[1199] = 4;
    exp_40_ram[1200] = 46;
    exp_40_ram[1201] = 44;
    exp_40_ram[1202] = 42;
    exp_40_ram[1203] = 40;
    exp_40_ram[1204] = 38;
    exp_40_ram[1205] = 34;
    exp_40_ram[1206] = 32;
    exp_40_ram[1207] = 5;
    exp_40_ram[1208] = 38;
    exp_40_ram[1209] = 39;
    exp_40_ram[1210] = 152;
    exp_40_ram[1211] = 39;
    exp_40_ram[1212] = 247;
    exp_40_ram[1213] = 34;
    exp_40_ram[1214] = 39;
    exp_40_ram[1215] = 247;
    exp_40_ram[1216] = 134;
    exp_40_ram[1217] = 39;
    exp_40_ram[1218] = 140;
    exp_40_ram[1219] = 39;
    exp_40_ram[1220] = 39;
    exp_40_ram[1221] = 119;
    exp_40_ram[1222] = 5;
    exp_40_ram[1223] = 71;
    exp_40_ram[1224] = 7;
    exp_40_ram[1225] = 234;
    exp_40_ram[1226] = 71;
    exp_40_ram[1227] = 135;
    exp_40_ram[1228] = 247;
    exp_40_ram[1229] = 0;
    exp_40_ram[1230] = 39;
    exp_40_ram[1231] = 247;
    exp_40_ram[1232] = 134;
    exp_40_ram[1233] = 7;
    exp_40_ram[1234] = 0;
    exp_40_ram[1235] = 7;
    exp_40_ram[1236] = 71;
    exp_40_ram[1237] = 135;
    exp_40_ram[1238] = 247;
    exp_40_ram[1239] = 135;
    exp_40_ram[1240] = 247;
    exp_40_ram[1241] = 39;
    exp_40_ram[1242] = 6;
    exp_40_ram[1243] = 38;
    exp_40_ram[1244] = 6;
    exp_40_ram[1245] = 135;
    exp_40_ram[1246] = 12;
    exp_40_ram[1247] = 39;
    exp_40_ram[1248] = 39;
    exp_40_ram[1249] = 87;
    exp_40_ram[1250] = 38;
    exp_40_ram[1251] = 39;
    exp_40_ram[1252] = 136;
    exp_40_ram[1253] = 39;
    exp_40_ram[1254] = 7;
    exp_40_ram[1255] = 248;
    exp_40_ram[1256] = 70;
    exp_40_ram[1257] = 7;
    exp_40_ram[1258] = 39;
    exp_40_ram[1259] = 36;
    exp_40_ram[1260] = 39;
    exp_40_ram[1261] = 34;
    exp_40_ram[1262] = 39;
    exp_40_ram[1263] = 32;
    exp_40_ram[1264] = 40;
    exp_40_ram[1265] = 136;
    exp_40_ram[1266] = 39;
    exp_40_ram[1267] = 38;
    exp_40_ram[1268] = 38;
    exp_40_ram[1269] = 37;
    exp_40_ram[1270] = 37;
    exp_40_ram[1271] = 240;
    exp_40_ram[1272] = 7;
    exp_40_ram[1273] = 133;
    exp_40_ram[1274] = 32;
    exp_40_ram[1275] = 36;
    exp_40_ram[1276] = 1;
    exp_40_ram[1277] = 128;
    exp_40_ram[1278] = 1;
    exp_40_ram[1279] = 46;
    exp_40_ram[1280] = 44;
    exp_40_ram[1281] = 4;
    exp_40_ram[1282] = 38;
    exp_40_ram[1283] = 36;
    exp_40_ram[1284] = 34;
    exp_40_ram[1285] = 32;
    exp_40_ram[1286] = 46;
    exp_40_ram[1287] = 46;
    exp_40_ram[1288] = 39;
    exp_40_ram[1289] = 158;
    exp_40_ram[1290] = 23;
    exp_40_ram[1291] = 135;
    exp_40_ram[1292] = 38;
    exp_40_ram[1293] = 0;
    exp_40_ram[1294] = 39;
    exp_40_ram[1295] = 199;
    exp_40_ram[1296] = 7;
    exp_40_ram[1297] = 14;
    exp_40_ram[1298] = 39;
    exp_40_ram[1299] = 197;
    exp_40_ram[1300] = 39;
    exp_40_ram[1301] = 135;
    exp_40_ram[1302] = 46;
    exp_40_ram[1303] = 39;
    exp_40_ram[1304] = 38;
    exp_40_ram[1305] = 134;
    exp_40_ram[1306] = 37;
    exp_40_ram[1307] = 0;
    exp_40_ram[1308] = 39;
    exp_40_ram[1309] = 135;
    exp_40_ram[1310] = 32;
    exp_40_ram[1311] = 0;
    exp_40_ram[1312] = 39;
    exp_40_ram[1313] = 135;
    exp_40_ram[1314] = 32;
    exp_40_ram[1315] = 38;
    exp_40_ram[1316] = 39;
    exp_40_ram[1317] = 199;
    exp_40_ram[1318] = 135;
    exp_40_ram[1319] = 7;
    exp_40_ram[1320] = 104;
    exp_40_ram[1321] = 151;
    exp_40_ram[1322] = 71;
    exp_40_ram[1323] = 135;
    exp_40_ram[1324] = 7;
    exp_40_ram[1325] = 167;
    exp_40_ram[1326] = 128;
    exp_40_ram[1327] = 39;
    exp_40_ram[1328] = 231;
    exp_40_ram[1329] = 38;
    exp_40_ram[1330] = 39;
    exp_40_ram[1331] = 135;
    exp_40_ram[1332] = 32;
    exp_40_ram[1333] = 7;
    exp_40_ram[1334] = 32;
    exp_40_ram[1335] = 0;
    exp_40_ram[1336] = 39;
    exp_40_ram[1337] = 231;
    exp_40_ram[1338] = 38;
    exp_40_ram[1339] = 39;
    exp_40_ram[1340] = 135;
    exp_40_ram[1341] = 32;
    exp_40_ram[1342] = 7;
    exp_40_ram[1343] = 32;
    exp_40_ram[1344] = 0;
    exp_40_ram[1345] = 39;
    exp_40_ram[1346] = 231;
    exp_40_ram[1347] = 38;
    exp_40_ram[1348] = 39;
    exp_40_ram[1349] = 135;
    exp_40_ram[1350] = 32;
    exp_40_ram[1351] = 7;
    exp_40_ram[1352] = 32;
    exp_40_ram[1353] = 0;
    exp_40_ram[1354] = 39;
    exp_40_ram[1355] = 231;
    exp_40_ram[1356] = 38;
    exp_40_ram[1357] = 39;
    exp_40_ram[1358] = 135;
    exp_40_ram[1359] = 32;
    exp_40_ram[1360] = 7;
    exp_40_ram[1361] = 32;
    exp_40_ram[1362] = 0;
    exp_40_ram[1363] = 39;
    exp_40_ram[1364] = 231;
    exp_40_ram[1365] = 38;
    exp_40_ram[1366] = 39;
    exp_40_ram[1367] = 135;
    exp_40_ram[1368] = 32;
    exp_40_ram[1369] = 7;
    exp_40_ram[1370] = 32;
    exp_40_ram[1371] = 0;
    exp_40_ram[1372] = 32;
    exp_40_ram[1373] = 0;
    exp_40_ram[1374] = 39;
    exp_40_ram[1375] = 154;
    exp_40_ram[1376] = 36;
    exp_40_ram[1377] = 39;
    exp_40_ram[1378] = 199;
    exp_40_ram[1379] = 133;
    exp_40_ram[1380] = 240;
    exp_40_ram[1381] = 7;
    exp_40_ram[1382] = 140;
    exp_40_ram[1383] = 7;
    exp_40_ram[1384] = 133;
    exp_40_ram[1385] = 240;
    exp_40_ram[1386] = 36;
    exp_40_ram[1387] = 0;
    exp_40_ram[1388] = 39;
    exp_40_ram[1389] = 199;
    exp_40_ram[1390] = 7;
    exp_40_ram[1391] = 24;
    exp_40_ram[1392] = 39;
    exp_40_ram[1393] = 135;
    exp_40_ram[1394] = 46;
    exp_40_ram[1395] = 167;
    exp_40_ram[1396] = 36;
    exp_40_ram[1397] = 39;
    exp_40_ram[1398] = 208;
    exp_40_ram[1399] = 39;
    exp_40_ram[1400] = 231;
    exp_40_ram[1401] = 38;
    exp_40_ram[1402] = 39;
    exp_40_ram[1403] = 7;
    exp_40_ram[1404] = 36;
    exp_40_ram[1405] = 0;
    exp_40_ram[1406] = 39;
    exp_40_ram[1407] = 36;
    exp_40_ram[1408] = 39;
    exp_40_ram[1409] = 135;
    exp_40_ram[1410] = 32;
    exp_40_ram[1411] = 34;
    exp_40_ram[1412] = 39;
    exp_40_ram[1413] = 199;
    exp_40_ram[1414] = 7;
    exp_40_ram[1415] = 20;
    exp_40_ram[1416] = 39;
    exp_40_ram[1417] = 231;
    exp_40_ram[1418] = 38;
    exp_40_ram[1419] = 39;
    exp_40_ram[1420] = 135;
    exp_40_ram[1421] = 32;
    exp_40_ram[1422] = 39;
    exp_40_ram[1423] = 199;
    exp_40_ram[1424] = 133;
    exp_40_ram[1425] = 240;
    exp_40_ram[1426] = 7;
    exp_40_ram[1427] = 140;
    exp_40_ram[1428] = 7;
    exp_40_ram[1429] = 133;
    exp_40_ram[1430] = 240;
    exp_40_ram[1431] = 34;
    exp_40_ram[1432] = 0;
    exp_40_ram[1433] = 39;
    exp_40_ram[1434] = 199;
    exp_40_ram[1435] = 7;
    exp_40_ram[1436] = 26;
    exp_40_ram[1437] = 39;
    exp_40_ram[1438] = 135;
    exp_40_ram[1439] = 46;
    exp_40_ram[1440] = 167;
    exp_40_ram[1441] = 34;
    exp_40_ram[1442] = 39;
    exp_40_ram[1443] = 212;
    exp_40_ram[1444] = 7;
    exp_40_ram[1445] = 34;
    exp_40_ram[1446] = 39;
    exp_40_ram[1447] = 135;
    exp_40_ram[1448] = 32;
    exp_40_ram[1449] = 39;
    exp_40_ram[1450] = 199;
    exp_40_ram[1451] = 135;
    exp_40_ram[1452] = 7;
    exp_40_ram[1453] = 108;
    exp_40_ram[1454] = 151;
    exp_40_ram[1455] = 71;
    exp_40_ram[1456] = 135;
    exp_40_ram[1457] = 7;
    exp_40_ram[1458] = 167;
    exp_40_ram[1459] = 128;
    exp_40_ram[1460] = 39;
    exp_40_ram[1461] = 231;
    exp_40_ram[1462] = 38;
    exp_40_ram[1463] = 39;
    exp_40_ram[1464] = 135;
    exp_40_ram[1465] = 32;
    exp_40_ram[1466] = 39;
    exp_40_ram[1467] = 199;
    exp_40_ram[1468] = 7;
    exp_40_ram[1469] = 16;
    exp_40_ram[1470] = 39;
    exp_40_ram[1471] = 231;
    exp_40_ram[1472] = 38;
    exp_40_ram[1473] = 39;
    exp_40_ram[1474] = 135;
    exp_40_ram[1475] = 32;
    exp_40_ram[1476] = 0;
    exp_40_ram[1477] = 39;
    exp_40_ram[1478] = 231;
    exp_40_ram[1479] = 38;
    exp_40_ram[1480] = 39;
    exp_40_ram[1481] = 135;
    exp_40_ram[1482] = 32;
    exp_40_ram[1483] = 39;
    exp_40_ram[1484] = 199;
    exp_40_ram[1485] = 7;
    exp_40_ram[1486] = 18;
    exp_40_ram[1487] = 39;
    exp_40_ram[1488] = 231;
    exp_40_ram[1489] = 38;
    exp_40_ram[1490] = 39;
    exp_40_ram[1491] = 135;
    exp_40_ram[1492] = 32;
    exp_40_ram[1493] = 0;
    exp_40_ram[1494] = 39;
    exp_40_ram[1495] = 231;
    exp_40_ram[1496] = 38;
    exp_40_ram[1497] = 39;
    exp_40_ram[1498] = 135;
    exp_40_ram[1499] = 32;
    exp_40_ram[1500] = 0;
    exp_40_ram[1501] = 39;
    exp_40_ram[1502] = 231;
    exp_40_ram[1503] = 38;
    exp_40_ram[1504] = 39;
    exp_40_ram[1505] = 135;
    exp_40_ram[1506] = 32;
    exp_40_ram[1507] = 0;
    exp_40_ram[1508] = 39;
    exp_40_ram[1509] = 231;
    exp_40_ram[1510] = 38;
    exp_40_ram[1511] = 39;
    exp_40_ram[1512] = 135;
    exp_40_ram[1513] = 32;
    exp_40_ram[1514] = 0;
    exp_40_ram[1515] = 0;
    exp_40_ram[1516] = 0;
    exp_40_ram[1517] = 0;
    exp_40_ram[1518] = 0;
    exp_40_ram[1519] = 0;
    exp_40_ram[1520] = 39;
    exp_40_ram[1521] = 199;
    exp_40_ram[1522] = 135;
    exp_40_ram[1523] = 7;
    exp_40_ram[1524] = 108;
    exp_40_ram[1525] = 151;
    exp_40_ram[1526] = 71;
    exp_40_ram[1527] = 135;
    exp_40_ram[1528] = 7;
    exp_40_ram[1529] = 167;
    exp_40_ram[1530] = 128;
    exp_40_ram[1531] = 39;
    exp_40_ram[1532] = 199;
    exp_40_ram[1533] = 7;
    exp_40_ram[1534] = 10;
    exp_40_ram[1535] = 39;
    exp_40_ram[1536] = 199;
    exp_40_ram[1537] = 7;
    exp_40_ram[1538] = 24;
    exp_40_ram[1539] = 7;
    exp_40_ram[1540] = 44;
    exp_40_ram[1541] = 0;
    exp_40_ram[1542] = 39;
    exp_40_ram[1543] = 199;
    exp_40_ram[1544] = 7;
    exp_40_ram[1545] = 24;
    exp_40_ram[1546] = 7;
    exp_40_ram[1547] = 44;
    exp_40_ram[1548] = 0;
    exp_40_ram[1549] = 39;
    exp_40_ram[1550] = 199;
    exp_40_ram[1551] = 7;
    exp_40_ram[1552] = 24;
    exp_40_ram[1553] = 7;
    exp_40_ram[1554] = 44;
    exp_40_ram[1555] = 0;
    exp_40_ram[1556] = 7;
    exp_40_ram[1557] = 44;
    exp_40_ram[1558] = 39;
    exp_40_ram[1559] = 247;
    exp_40_ram[1560] = 38;
    exp_40_ram[1561] = 39;
    exp_40_ram[1562] = 199;
    exp_40_ram[1563] = 7;
    exp_40_ram[1564] = 24;
    exp_40_ram[1565] = 39;
    exp_40_ram[1566] = 231;
    exp_40_ram[1567] = 38;
    exp_40_ram[1568] = 39;
    exp_40_ram[1569] = 199;
    exp_40_ram[1570] = 7;
    exp_40_ram[1571] = 0;
    exp_40_ram[1572] = 39;
    exp_40_ram[1573] = 199;
    exp_40_ram[1574] = 7;
    exp_40_ram[1575] = 8;
    exp_40_ram[1576] = 39;
    exp_40_ram[1577] = 247;
    exp_40_ram[1578] = 38;
    exp_40_ram[1579] = 39;
    exp_40_ram[1580] = 247;
    exp_40_ram[1581] = 136;
    exp_40_ram[1582] = 39;
    exp_40_ram[1583] = 247;
    exp_40_ram[1584] = 38;
    exp_40_ram[1585] = 39;
    exp_40_ram[1586] = 199;
    exp_40_ram[1587] = 7;
    exp_40_ram[1588] = 10;
    exp_40_ram[1589] = 39;
    exp_40_ram[1590] = 199;
    exp_40_ram[1591] = 7;
    exp_40_ram[1592] = 24;
    exp_40_ram[1593] = 39;
    exp_40_ram[1594] = 247;
    exp_40_ram[1595] = 158;
    exp_40_ram[1596] = 39;
    exp_40_ram[1597] = 247;
    exp_40_ram[1598] = 140;
    exp_40_ram[1599] = 39;
    exp_40_ram[1600] = 135;
    exp_40_ram[1601] = 46;
    exp_40_ram[1602] = 167;
    exp_40_ram[1603] = 44;
    exp_40_ram[1604] = 39;
    exp_40_ram[1605] = 215;
    exp_40_ram[1606] = 39;
    exp_40_ram[1607] = 71;
    exp_40_ram[1608] = 135;
    exp_40_ram[1609] = 134;
    exp_40_ram[1610] = 39;
    exp_40_ram[1611] = 215;
    exp_40_ram[1612] = 247;
    exp_40_ram[1613] = 39;
    exp_40_ram[1614] = 34;
    exp_40_ram[1615] = 39;
    exp_40_ram[1616] = 32;
    exp_40_ram[1617] = 40;
    exp_40_ram[1618] = 40;
    exp_40_ram[1619] = 7;
    exp_40_ram[1620] = 135;
    exp_40_ram[1621] = 38;
    exp_40_ram[1622] = 38;
    exp_40_ram[1623] = 37;
    exp_40_ram[1624] = 37;
    exp_40_ram[1625] = 240;
    exp_40_ram[1626] = 46;
    exp_40_ram[1627] = 0;
    exp_40_ram[1628] = 39;
    exp_40_ram[1629] = 247;
    exp_40_ram[1630] = 142;
    exp_40_ram[1631] = 39;
    exp_40_ram[1632] = 135;
    exp_40_ram[1633] = 46;
    exp_40_ram[1634] = 167;
    exp_40_ram[1635] = 247;
    exp_40_ram[1636] = 0;
    exp_40_ram[1637] = 39;
    exp_40_ram[1638] = 247;
    exp_40_ram[1639] = 128;
    exp_40_ram[1640] = 39;
    exp_40_ram[1641] = 135;
    exp_40_ram[1642] = 46;
    exp_40_ram[1643] = 167;
    exp_40_ram[1644] = 151;
    exp_40_ram[1645] = 215;
    exp_40_ram[1646] = 0;
    exp_40_ram[1647] = 39;
    exp_40_ram[1648] = 135;
    exp_40_ram[1649] = 46;
    exp_40_ram[1650] = 167;
    exp_40_ram[1651] = 46;
    exp_40_ram[1652] = 39;
    exp_40_ram[1653] = 215;
    exp_40_ram[1654] = 39;
    exp_40_ram[1655] = 71;
    exp_40_ram[1656] = 135;
    exp_40_ram[1657] = 134;
    exp_40_ram[1658] = 39;
    exp_40_ram[1659] = 215;
    exp_40_ram[1660] = 247;
    exp_40_ram[1661] = 39;
    exp_40_ram[1662] = 34;
    exp_40_ram[1663] = 39;
    exp_40_ram[1664] = 32;
    exp_40_ram[1665] = 40;
    exp_40_ram[1666] = 40;
    exp_40_ram[1667] = 7;
    exp_40_ram[1668] = 135;
    exp_40_ram[1669] = 38;
    exp_40_ram[1670] = 38;
    exp_40_ram[1671] = 37;
    exp_40_ram[1672] = 37;
    exp_40_ram[1673] = 240;
    exp_40_ram[1674] = 46;
    exp_40_ram[1675] = 0;
    exp_40_ram[1676] = 39;
    exp_40_ram[1677] = 247;
    exp_40_ram[1678] = 152;
    exp_40_ram[1679] = 39;
    exp_40_ram[1680] = 247;
    exp_40_ram[1681] = 134;
    exp_40_ram[1682] = 39;
    exp_40_ram[1683] = 135;
    exp_40_ram[1684] = 46;
    exp_40_ram[1685] = 167;
    exp_40_ram[1686] = 39;
    exp_40_ram[1687] = 34;
    exp_40_ram[1688] = 39;
    exp_40_ram[1689] = 32;
    exp_40_ram[1690] = 40;
    exp_40_ram[1691] = 40;
    exp_40_ram[1692] = 7;
    exp_40_ram[1693] = 38;
    exp_40_ram[1694] = 38;
    exp_40_ram[1695] = 37;
    exp_40_ram[1696] = 37;
    exp_40_ram[1697] = 240;
    exp_40_ram[1698] = 46;
    exp_40_ram[1699] = 0;
    exp_40_ram[1700] = 39;
    exp_40_ram[1701] = 247;
    exp_40_ram[1702] = 142;
    exp_40_ram[1703] = 39;
    exp_40_ram[1704] = 135;
    exp_40_ram[1705] = 46;
    exp_40_ram[1706] = 167;
    exp_40_ram[1707] = 247;
    exp_40_ram[1708] = 0;
    exp_40_ram[1709] = 39;
    exp_40_ram[1710] = 247;
    exp_40_ram[1711] = 128;
    exp_40_ram[1712] = 39;
    exp_40_ram[1713] = 135;
    exp_40_ram[1714] = 46;
    exp_40_ram[1715] = 167;
    exp_40_ram[1716] = 151;
    exp_40_ram[1717] = 215;
    exp_40_ram[1718] = 0;
    exp_40_ram[1719] = 39;
    exp_40_ram[1720] = 135;
    exp_40_ram[1721] = 46;
    exp_40_ram[1722] = 167;
    exp_40_ram[1723] = 32;
    exp_40_ram[1724] = 39;
    exp_40_ram[1725] = 34;
    exp_40_ram[1726] = 39;
    exp_40_ram[1727] = 32;
    exp_40_ram[1728] = 40;
    exp_40_ram[1729] = 40;
    exp_40_ram[1730] = 7;
    exp_40_ram[1731] = 39;
    exp_40_ram[1732] = 38;
    exp_40_ram[1733] = 38;
    exp_40_ram[1734] = 37;
    exp_40_ram[1735] = 37;
    exp_40_ram[1736] = 240;
    exp_40_ram[1737] = 46;
    exp_40_ram[1738] = 39;
    exp_40_ram[1739] = 135;
    exp_40_ram[1740] = 32;
    exp_40_ram[1741] = 0;
    exp_40_ram[1742] = 7;
    exp_40_ram[1743] = 42;
    exp_40_ram[1744] = 39;
    exp_40_ram[1745] = 247;
    exp_40_ram[1746] = 144;
    exp_40_ram[1747] = 0;
    exp_40_ram[1748] = 39;
    exp_40_ram[1749] = 135;
    exp_40_ram[1750] = 46;
    exp_40_ram[1751] = 39;
    exp_40_ram[1752] = 38;
    exp_40_ram[1753] = 134;
    exp_40_ram[1754] = 37;
    exp_40_ram[1755] = 5;
    exp_40_ram[1756] = 0;
    exp_40_ram[1757] = 39;
    exp_40_ram[1758] = 135;
    exp_40_ram[1759] = 42;
    exp_40_ram[1760] = 39;
    exp_40_ram[1761] = 230;
    exp_40_ram[1762] = 39;
    exp_40_ram[1763] = 135;
    exp_40_ram[1764] = 46;
    exp_40_ram[1765] = 167;
    exp_40_ram[1766] = 245;
    exp_40_ram[1767] = 39;
    exp_40_ram[1768] = 135;
    exp_40_ram[1769] = 46;
    exp_40_ram[1770] = 39;
    exp_40_ram[1771] = 38;
    exp_40_ram[1772] = 134;
    exp_40_ram[1773] = 37;
    exp_40_ram[1774] = 0;
    exp_40_ram[1775] = 39;
    exp_40_ram[1776] = 247;
    exp_40_ram[1777] = 128;
    exp_40_ram[1778] = 0;
    exp_40_ram[1779] = 39;
    exp_40_ram[1780] = 135;
    exp_40_ram[1781] = 46;
    exp_40_ram[1782] = 39;
    exp_40_ram[1783] = 38;
    exp_40_ram[1784] = 134;
    exp_40_ram[1785] = 37;
    exp_40_ram[1786] = 5;
    exp_40_ram[1787] = 0;
    exp_40_ram[1788] = 39;
    exp_40_ram[1789] = 135;
    exp_40_ram[1790] = 42;
    exp_40_ram[1791] = 39;
    exp_40_ram[1792] = 230;
    exp_40_ram[1793] = 39;
    exp_40_ram[1794] = 135;
    exp_40_ram[1795] = 32;
    exp_40_ram[1796] = 0;
    exp_40_ram[1797] = 39;
    exp_40_ram[1798] = 135;
    exp_40_ram[1799] = 46;
    exp_40_ram[1800] = 167;
    exp_40_ram[1801] = 40;
    exp_40_ram[1802] = 39;
    exp_40_ram[1803] = 134;
    exp_40_ram[1804] = 39;
    exp_40_ram[1805] = 0;
    exp_40_ram[1806] = 7;
    exp_40_ram[1807] = 133;
    exp_40_ram[1808] = 37;
    exp_40_ram[1809] = 240;
    exp_40_ram[1810] = 38;
    exp_40_ram[1811] = 39;
    exp_40_ram[1812] = 247;
    exp_40_ram[1813] = 140;
    exp_40_ram[1814] = 39;
    exp_40_ram[1815] = 39;
    exp_40_ram[1816] = 116;
    exp_40_ram[1817] = 7;
    exp_40_ram[1818] = 38;
    exp_40_ram[1819] = 39;
    exp_40_ram[1820] = 247;
    exp_40_ram[1821] = 154;
    exp_40_ram[1822] = 0;
    exp_40_ram[1823] = 39;
    exp_40_ram[1824] = 135;
    exp_40_ram[1825] = 46;
    exp_40_ram[1826] = 39;
    exp_40_ram[1827] = 38;
    exp_40_ram[1828] = 134;
    exp_40_ram[1829] = 37;
    exp_40_ram[1830] = 5;
    exp_40_ram[1831] = 0;
    exp_40_ram[1832] = 39;
    exp_40_ram[1833] = 135;
    exp_40_ram[1834] = 38;
    exp_40_ram[1835] = 39;
    exp_40_ram[1836] = 230;
    exp_40_ram[1837] = 0;
    exp_40_ram[1838] = 39;
    exp_40_ram[1839] = 135;
    exp_40_ram[1840] = 40;
    exp_40_ram[1841] = 197;
    exp_40_ram[1842] = 39;
    exp_40_ram[1843] = 135;
    exp_40_ram[1844] = 46;
    exp_40_ram[1845] = 39;
    exp_40_ram[1846] = 38;
    exp_40_ram[1847] = 134;
    exp_40_ram[1848] = 37;
    exp_40_ram[1849] = 0;
    exp_40_ram[1850] = 39;
    exp_40_ram[1851] = 199;
    exp_40_ram[1852] = 128;
    exp_40_ram[1853] = 39;
    exp_40_ram[1854] = 247;
    exp_40_ram[1855] = 142;
    exp_40_ram[1856] = 39;
    exp_40_ram[1857] = 135;
    exp_40_ram[1858] = 34;
    exp_40_ram[1859] = 150;
    exp_40_ram[1860] = 39;
    exp_40_ram[1861] = 247;
    exp_40_ram[1862] = 128;
    exp_40_ram[1863] = 0;
    exp_40_ram[1864] = 39;
    exp_40_ram[1865] = 135;
    exp_40_ram[1866] = 46;
    exp_40_ram[1867] = 39;
    exp_40_ram[1868] = 38;
    exp_40_ram[1869] = 134;
    exp_40_ram[1870] = 37;
    exp_40_ram[1871] = 5;
    exp_40_ram[1872] = 0;
    exp_40_ram[1873] = 39;
    exp_40_ram[1874] = 135;
    exp_40_ram[1875] = 38;
    exp_40_ram[1876] = 39;
    exp_40_ram[1877] = 230;
    exp_40_ram[1878] = 39;
    exp_40_ram[1879] = 135;
    exp_40_ram[1880] = 32;
    exp_40_ram[1881] = 0;
    exp_40_ram[1882] = 7;
    exp_40_ram[1883] = 36;
    exp_40_ram[1884] = 39;
    exp_40_ram[1885] = 231;
    exp_40_ram[1886] = 38;
    exp_40_ram[1887] = 39;
    exp_40_ram[1888] = 135;
    exp_40_ram[1889] = 46;
    exp_40_ram[1890] = 167;
    exp_40_ram[1891] = 135;
    exp_40_ram[1892] = 39;
    exp_40_ram[1893] = 34;
    exp_40_ram[1894] = 39;
    exp_40_ram[1895] = 32;
    exp_40_ram[1896] = 40;
    exp_40_ram[1897] = 8;
    exp_40_ram[1898] = 7;
    exp_40_ram[1899] = 38;
    exp_40_ram[1900] = 38;
    exp_40_ram[1901] = 37;
    exp_40_ram[1902] = 37;
    exp_40_ram[1903] = 240;
    exp_40_ram[1904] = 46;
    exp_40_ram[1905] = 39;
    exp_40_ram[1906] = 135;
    exp_40_ram[1907] = 32;
    exp_40_ram[1908] = 0;
    exp_40_ram[1909] = 39;
    exp_40_ram[1910] = 135;
    exp_40_ram[1911] = 46;
    exp_40_ram[1912] = 39;
    exp_40_ram[1913] = 38;
    exp_40_ram[1914] = 134;
    exp_40_ram[1915] = 37;
    exp_40_ram[1916] = 5;
    exp_40_ram[1917] = 0;
    exp_40_ram[1918] = 39;
    exp_40_ram[1919] = 135;
    exp_40_ram[1920] = 32;
    exp_40_ram[1921] = 0;
    exp_40_ram[1922] = 39;
    exp_40_ram[1923] = 197;
    exp_40_ram[1924] = 39;
    exp_40_ram[1925] = 135;
    exp_40_ram[1926] = 46;
    exp_40_ram[1927] = 39;
    exp_40_ram[1928] = 38;
    exp_40_ram[1929] = 134;
    exp_40_ram[1930] = 37;
    exp_40_ram[1931] = 0;
    exp_40_ram[1932] = 39;
    exp_40_ram[1933] = 135;
    exp_40_ram[1934] = 32;
    exp_40_ram[1935] = 0;
    exp_40_ram[1936] = 39;
    exp_40_ram[1937] = 199;
    exp_40_ram[1938] = 152;
    exp_40_ram[1939] = 39;
    exp_40_ram[1940] = 39;
    exp_40_ram[1941] = 104;
    exp_40_ram[1942] = 39;
    exp_40_ram[1943] = 135;
    exp_40_ram[1944] = 0;
    exp_40_ram[1945] = 39;
    exp_40_ram[1946] = 39;
    exp_40_ram[1947] = 38;
    exp_40_ram[1948] = 134;
    exp_40_ram[1949] = 37;
    exp_40_ram[1950] = 5;
    exp_40_ram[1951] = 0;
    exp_40_ram[1952] = 39;
    exp_40_ram[1953] = 133;
    exp_40_ram[1954] = 32;
    exp_40_ram[1955] = 36;
    exp_40_ram[1956] = 1;
    exp_40_ram[1957] = 128;
    exp_40_ram[1958] = 1;
    exp_40_ram[1959] = 38;
    exp_40_ram[1960] = 36;
    exp_40_ram[1961] = 4;
    exp_40_ram[1962] = 46;
    exp_40_ram[1963] = 34;
    exp_40_ram[1964] = 36;
    exp_40_ram[1965] = 38;
    exp_40_ram[1966] = 40;
    exp_40_ram[1967] = 42;
    exp_40_ram[1968] = 44;
    exp_40_ram[1969] = 46;
    exp_40_ram[1970] = 7;
    exp_40_ram[1971] = 44;
    exp_40_ram[1972] = 39;
    exp_40_ram[1973] = 135;
    exp_40_ram[1974] = 36;
    exp_40_ram[1975] = 39;
    exp_40_ram[1976] = 7;
    exp_40_ram[1977] = 38;
    exp_40_ram[1978] = 6;
    exp_40_ram[1979] = 133;
    exp_40_ram[1980] = 23;
    exp_40_ram[1981] = 133;
    exp_40_ram[1982] = 240;
    exp_40_ram[1983] = 38;
    exp_40_ram[1984] = 39;
    exp_40_ram[1985] = 133;
    exp_40_ram[1986] = 32;
    exp_40_ram[1987] = 36;
    exp_40_ram[1988] = 1;
    exp_40_ram[1989] = 128;
    exp_40_ram[1990] = 1;
    exp_40_ram[1991] = 46;
    exp_40_ram[1992] = 44;
    exp_40_ram[1993] = 4;
    exp_40_ram[1994] = 7;
    exp_40_ram[1995] = 7;
    exp_40_ram[1996] = 71;
    exp_40_ram[1997] = 71;
    exp_40_ram[1998] = 167;
    exp_40_ram[1999] = 133;
    exp_40_ram[2000] = 5;
    exp_40_ram[2001] = 224;
    exp_40_ram[2002] = 0;
    exp_40_ram[2003] = 32;
    exp_40_ram[2004] = 36;
    exp_40_ram[2005] = 1;
    exp_40_ram[2006] = 128;
    exp_40_ram[2007] = 1;
    exp_40_ram[2008] = 46;
    exp_40_ram[2009] = 44;
    exp_40_ram[2010] = 42;
    exp_40_ram[2011] = 4;
    exp_40_ram[2012] = 4;
    exp_40_ram[2013] = 167;
    exp_40_ram[2014] = 36;
    exp_40_ram[2015] = 7;
    exp_40_ram[2016] = 34;
    exp_40_ram[2017] = 7;
    exp_40_ram[2018] = 32;
    exp_40_ram[2019] = 7;
    exp_40_ram[2020] = 46;
    exp_40_ram[2021] = 44;
    exp_40_ram[2022] = 42;
    exp_40_ram[2023] = 42;
    exp_40_ram[2024] = 35;
    exp_40_ram[2025] = 40;
    exp_40_ram[2026] = 40;
    exp_40_ram[2027] = 37;
    exp_40_ram[2028] = 37;
    exp_40_ram[2029] = 38;
    exp_40_ram[2030] = 38;
    exp_40_ram[2031] = 39;
    exp_40_ram[2032] = 39;
    exp_40_ram[2033] = 32;
    exp_40_ram[2034] = 34;
    exp_40_ram[2035] = 36;
    exp_40_ram[2036] = 38;
    exp_40_ram[2037] = 40;
    exp_40_ram[2038] = 42;
    exp_40_ram[2039] = 44;
    exp_40_ram[2040] = 46;
    exp_40_ram[2041] = 32;
    exp_40_ram[2042] = 7;
    exp_40_ram[2043] = 133;
    exp_40_ram[2044] = 0;
    exp_40_ram[2045] = 36;
    exp_40_ram[2046] = 38;
    exp_40_ram[2047] = 7;
    exp_40_ram[2048] = 37;
    exp_40_ram[2049] = 38;
    exp_40_ram[2050] = 133;
    exp_40_ram[2051] = 16;
    exp_40_ram[2052] = 39;
    exp_40_ram[2053] = 39;
    exp_40_ram[2054] = 7;
    exp_40_ram[2055] = 32;
    exp_40_ram[2056] = 35;
    exp_40_ram[2057] = 40;
    exp_40_ram[2058] = 40;
    exp_40_ram[2059] = 37;
    exp_40_ram[2060] = 37;
    exp_40_ram[2061] = 38;
    exp_40_ram[2062] = 38;
    exp_40_ram[2063] = 39;
    exp_40_ram[2064] = 39;
    exp_40_ram[2065] = 32;
    exp_40_ram[2066] = 34;
    exp_40_ram[2067] = 36;
    exp_40_ram[2068] = 38;
    exp_40_ram[2069] = 40;
    exp_40_ram[2070] = 42;
    exp_40_ram[2071] = 44;
    exp_40_ram[2072] = 46;
    exp_40_ram[2073] = 32;
    exp_40_ram[2074] = 7;
    exp_40_ram[2075] = 133;
    exp_40_ram[2076] = 0;
    exp_40_ram[2077] = 36;
    exp_40_ram[2078] = 38;
    exp_40_ram[2079] = 167;
    exp_40_ram[2080] = 34;
    exp_40_ram[2081] = 7;
    exp_40_ram[2082] = 32;
    exp_40_ram[2083] = 7;
    exp_40_ram[2084] = 46;
    exp_40_ram[2085] = 7;
    exp_40_ram[2086] = 44;
    exp_40_ram[2087] = 42;
    exp_40_ram[2088] = 40;
    exp_40_ram[2089] = 42;
    exp_40_ram[2090] = 35;
    exp_40_ram[2091] = 40;
    exp_40_ram[2092] = 40;
    exp_40_ram[2093] = 37;
    exp_40_ram[2094] = 37;
    exp_40_ram[2095] = 38;
    exp_40_ram[2096] = 38;
    exp_40_ram[2097] = 39;
    exp_40_ram[2098] = 39;
    exp_40_ram[2099] = 32;
    exp_40_ram[2100] = 34;
    exp_40_ram[2101] = 36;
    exp_40_ram[2102] = 38;
    exp_40_ram[2103] = 40;
    exp_40_ram[2104] = 42;
    exp_40_ram[2105] = 44;
    exp_40_ram[2106] = 46;
    exp_40_ram[2107] = 32;
    exp_40_ram[2108] = 7;
    exp_40_ram[2109] = 133;
    exp_40_ram[2110] = 0;
    exp_40_ram[2111] = 32;
    exp_40_ram[2112] = 34;
    exp_40_ram[2113] = 7;
    exp_40_ram[2114] = 37;
    exp_40_ram[2115] = 38;
    exp_40_ram[2116] = 133;
    exp_40_ram[2117] = 0;
    exp_40_ram[2118] = 39;
    exp_40_ram[2119] = 39;
    exp_40_ram[2120] = 7;
    exp_40_ram[2121] = 46;
    exp_40_ram[2122] = 35;
    exp_40_ram[2123] = 40;
    exp_40_ram[2124] = 40;
    exp_40_ram[2125] = 37;
    exp_40_ram[2126] = 37;
    exp_40_ram[2127] = 38;
    exp_40_ram[2128] = 38;
    exp_40_ram[2129] = 39;
    exp_40_ram[2130] = 39;
    exp_40_ram[2131] = 32;
    exp_40_ram[2132] = 34;
    exp_40_ram[2133] = 36;
    exp_40_ram[2134] = 38;
    exp_40_ram[2135] = 40;
    exp_40_ram[2136] = 42;
    exp_40_ram[2137] = 44;
    exp_40_ram[2138] = 46;
    exp_40_ram[2139] = 32;
    exp_40_ram[2140] = 7;
    exp_40_ram[2141] = 133;
    exp_40_ram[2142] = 0;
    exp_40_ram[2143] = 32;
    exp_40_ram[2144] = 34;
    exp_40_ram[2145] = 163;
    exp_40_ram[2146] = 168;
    exp_40_ram[2147] = 168;
    exp_40_ram[2148] = 165;
    exp_40_ram[2149] = 165;
    exp_40_ram[2150] = 166;
    exp_40_ram[2151] = 166;
    exp_40_ram[2152] = 167;
    exp_40_ram[2153] = 167;
    exp_40_ram[2154] = 32;
    exp_40_ram[2155] = 34;
    exp_40_ram[2156] = 36;
    exp_40_ram[2157] = 38;
    exp_40_ram[2158] = 40;
    exp_40_ram[2159] = 42;
    exp_40_ram[2160] = 44;
    exp_40_ram[2161] = 46;
    exp_40_ram[2162] = 32;
    exp_40_ram[2163] = 7;
    exp_40_ram[2164] = 133;
    exp_40_ram[2165] = 0;
    exp_40_ram[2166] = 44;
    exp_40_ram[2167] = 46;
    exp_40_ram[2168] = 39;
    exp_40_ram[2169] = 39;
    exp_40_ram[2170] = 228;
    exp_40_ram[2171] = 39;
    exp_40_ram[2172] = 39;
    exp_40_ram[2173] = 24;
    exp_40_ram[2174] = 39;
    exp_40_ram[2175] = 39;
    exp_40_ram[2176] = 232;
    exp_40_ram[2177] = 39;
    exp_40_ram[2178] = 39;
    exp_40_ram[2179] = 238;
    exp_40_ram[2180] = 39;
    exp_40_ram[2181] = 39;
    exp_40_ram[2182] = 28;
    exp_40_ram[2183] = 39;
    exp_40_ram[2184] = 39;
    exp_40_ram[2185] = 246;
    exp_40_ram[2186] = 7;
    exp_40_ram[2187] = 0;
    exp_40_ram[2188] = 7;
    exp_40_ram[2189] = 133;
    exp_40_ram[2190] = 32;
    exp_40_ram[2191] = 36;
    exp_40_ram[2192] = 36;
    exp_40_ram[2193] = 1;
    exp_40_ram[2194] = 128;
    exp_40_ram[2195] = 1;
    exp_40_ram[2196] = 46;
    exp_40_ram[2197] = 44;
    exp_40_ram[2198] = 4;
    exp_40_ram[2199] = 44;
    exp_40_ram[2200] = 46;
    exp_40_ram[2201] = 7;
    exp_40_ram[2202] = 37;
    exp_40_ram[2203] = 38;
    exp_40_ram[2204] = 133;
    exp_40_ram[2205] = 0;
    exp_40_ram[2206] = 35;
    exp_40_ram[2207] = 40;
    exp_40_ram[2208] = 40;
    exp_40_ram[2209] = 37;
    exp_40_ram[2210] = 37;
    exp_40_ram[2211] = 38;
    exp_40_ram[2212] = 38;
    exp_40_ram[2213] = 39;
    exp_40_ram[2214] = 39;
    exp_40_ram[2215] = 32;
    exp_40_ram[2216] = 34;
    exp_40_ram[2217] = 36;
    exp_40_ram[2218] = 38;
    exp_40_ram[2219] = 40;
    exp_40_ram[2220] = 42;
    exp_40_ram[2221] = 44;
    exp_40_ram[2222] = 46;
    exp_40_ram[2223] = 32;
    exp_40_ram[2224] = 7;
    exp_40_ram[2225] = 133;
    exp_40_ram[2226] = 240;
    exp_40_ram[2227] = 7;
    exp_40_ram[2228] = 133;
    exp_40_ram[2229] = 32;
    exp_40_ram[2230] = 36;
    exp_40_ram[2231] = 1;
    exp_40_ram[2232] = 128;
    exp_40_ram[2233] = 1;
    exp_40_ram[2234] = 46;
    exp_40_ram[2235] = 4;
    exp_40_ram[2236] = 6;
    exp_40_ram[2237] = 38;
    exp_40_ram[2238] = 6;
    exp_40_ram[2239] = 134;
    exp_40_ram[2240] = 36;
    exp_40_ram[2241] = 38;
    exp_40_ram[2242] = 166;
    exp_40_ram[2243] = 166;
    exp_40_ram[2244] = 40;
    exp_40_ram[2245] = 40;
    exp_40_ram[2246] = 40;
    exp_40_ram[2247] = 23;
    exp_40_ram[2248] = 7;
    exp_40_ram[2249] = 101;
    exp_40_ram[2250] = 229;
    exp_40_ram[2251] = 7;
    exp_40_ram[2252] = 135;
    exp_40_ram[2253] = 5;
    exp_40_ram[2254] = 133;
    exp_40_ram[2255] = 36;
    exp_40_ram[2256] = 1;
    exp_40_ram[2257] = 128;
    exp_40_ram[2258] = 1;
    exp_40_ram[2259] = 46;
    exp_40_ram[2260] = 44;
    exp_40_ram[2261] = 4;
    exp_40_ram[2262] = 36;
    exp_40_ram[2263] = 38;
    exp_40_ram[2264] = 32;
    exp_40_ram[2265] = 34;
    exp_40_ram[2266] = 39;
    exp_40_ram[2267] = 39;
    exp_40_ram[2268] = 37;
    exp_40_ram[2269] = 37;
    exp_40_ram[2270] = 6;
    exp_40_ram[2271] = 8;
    exp_40_ram[2272] = 56;
    exp_40_ram[2273] = 134;
    exp_40_ram[2274] = 135;
    exp_40_ram[2275] = 134;
    exp_40_ram[2276] = 7;
    exp_40_ram[2277] = 135;
    exp_40_ram[2278] = 5;
    exp_40_ram[2279] = 133;
    exp_40_ram[2280] = 224;
    exp_40_ram[2281] = 7;
    exp_40_ram[2282] = 135;
    exp_40_ram[2283] = 5;
    exp_40_ram[2284] = 133;
    exp_40_ram[2285] = 32;
    exp_40_ram[2286] = 36;
    exp_40_ram[2287] = 1;
    exp_40_ram[2288] = 128;
    exp_40_ram[2289] = 1;
    exp_40_ram[2290] = 46;
    exp_40_ram[2291] = 4;
    exp_40_ram[2292] = 38;
    exp_40_ram[2293] = 39;
    exp_40_ram[2294] = 247;
    exp_40_ram[2295] = 150;
    exp_40_ram[2296] = 39;
    exp_40_ram[2297] = 7;
    exp_40_ram[2298] = 119;
    exp_40_ram[2299] = 154;
    exp_40_ram[2300] = 39;
    exp_40_ram[2301] = 7;
    exp_40_ram[2302] = 119;
    exp_40_ram[2303] = 150;
    exp_40_ram[2304] = 7;
    exp_40_ram[2305] = 0;
    exp_40_ram[2306] = 7;
    exp_40_ram[2307] = 133;
    exp_40_ram[2308] = 36;
    exp_40_ram[2309] = 1;
    exp_40_ram[2310] = 128;
    exp_40_ram[2311] = 1;
    exp_40_ram[2312] = 46;
    exp_40_ram[2313] = 44;
    exp_40_ram[2314] = 4;
    exp_40_ram[2315] = 38;
    exp_40_ram[2316] = 37;
    exp_40_ram[2317] = 240;
    exp_40_ram[2318] = 7;
    exp_40_ram[2319] = 134;
    exp_40_ram[2320] = 7;
    exp_40_ram[2321] = 0;
    exp_40_ram[2322] = 7;
    exp_40_ram[2323] = 133;
    exp_40_ram[2324] = 32;
    exp_40_ram[2325] = 36;
    exp_40_ram[2326] = 1;
    exp_40_ram[2327] = 128;
    exp_40_ram[2328] = 1;
    exp_40_ram[2329] = 46;
    exp_40_ram[2330] = 44;
    exp_40_ram[2331] = 4;
    exp_40_ram[2332] = 38;
    exp_40_ram[2333] = 36;
    exp_40_ram[2334] = 39;
    exp_40_ram[2335] = 7;
    exp_40_ram[2336] = 4;
    exp_40_ram[2337] = 39;
    exp_40_ram[2338] = 7;
    exp_40_ram[2339] = 14;
    exp_40_ram[2340] = 39;
    exp_40_ram[2341] = 7;
    exp_40_ram[2342] = 8;
    exp_40_ram[2343] = 39;
    exp_40_ram[2344] = 7;
    exp_40_ram[2345] = 22;
    exp_40_ram[2346] = 7;
    exp_40_ram[2347] = 0;
    exp_40_ram[2348] = 39;
    exp_40_ram[2349] = 7;
    exp_40_ram[2350] = 18;
    exp_40_ram[2351] = 37;
    exp_40_ram[2352] = 240;
    exp_40_ram[2353] = 7;
    exp_40_ram[2354] = 134;
    exp_40_ram[2355] = 7;
    exp_40_ram[2356] = 0;
    exp_40_ram[2357] = 7;
    exp_40_ram[2358] = 0;
    exp_40_ram[2359] = 7;
    exp_40_ram[2360] = 133;
    exp_40_ram[2361] = 32;
    exp_40_ram[2362] = 36;
    exp_40_ram[2363] = 1;
    exp_40_ram[2364] = 128;
    exp_40_ram[2365] = 1;
    exp_40_ram[2366] = 38;
    exp_40_ram[2367] = 36;
    exp_40_ram[2368] = 34;
    exp_40_ram[2369] = 32;
    exp_40_ram[2370] = 46;
    exp_40_ram[2371] = 44;
    exp_40_ram[2372] = 42;
    exp_40_ram[2373] = 40;
    exp_40_ram[2374] = 38;
    exp_40_ram[2375] = 36;
    exp_40_ram[2376] = 34;
    exp_40_ram[2377] = 32;
    exp_40_ram[2378] = 46;
    exp_40_ram[2379] = 4;
    exp_40_ram[2380] = 4;
    exp_40_ram[2381] = 7;
    exp_40_ram[2382] = 8;
    exp_40_ram[2383] = 44;
    exp_40_ram[2384] = 46;
    exp_40_ram[2385] = 7;
    exp_40_ram[2386] = 42;
    exp_40_ram[2387] = 167;
    exp_40_ram[2388] = 38;
    exp_40_ram[2389] = 39;
    exp_40_ram[2390] = 135;
    exp_40_ram[2391] = 39;
    exp_40_ram[2392] = 6;
    exp_40_ram[2393] = 37;
    exp_40_ram[2394] = 240;
    exp_40_ram[2395] = 7;
    exp_40_ram[2396] = 87;
    exp_40_ram[2397] = 135;
    exp_40_ram[2398] = 7;
    exp_40_ram[2399] = 44;
    exp_40_ram[2400] = 46;
    exp_40_ram[2401] = 38;
    exp_40_ram[2402] = 38;
    exp_40_ram[2403] = 40;
    exp_40_ram[2404] = 40;
    exp_40_ram[2405] = 5;
    exp_40_ram[2406] = 7;
    exp_40_ram[2407] = 5;
    exp_40_ram[2408] = 181;
    exp_40_ram[2409] = 133;
    exp_40_ram[2410] = 135;
    exp_40_ram[2411] = 134;
    exp_40_ram[2412] = 135;
    exp_40_ram[2413] = 44;
    exp_40_ram[2414] = 46;
    exp_40_ram[2415] = 39;
    exp_40_ram[2416] = 135;
    exp_40_ram[2417] = 42;
    exp_40_ram[2418] = 240;
    exp_40_ram[2419] = 0;
    exp_40_ram[2420] = 40;
    exp_40_ram[2421] = 167;
    exp_40_ram[2422] = 135;
    exp_40_ram[2423] = 39;
    exp_40_ram[2424] = 128;
    exp_40_ram[2425] = 37;
    exp_40_ram[2426] = 37;
    exp_40_ram[2427] = 240;
    exp_40_ram[2428] = 7;
    exp_40_ram[2429] = 87;
    exp_40_ram[2430] = 135;
    exp_40_ram[2431] = 7;
    exp_40_ram[2432] = 141;
    exp_40_ram[2433] = 13;
    exp_40_ram[2434] = 38;
    exp_40_ram[2435] = 38;
    exp_40_ram[2436] = 7;
    exp_40_ram[2437] = 5;
    exp_40_ram[2438] = 181;
    exp_40_ram[2439] = 135;
    exp_40_ram[2440] = 134;
    exp_40_ram[2441] = 135;
    exp_40_ram[2442] = 44;
    exp_40_ram[2443] = 46;
    exp_40_ram[2444] = 39;
    exp_40_ram[2445] = 135;
    exp_40_ram[2446] = 40;
    exp_40_ram[2447] = 240;
    exp_40_ram[2448] = 0;
    exp_40_ram[2449] = 167;
    exp_40_ram[2450] = 135;
    exp_40_ram[2451] = 87;
    exp_40_ram[2452] = 135;
    exp_40_ram[2453] = 7;
    exp_40_ram[2454] = 140;
    exp_40_ram[2455] = 215;
    exp_40_ram[2456] = 140;
    exp_40_ram[2457] = 38;
    exp_40_ram[2458] = 38;
    exp_40_ram[2459] = 7;
    exp_40_ram[2460] = 5;
    exp_40_ram[2461] = 181;
    exp_40_ram[2462] = 135;
    exp_40_ram[2463] = 134;
    exp_40_ram[2464] = 135;
    exp_40_ram[2465] = 44;
    exp_40_ram[2466] = 46;
    exp_40_ram[2467] = 167;
    exp_40_ram[2468] = 23;
    exp_40_ram[2469] = 135;
    exp_40_ram[2470] = 7;
    exp_40_ram[2471] = 139;
    exp_40_ram[2472] = 215;
    exp_40_ram[2473] = 139;
    exp_40_ram[2474] = 38;
    exp_40_ram[2475] = 38;
    exp_40_ram[2476] = 7;
    exp_40_ram[2477] = 5;
    exp_40_ram[2478] = 181;
    exp_40_ram[2479] = 135;
    exp_40_ram[2480] = 134;
    exp_40_ram[2481] = 135;
    exp_40_ram[2482] = 44;
    exp_40_ram[2483] = 46;
    exp_40_ram[2484] = 167;
    exp_40_ram[2485] = 7;
    exp_40_ram[2486] = 151;
    exp_40_ram[2487] = 135;
    exp_40_ram[2488] = 151;
    exp_40_ram[2489] = 138;
    exp_40_ram[2490] = 215;
    exp_40_ram[2491] = 138;
    exp_40_ram[2492] = 38;
    exp_40_ram[2493] = 38;
    exp_40_ram[2494] = 7;
    exp_40_ram[2495] = 5;
    exp_40_ram[2496] = 181;
    exp_40_ram[2497] = 135;
    exp_40_ram[2498] = 134;
    exp_40_ram[2499] = 135;
    exp_40_ram[2500] = 44;
    exp_40_ram[2501] = 46;
    exp_40_ram[2502] = 167;
    exp_40_ram[2503] = 137;
    exp_40_ram[2504] = 215;
    exp_40_ram[2505] = 137;
    exp_40_ram[2506] = 38;
    exp_40_ram[2507] = 38;
    exp_40_ram[2508] = 7;
    exp_40_ram[2509] = 5;
    exp_40_ram[2510] = 181;
    exp_40_ram[2511] = 135;
    exp_40_ram[2512] = 134;
    exp_40_ram[2513] = 135;
    exp_40_ram[2514] = 44;
    exp_40_ram[2515] = 46;
    exp_40_ram[2516] = 39;
    exp_40_ram[2517] = 39;
    exp_40_ram[2518] = 5;
    exp_40_ram[2519] = 133;
    exp_40_ram[2520] = 32;
    exp_40_ram[2521] = 36;
    exp_40_ram[2522] = 36;
    exp_40_ram[2523] = 41;
    exp_40_ram[2524] = 41;
    exp_40_ram[2525] = 42;
    exp_40_ram[2526] = 42;
    exp_40_ram[2527] = 43;
    exp_40_ram[2528] = 43;
    exp_40_ram[2529] = 44;
    exp_40_ram[2530] = 44;
    exp_40_ram[2531] = 45;
    exp_40_ram[2532] = 45;
    exp_40_ram[2533] = 1;
    exp_40_ram[2534] = 128;
    exp_40_ram[2535] = 1;
    exp_40_ram[2536] = 46;
    exp_40_ram[2537] = 44;
    exp_40_ram[2538] = 42;
    exp_40_ram[2539] = 40;
    exp_40_ram[2540] = 38;
    exp_40_ram[2541] = 4;
    exp_40_ram[2542] = 46;
    exp_40_ram[2543] = 39;
    exp_40_ram[2544] = 163;
    exp_40_ram[2545] = 168;
    exp_40_ram[2546] = 168;
    exp_40_ram[2547] = 165;
    exp_40_ram[2548] = 165;
    exp_40_ram[2549] = 166;
    exp_40_ram[2550] = 166;
    exp_40_ram[2551] = 167;
    exp_40_ram[2552] = 167;
    exp_40_ram[2553] = 38;
    exp_40_ram[2554] = 40;
    exp_40_ram[2555] = 42;
    exp_40_ram[2556] = 44;
    exp_40_ram[2557] = 46;
    exp_40_ram[2558] = 32;
    exp_40_ram[2559] = 34;
    exp_40_ram[2560] = 36;
    exp_40_ram[2561] = 38;
    exp_40_ram[2562] = 35;
    exp_40_ram[2563] = 40;
    exp_40_ram[2564] = 40;
    exp_40_ram[2565] = 37;
    exp_40_ram[2566] = 37;
    exp_40_ram[2567] = 38;
    exp_40_ram[2568] = 38;
    exp_40_ram[2569] = 39;
    exp_40_ram[2570] = 39;
    exp_40_ram[2571] = 32;
    exp_40_ram[2572] = 34;
    exp_40_ram[2573] = 36;
    exp_40_ram[2574] = 38;
    exp_40_ram[2575] = 40;
    exp_40_ram[2576] = 42;
    exp_40_ram[2577] = 44;
    exp_40_ram[2578] = 46;
    exp_40_ram[2579] = 32;
    exp_40_ram[2580] = 7;
    exp_40_ram[2581] = 133;
    exp_40_ram[2582] = 240;
    exp_40_ram[2583] = 40;
    exp_40_ram[2584] = 42;
    exp_40_ram[2585] = 39;
    exp_40_ram[2586] = 94;
    exp_40_ram[2587] = 38;
    exp_40_ram[2588] = 38;
    exp_40_ram[2589] = 245;
    exp_40_ram[2590] = 5;
    exp_40_ram[2591] = 5;
    exp_40_ram[2592] = 7;
    exp_40_ram[2593] = 8;
    exp_40_ram[2594] = 56;
    exp_40_ram[2595] = 135;
    exp_40_ram[2596] = 6;
    exp_40_ram[2597] = 135;
    exp_40_ram[2598] = 44;
    exp_40_ram[2599] = 46;
    exp_40_ram[2600] = 0;
    exp_40_ram[2601] = 39;
    exp_40_ram[2602] = 210;
    exp_40_ram[2603] = 35;
    exp_40_ram[2604] = 40;
    exp_40_ram[2605] = 40;
    exp_40_ram[2606] = 37;
    exp_40_ram[2607] = 37;
    exp_40_ram[2608] = 38;
    exp_40_ram[2609] = 38;
    exp_40_ram[2610] = 39;
    exp_40_ram[2611] = 39;
    exp_40_ram[2612] = 32;
    exp_40_ram[2613] = 34;
    exp_40_ram[2614] = 36;
    exp_40_ram[2615] = 38;
    exp_40_ram[2616] = 40;
    exp_40_ram[2617] = 42;
    exp_40_ram[2618] = 44;
    exp_40_ram[2619] = 46;
    exp_40_ram[2620] = 32;
    exp_40_ram[2621] = 7;
    exp_40_ram[2622] = 133;
    exp_40_ram[2623] = 240;
    exp_40_ram[2624] = 7;
    exp_40_ram[2625] = 138;
    exp_40_ram[2626] = 22;
    exp_40_ram[2627] = 6;
    exp_40_ram[2628] = 6;
    exp_40_ram[2629] = 0;
    exp_40_ram[2630] = 6;
    exp_40_ram[2631] = 6;
    exp_40_ram[2632] = 37;
    exp_40_ram[2633] = 37;
    exp_40_ram[2634] = 7;
    exp_40_ram[2635] = 8;
    exp_40_ram[2636] = 56;
    exp_40_ram[2637] = 135;
    exp_40_ram[2638] = 134;
    exp_40_ram[2639] = 135;
    exp_40_ram[2640] = 44;
    exp_40_ram[2641] = 46;
    exp_40_ram[2642] = 0;
    exp_40_ram[2643] = 39;
    exp_40_ram[2644] = 39;
    exp_40_ram[2645] = 44;
    exp_40_ram[2646] = 46;
    exp_40_ram[2647] = 71;
    exp_40_ram[2648] = 167;
    exp_40_ram[2649] = 137;
    exp_40_ram[2650] = 215;
    exp_40_ram[2651] = 137;
    exp_40_ram[2652] = 38;
    exp_40_ram[2653] = 38;
    exp_40_ram[2654] = 7;
    exp_40_ram[2655] = 5;
    exp_40_ram[2656] = 53;
    exp_40_ram[2657] = 135;
    exp_40_ram[2658] = 134;
    exp_40_ram[2659] = 135;
    exp_40_ram[2660] = 44;
    exp_40_ram[2661] = 46;
    exp_40_ram[2662] = 36;
    exp_40_ram[2663] = 7;
    exp_40_ram[2664] = 37;
    exp_40_ram[2665] = 38;
    exp_40_ram[2666] = 133;
    exp_40_ram[2667] = 0;
    exp_40_ram[2668] = 35;
    exp_40_ram[2669] = 40;
    exp_40_ram[2670] = 40;
    exp_40_ram[2671] = 37;
    exp_40_ram[2672] = 37;
    exp_40_ram[2673] = 38;
    exp_40_ram[2674] = 38;
    exp_40_ram[2675] = 39;
    exp_40_ram[2676] = 39;
    exp_40_ram[2677] = 160;
    exp_40_ram[2678] = 162;
    exp_40_ram[2679] = 164;
    exp_40_ram[2680] = 166;
    exp_40_ram[2681] = 168;
    exp_40_ram[2682] = 170;
    exp_40_ram[2683] = 172;
    exp_40_ram[2684] = 174;
    exp_40_ram[2685] = 160;
    exp_40_ram[2686] = 39;
    exp_40_ram[2687] = 90;
    exp_40_ram[2688] = 39;
    exp_40_ram[2689] = 7;
    exp_40_ram[2690] = 160;
    exp_40_ram[2691] = 0;
    exp_40_ram[2692] = 39;
    exp_40_ram[2693] = 212;
    exp_40_ram[2694] = 35;
    exp_40_ram[2695] = 40;
    exp_40_ram[2696] = 40;
    exp_40_ram[2697] = 37;
    exp_40_ram[2698] = 37;
    exp_40_ram[2699] = 38;
    exp_40_ram[2700] = 38;
    exp_40_ram[2701] = 39;
    exp_40_ram[2702] = 39;
    exp_40_ram[2703] = 32;
    exp_40_ram[2704] = 34;
    exp_40_ram[2705] = 36;
    exp_40_ram[2706] = 38;
    exp_40_ram[2707] = 40;
    exp_40_ram[2708] = 42;
    exp_40_ram[2709] = 44;
    exp_40_ram[2710] = 46;
    exp_40_ram[2711] = 32;
    exp_40_ram[2712] = 7;
    exp_40_ram[2713] = 133;
    exp_40_ram[2714] = 240;
    exp_40_ram[2715] = 7;
    exp_40_ram[2716] = 39;
    exp_40_ram[2717] = 160;
    exp_40_ram[2718] = 0;
    exp_40_ram[2719] = 39;
    exp_40_ram[2720] = 160;
    exp_40_ram[2721] = 39;
    exp_40_ram[2722] = 39;
    exp_40_ram[2723] = 5;
    exp_40_ram[2724] = 133;
    exp_40_ram[2725] = 32;
    exp_40_ram[2726] = 36;
    exp_40_ram[2727] = 36;
    exp_40_ram[2728] = 41;
    exp_40_ram[2729] = 41;
    exp_40_ram[2730] = 1;
    exp_40_ram[2731] = 128;
    exp_40_ram[2732] = 1;
    exp_40_ram[2733] = 46;
    exp_40_ram[2734] = 44;
    exp_40_ram[2735] = 42;
    exp_40_ram[2736] = 40;
    exp_40_ram[2737] = 38;
    exp_40_ram[2738] = 36;
    exp_40_ram[2739] = 34;
    exp_40_ram[2740] = 32;
    exp_40_ram[2741] = 4;
    exp_40_ram[2742] = 38;
    exp_40_ram[2743] = 240;
    exp_40_ram[2744] = 7;
    exp_40_ram[2745] = 135;
    exp_40_ram[2746] = 70;
    exp_40_ram[2747] = 166;
    exp_40_ram[2748] = 138;
    exp_40_ram[2749] = 10;
    exp_40_ram[2750] = 6;
    exp_40_ram[2751] = 134;
    exp_40_ram[2752] = 5;
    exp_40_ram[2753] = 133;
    exp_40_ram[2754] = 208;
    exp_40_ram[2755] = 7;
    exp_40_ram[2756] = 135;
    exp_40_ram[2757] = 46;
    exp_40_ram[2758] = 71;
    exp_40_ram[2759] = 167;
    exp_40_ram[2760] = 167;
    exp_40_ram[2761] = 39;
    exp_40_ram[2762] = 135;
    exp_40_ram[2763] = 46;
    exp_40_ram[2764] = 39;
    exp_40_ram[2765] = 142;
    exp_40_ram[2766] = 39;
    exp_40_ram[2767] = 137;
    exp_40_ram[2768] = 9;
    exp_40_ram[2769] = 39;
    exp_40_ram[2770] = 160;
    exp_40_ram[2771] = 162;
    exp_40_ram[2772] = 39;
    exp_40_ram[2773] = 139;
    exp_40_ram[2774] = 11;
    exp_40_ram[2775] = 7;
    exp_40_ram[2776] = 135;
    exp_40_ram[2777] = 5;
    exp_40_ram[2778] = 133;
    exp_40_ram[2779] = 32;
    exp_40_ram[2780] = 36;
    exp_40_ram[2781] = 41;
    exp_40_ram[2782] = 41;
    exp_40_ram[2783] = 42;
    exp_40_ram[2784] = 42;
    exp_40_ram[2785] = 43;
    exp_40_ram[2786] = 43;
    exp_40_ram[2787] = 1;
    exp_40_ram[2788] = 128;
    exp_40_ram[2789] = 1;
    exp_40_ram[2790] = 38;
    exp_40_ram[2791] = 36;
    exp_40_ram[2792] = 34;
    exp_40_ram[2793] = 32;
    exp_40_ram[2794] = 4;
    exp_40_ram[2795] = 44;
    exp_40_ram[2796] = 46;
    exp_40_ram[2797] = 240;
    exp_40_ram[2798] = 7;
    exp_40_ram[2799] = 135;
    exp_40_ram[2800] = 70;
    exp_40_ram[2801] = 166;
    exp_40_ram[2802] = 137;
    exp_40_ram[2803] = 9;
    exp_40_ram[2804] = 6;
    exp_40_ram[2805] = 134;
    exp_40_ram[2806] = 5;
    exp_40_ram[2807] = 133;
    exp_40_ram[2808] = 208;
    exp_40_ram[2809] = 7;
    exp_40_ram[2810] = 135;
    exp_40_ram[2811] = 36;
    exp_40_ram[2812] = 38;
    exp_40_ram[2813] = 39;
    exp_40_ram[2814] = 39;
    exp_40_ram[2815] = 37;
    exp_40_ram[2816] = 37;
    exp_40_ram[2817] = 6;
    exp_40_ram[2818] = 8;
    exp_40_ram[2819] = 56;
    exp_40_ram[2820] = 134;
    exp_40_ram[2821] = 135;
    exp_40_ram[2822] = 134;
    exp_40_ram[2823] = 7;
    exp_40_ram[2824] = 135;
    exp_40_ram[2825] = 70;
    exp_40_ram[2826] = 164;
    exp_40_ram[2827] = 166;
    exp_40_ram[2828] = 0;
    exp_40_ram[2829] = 32;
    exp_40_ram[2830] = 36;
    exp_40_ram[2831] = 41;
    exp_40_ram[2832] = 41;
    exp_40_ram[2833] = 1;
    exp_40_ram[2834] = 128;
    exp_40_ram[2835] = 1;
    exp_40_ram[2836] = 38;
    exp_40_ram[2837] = 36;
    exp_40_ram[2838] = 4;
    exp_40_ram[2839] = 46;
    exp_40_ram[2840] = 23;
    exp_40_ram[2841] = 135;
    exp_40_ram[2842] = 165;
    exp_40_ram[2843] = 165;
    exp_40_ram[2844] = 166;
    exp_40_ram[2845] = 166;
    exp_40_ram[2846] = 167;
    exp_40_ram[2847] = 42;
    exp_40_ram[2848] = 44;
    exp_40_ram[2849] = 46;
    exp_40_ram[2850] = 32;
    exp_40_ram[2851] = 34;
    exp_40_ram[2852] = 215;
    exp_40_ram[2853] = 20;
    exp_40_ram[2854] = 23;
    exp_40_ram[2855] = 135;
    exp_40_ram[2856] = 174;
    exp_40_ram[2857] = 163;
    exp_40_ram[2858] = 168;
    exp_40_ram[2859] = 168;
    exp_40_ram[2860] = 165;
    exp_40_ram[2861] = 165;
    exp_40_ram[2862] = 166;
    exp_40_ram[2863] = 166;
    exp_40_ram[2864] = 167;
    exp_40_ram[2865] = 38;
    exp_40_ram[2866] = 40;
    exp_40_ram[2867] = 42;
    exp_40_ram[2868] = 44;
    exp_40_ram[2869] = 46;
    exp_40_ram[2870] = 32;
    exp_40_ram[2871] = 34;
    exp_40_ram[2872] = 36;
    exp_40_ram[2873] = 38;
    exp_40_ram[2874] = 199;
    exp_40_ram[2875] = 8;
    exp_40_ram[2876] = 38;
    exp_40_ram[2877] = 0;
    exp_40_ram[2878] = 39;
    exp_40_ram[2879] = 167;
    exp_40_ram[2880] = 7;
    exp_40_ram[2881] = 151;
    exp_40_ram[2882] = 135;
    exp_40_ram[2883] = 39;
    exp_40_ram[2884] = 7;
    exp_40_ram[2885] = 7;
    exp_40_ram[2886] = 7;
    exp_40_ram[2887] = 199;
    exp_40_ram[2888] = 71;
    exp_40_ram[2889] = 134;
    exp_40_ram[2890] = 39;
    exp_40_ram[2891] = 135;
    exp_40_ram[2892] = 128;
    exp_40_ram[2893] = 39;
    exp_40_ram[2894] = 135;
    exp_40_ram[2895] = 38;
    exp_40_ram[2896] = 39;
    exp_40_ram[2897] = 7;
    exp_40_ram[2898] = 216;
    exp_40_ram[2899] = 71;
    exp_40_ram[2900] = 135;
    exp_40_ram[2901] = 7;
    exp_40_ram[2902] = 129;
    exp_40_ram[2903] = 38;
    exp_40_ram[2904] = 0;
    exp_40_ram[2905] = 39;
    exp_40_ram[2906] = 167;
    exp_40_ram[2907] = 7;
    exp_40_ram[2908] = 151;
    exp_40_ram[2909] = 135;
    exp_40_ram[2910] = 39;
    exp_40_ram[2911] = 7;
    exp_40_ram[2912] = 39;
    exp_40_ram[2913] = 135;
    exp_40_ram[2914] = 6;
    exp_40_ram[2915] = 135;
    exp_40_ram[2916] = 71;
    exp_40_ram[2917] = 70;
    exp_40_ram[2918] = 134;
    exp_40_ram[2919] = 135;
    exp_40_ram[2920] = 128;
    exp_40_ram[2921] = 39;
    exp_40_ram[2922] = 135;
    exp_40_ram[2923] = 38;
    exp_40_ram[2924] = 39;
    exp_40_ram[2925] = 7;
    exp_40_ram[2926] = 214;
    exp_40_ram[2927] = 71;
    exp_40_ram[2928] = 135;
    exp_40_ram[2929] = 7;
    exp_40_ram[2930] = 131;
    exp_40_ram[2931] = 39;
    exp_40_ram[2932] = 167;
    exp_40_ram[2933] = 5;
    exp_40_ram[2934] = 133;
    exp_40_ram[2935] = 16;
    exp_40_ram[2936] = 7;
    exp_40_ram[2937] = 135;
    exp_40_ram[2938] = 34;
    exp_40_ram[2939] = 36;
    exp_40_ram[2940] = 39;
    exp_40_ram[2941] = 247;
    exp_40_ram[2942] = 135;
    exp_40_ram[2943] = 247;
    exp_40_ram[2944] = 71;
    exp_40_ram[2945] = 135;
    exp_40_ram[2946] = 132;
    exp_40_ram[2947] = 39;
    exp_40_ram[2948] = 247;
    exp_40_ram[2949] = 135;
    exp_40_ram[2950] = 247;
    exp_40_ram[2951] = 71;
    exp_40_ram[2952] = 135;
    exp_40_ram[2953] = 132;
    exp_40_ram[2954] = 71;
    exp_40_ram[2955] = 135;
    exp_40_ram[2956] = 7;
    exp_40_ram[2957] = 133;
    exp_40_ram[2958] = 39;
    exp_40_ram[2959] = 167;
    exp_40_ram[2960] = 5;
    exp_40_ram[2961] = 133;
    exp_40_ram[2962] = 16;
    exp_40_ram[2963] = 7;
    exp_40_ram[2964] = 135;
    exp_40_ram[2965] = 34;
    exp_40_ram[2966] = 36;
    exp_40_ram[2967] = 39;
    exp_40_ram[2968] = 247;
    exp_40_ram[2969] = 135;
    exp_40_ram[2970] = 247;
    exp_40_ram[2971] = 71;
    exp_40_ram[2972] = 135;
    exp_40_ram[2973] = 133;
    exp_40_ram[2974] = 39;
    exp_40_ram[2975] = 247;
    exp_40_ram[2976] = 135;
    exp_40_ram[2977] = 247;
    exp_40_ram[2978] = 71;
    exp_40_ram[2979] = 135;
    exp_40_ram[2980] = 134;
    exp_40_ram[2981] = 71;
    exp_40_ram[2982] = 135;
    exp_40_ram[2983] = 7;
    exp_40_ram[2984] = 134;
    exp_40_ram[2985] = 39;
    exp_40_ram[2986] = 167;
    exp_40_ram[2987] = 5;
    exp_40_ram[2988] = 133;
    exp_40_ram[2989] = 16;
    exp_40_ram[2990] = 7;
    exp_40_ram[2991] = 135;
    exp_40_ram[2992] = 34;
    exp_40_ram[2993] = 36;
    exp_40_ram[2994] = 39;
    exp_40_ram[2995] = 247;
    exp_40_ram[2996] = 135;
    exp_40_ram[2997] = 247;
    exp_40_ram[2998] = 71;
    exp_40_ram[2999] = 135;
    exp_40_ram[3000] = 135;
    exp_40_ram[3001] = 39;
    exp_40_ram[3002] = 247;
    exp_40_ram[3003] = 135;
    exp_40_ram[3004] = 247;
    exp_40_ram[3005] = 71;
    exp_40_ram[3006] = 135;
    exp_40_ram[3007] = 135;
    exp_40_ram[3008] = 71;
    exp_40_ram[3009] = 135;
    exp_40_ram[3010] = 7;
    exp_40_ram[3011] = 136;
    exp_40_ram[3012] = 39;
    exp_40_ram[3013] = 167;
    exp_40_ram[3014] = 5;
    exp_40_ram[3015] = 133;
    exp_40_ram[3016] = 16;
    exp_40_ram[3017] = 7;
    exp_40_ram[3018] = 135;
    exp_40_ram[3019] = 34;
    exp_40_ram[3020] = 36;
    exp_40_ram[3021] = 39;
    exp_40_ram[3022] = 247;
    exp_40_ram[3023] = 135;
    exp_40_ram[3024] = 247;
    exp_40_ram[3025] = 71;
    exp_40_ram[3026] = 135;
    exp_40_ram[3027] = 136;
    exp_40_ram[3028] = 39;
    exp_40_ram[3029] = 247;
    exp_40_ram[3030] = 135;
    exp_40_ram[3031] = 247;
    exp_40_ram[3032] = 71;
    exp_40_ram[3033] = 135;
    exp_40_ram[3034] = 137;
    exp_40_ram[3035] = 71;
    exp_40_ram[3036] = 135;
    exp_40_ram[3037] = 7;
    exp_40_ram[3038] = 137;
    exp_40_ram[3039] = 39;
    exp_40_ram[3040] = 167;
    exp_40_ram[3041] = 135;
    exp_40_ram[3042] = 5;
    exp_40_ram[3043] = 133;
    exp_40_ram[3044] = 16;
    exp_40_ram[3045] = 7;
    exp_40_ram[3046] = 135;
    exp_40_ram[3047] = 34;
    exp_40_ram[3048] = 36;
    exp_40_ram[3049] = 39;
    exp_40_ram[3050] = 247;
    exp_40_ram[3051] = 135;
    exp_40_ram[3052] = 247;
    exp_40_ram[3053] = 71;
    exp_40_ram[3054] = 135;
    exp_40_ram[3055] = 138;
    exp_40_ram[3056] = 39;
    exp_40_ram[3057] = 5;
    exp_40_ram[3058] = 133;
    exp_40_ram[3059] = 16;
    exp_40_ram[3060] = 7;
    exp_40_ram[3061] = 135;
    exp_40_ram[3062] = 34;
    exp_40_ram[3063] = 36;
    exp_40_ram[3064] = 39;
    exp_40_ram[3065] = 247;
    exp_40_ram[3066] = 135;
    exp_40_ram[3067] = 247;
    exp_40_ram[3068] = 71;
    exp_40_ram[3069] = 135;
    exp_40_ram[3070] = 138;
    exp_40_ram[3071] = 39;
    exp_40_ram[3072] = 5;
    exp_40_ram[3073] = 133;
    exp_40_ram[3074] = 16;
    exp_40_ram[3075] = 7;
    exp_40_ram[3076] = 135;
    exp_40_ram[3077] = 34;
    exp_40_ram[3078] = 36;
    exp_40_ram[3079] = 39;
    exp_40_ram[3080] = 247;
    exp_40_ram[3081] = 135;
    exp_40_ram[3082] = 247;
    exp_40_ram[3083] = 71;
    exp_40_ram[3084] = 135;
    exp_40_ram[3085] = 139;
    exp_40_ram[3086] = 39;
    exp_40_ram[3087] = 247;
    exp_40_ram[3088] = 135;
    exp_40_ram[3089] = 247;
    exp_40_ram[3090] = 71;
    exp_40_ram[3091] = 135;
    exp_40_ram[3092] = 139;
    exp_40_ram[3093] = 71;
    exp_40_ram[3094] = 135;
    exp_40_ram[3095] = 7;
    exp_40_ram[3096] = 140;
    exp_40_ram[3097] = 71;
    exp_40_ram[3098] = 135;
    exp_40_ram[3099] = 140;
    exp_40_ram[3100] = 71;
    exp_40_ram[3101] = 135;
    exp_40_ram[3102] = 133;
    exp_40_ram[3103] = 32;
    exp_40_ram[3104] = 36;
    exp_40_ram[3105] = 1;
    exp_40_ram[3106] = 128;
    exp_40_ram[3107] = 1;
    exp_40_ram[3108] = 46;
    exp_40_ram[3109] = 44;
    exp_40_ram[3110] = 4;
    exp_40_ram[3111] = 38;
    exp_40_ram[3112] = 37;
    exp_40_ram[3113] = 0;
    exp_40_ram[3114] = 7;
    exp_40_ram[3115] = 133;
    exp_40_ram[3116] = 240;
    exp_40_ram[3117] = 7;
    exp_40_ram[3118] = 133;
    exp_40_ram[3119] = 32;
    exp_40_ram[3120] = 36;
    exp_40_ram[3121] = 1;
    exp_40_ram[3122] = 128;
    exp_40_ram[3123] = 1;
    exp_40_ram[3124] = 46;
    exp_40_ram[3125] = 44;
    exp_40_ram[3126] = 42;
    exp_40_ram[3127] = 40;
    exp_40_ram[3128] = 38;
    exp_40_ram[3129] = 36;
    exp_40_ram[3130] = 34;
    exp_40_ram[3131] = 32;
    exp_40_ram[3132] = 46;
    exp_40_ram[3133] = 44;
    exp_40_ram[3134] = 4;
    exp_40_ram[3135] = 38;
    exp_40_ram[3136] = 32;
    exp_40_ram[3137] = 34;
    exp_40_ram[3138] = 7;
    exp_40_ram[3139] = 44;
    exp_40_ram[3140] = 7;
    exp_40_ram[3141] = 46;
    exp_40_ram[3142] = 39;
    exp_40_ram[3143] = 133;
    exp_40_ram[3144] = 240;
    exp_40_ram[3145] = 38;
    exp_40_ram[3146] = 39;
    exp_40_ram[3147] = 87;
    exp_40_ram[3148] = 135;
    exp_40_ram[3149] = 7;
    exp_40_ram[3150] = 36;
    exp_40_ram[3151] = 39;
    exp_40_ram[3152] = 140;
    exp_40_ram[3153] = 12;
    exp_40_ram[3154] = 39;
    exp_40_ram[3155] = 135;
    exp_40_ram[3156] = 234;
    exp_40_ram[3157] = 39;
    exp_40_ram[3158] = 135;
    exp_40_ram[3159] = 152;
    exp_40_ram[3160] = 39;
    exp_40_ram[3161] = 7;
    exp_40_ram[3162] = 238;
    exp_40_ram[3163] = 39;
    exp_40_ram[3164] = 135;
    exp_40_ram[3165] = 44;
    exp_40_ram[3166] = 39;
    exp_40_ram[3167] = 135;
    exp_40_ram[3168] = 39;
    exp_40_ram[3169] = 7;
    exp_40_ram[3170] = 46;
    exp_40_ram[3171] = 39;
    exp_40_ram[3172] = 138;
    exp_40_ram[3173] = 10;
    exp_40_ram[3174] = 38;
    exp_40_ram[3175] = 38;
    exp_40_ram[3176] = 7;
    exp_40_ram[3177] = 5;
    exp_40_ram[3178] = 53;
    exp_40_ram[3179] = 135;
    exp_40_ram[3180] = 134;
    exp_40_ram[3181] = 135;
    exp_40_ram[3182] = 32;
    exp_40_ram[3183] = 34;
    exp_40_ram[3184] = 240;
    exp_40_ram[3185] = 0;
    exp_40_ram[3186] = 42;
    exp_40_ram[3187] = 32;
    exp_40_ram[3188] = 39;
    exp_40_ram[3189] = 135;
    exp_40_ram[3190] = 39;
    exp_40_ram[3191] = 133;
    exp_40_ram[3192] = 5;
    exp_40_ram[3193] = 240;
    exp_40_ram[3194] = 38;
    exp_40_ram[3195] = 39;
    exp_40_ram[3196] = 87;
    exp_40_ram[3197] = 135;
    exp_40_ram[3198] = 7;
    exp_40_ram[3199] = 36;
    exp_40_ram[3200] = 39;
    exp_40_ram[3201] = 139;
    exp_40_ram[3202] = 11;
    exp_40_ram[3203] = 39;
    exp_40_ram[3204] = 135;
    exp_40_ram[3205] = 228;
    exp_40_ram[3206] = 39;
    exp_40_ram[3207] = 135;
    exp_40_ram[3208] = 152;
    exp_40_ram[3209] = 39;
    exp_40_ram[3210] = 7;
    exp_40_ram[3211] = 232;
    exp_40_ram[3212] = 39;
    exp_40_ram[3213] = 135;
    exp_40_ram[3214] = 42;
    exp_40_ram[3215] = 39;
    exp_40_ram[3216] = 135;
    exp_40_ram[3217] = 39;
    exp_40_ram[3218] = 7;
    exp_40_ram[3219] = 46;
    exp_40_ram[3220] = 39;
    exp_40_ram[3221] = 135;
    exp_40_ram[3222] = 39;
    exp_40_ram[3223] = 7;
    exp_40_ram[3224] = 32;
    exp_40_ram[3225] = 39;
    exp_40_ram[3226] = 137;
    exp_40_ram[3227] = 9;
    exp_40_ram[3228] = 38;
    exp_40_ram[3229] = 38;
    exp_40_ram[3230] = 7;
    exp_40_ram[3231] = 5;
    exp_40_ram[3232] = 53;
    exp_40_ram[3233] = 135;
    exp_40_ram[3234] = 134;
    exp_40_ram[3235] = 135;
    exp_40_ram[3236] = 32;
    exp_40_ram[3237] = 34;
    exp_40_ram[3238] = 240;
    exp_40_ram[3239] = 0;
    exp_40_ram[3240] = 39;
    exp_40_ram[3241] = 135;
    exp_40_ram[3242] = 44;
    exp_40_ram[3243] = 39;
    exp_40_ram[3244] = 87;
    exp_40_ram[3245] = 133;
    exp_40_ram[3246] = 5;
    exp_40_ram[3247] = 0;
    exp_40_ram[3248] = 7;
    exp_40_ram[3249] = 135;
    exp_40_ram[3250] = 46;
    exp_40_ram[3251] = 32;
    exp_40_ram[3252] = 39;
    exp_40_ram[3253] = 135;
    exp_40_ram[3254] = 40;
    exp_40_ram[3255] = 39;
    exp_40_ram[3256] = 39;
    exp_40_ram[3257] = 7;
    exp_40_ram[3258] = 46;
    exp_40_ram[3259] = 39;
    exp_40_ram[3260] = 7;
    exp_40_ram[3261] = 103;
    exp_40_ram[3262] = 46;
    exp_40_ram[3263] = 39;
    exp_40_ram[3264] = 39;
    exp_40_ram[3265] = 7;
    exp_40_ram[3266] = 32;
    exp_40_ram[3267] = 39;
    exp_40_ram[3268] = 32;
    exp_40_ram[3269] = 215;
    exp_40_ram[3270] = 34;
    exp_40_ram[3271] = 39;
    exp_40_ram[3272] = 23;
    exp_40_ram[3273] = 133;
    exp_40_ram[3274] = 5;
    exp_40_ram[3275] = 0;
    exp_40_ram[3276] = 7;
    exp_40_ram[3277] = 135;
    exp_40_ram[3278] = 46;
    exp_40_ram[3279] = 32;
    exp_40_ram[3280] = 39;
    exp_40_ram[3281] = 38;
    exp_40_ram[3282] = 39;
    exp_40_ram[3283] = 32;
    exp_40_ram[3284] = 215;
    exp_40_ram[3285] = 34;
    exp_40_ram[3286] = 39;
    exp_40_ram[3287] = 5;
    exp_40_ram[3288] = 133;
    exp_40_ram[3289] = 0;
    exp_40_ram[3290] = 7;
    exp_40_ram[3291] = 135;
    exp_40_ram[3292] = 46;
    exp_40_ram[3293] = 32;
    exp_40_ram[3294] = 39;
    exp_40_ram[3295] = 36;
    exp_40_ram[3296] = 39;
    exp_40_ram[3297] = 32;
    exp_40_ram[3298] = 215;
    exp_40_ram[3299] = 34;
    exp_40_ram[3300] = 39;
    exp_40_ram[3301] = 34;
    exp_40_ram[3302] = 39;
    exp_40_ram[3303] = 46;
    exp_40_ram[3304] = 35;
    exp_40_ram[3305] = 40;
    exp_40_ram[3306] = 40;
    exp_40_ram[3307] = 37;
    exp_40_ram[3308] = 37;
    exp_40_ram[3309] = 38;
    exp_40_ram[3310] = 38;
    exp_40_ram[3311] = 39;
    exp_40_ram[3312] = 160;
    exp_40_ram[3313] = 162;
    exp_40_ram[3314] = 164;
    exp_40_ram[3315] = 166;
    exp_40_ram[3316] = 168;
    exp_40_ram[3317] = 170;
    exp_40_ram[3318] = 172;
    exp_40_ram[3319] = 174;
    exp_40_ram[3320] = 160;
    exp_40_ram[3321] = 37;
    exp_40_ram[3322] = 32;
    exp_40_ram[3323] = 36;
    exp_40_ram[3324] = 41;
    exp_40_ram[3325] = 41;
    exp_40_ram[3326] = 42;
    exp_40_ram[3327] = 42;
    exp_40_ram[3328] = 43;
    exp_40_ram[3329] = 43;
    exp_40_ram[3330] = 44;
    exp_40_ram[3331] = 44;
    exp_40_ram[3332] = 1;
    exp_40_ram[3333] = 128;
    exp_40_ram[3334] = 1;
    exp_40_ram[3335] = 46;
    exp_40_ram[3336] = 44;
    exp_40_ram[3337] = 42;
    exp_40_ram[3338] = 40;
    exp_40_ram[3339] = 38;
    exp_40_ram[3340] = 4;
    exp_40_ram[3341] = 46;
    exp_40_ram[3342] = 7;
    exp_40_ram[3343] = 8;
    exp_40_ram[3344] = 44;
    exp_40_ram[3345] = 46;
    exp_40_ram[3346] = 39;
    exp_40_ram[3347] = 167;
    exp_40_ram[3348] = 167;
    exp_40_ram[3349] = 40;
    exp_40_ram[3350] = 42;
    exp_40_ram[3351] = 37;
    exp_40_ram[3352] = 37;
    exp_40_ram[3353] = 224;
    exp_40_ram[3354] = 7;
    exp_40_ram[3355] = 140;
    exp_40_ram[3356] = 23;
    exp_40_ram[3357] = 7;
    exp_40_ram[3358] = 7;
    exp_40_ram[3359] = 44;
    exp_40_ram[3360] = 46;
    exp_40_ram[3361] = 71;
    exp_40_ram[3362] = 167;
    exp_40_ram[3363] = 137;
    exp_40_ram[3364] = 215;
    exp_40_ram[3365] = 137;
    exp_40_ram[3366] = 38;
    exp_40_ram[3367] = 38;
    exp_40_ram[3368] = 7;
    exp_40_ram[3369] = 5;
    exp_40_ram[3370] = 181;
    exp_40_ram[3371] = 135;
    exp_40_ram[3372] = 134;
    exp_40_ram[3373] = 135;
    exp_40_ram[3374] = 5;
    exp_40_ram[3375] = 133;
    exp_40_ram[3376] = 38;
    exp_40_ram[3377] = 38;
    exp_40_ram[3378] = 7;
    exp_40_ram[3379] = 8;
    exp_40_ram[3380] = 56;
    exp_40_ram[3381] = 135;
    exp_40_ram[3382] = 6;
    exp_40_ram[3383] = 135;
    exp_40_ram[3384] = 36;
    exp_40_ram[3385] = 38;
    exp_40_ram[3386] = 71;
    exp_40_ram[3387] = 132;
    exp_40_ram[3388] = 7;
    exp_40_ram[3389] = 37;
    exp_40_ram[3390] = 38;
    exp_40_ram[3391] = 133;
    exp_40_ram[3392] = 240;
    exp_40_ram[3393] = 35;
    exp_40_ram[3394] = 40;
    exp_40_ram[3395] = 40;
    exp_40_ram[3396] = 37;
    exp_40_ram[3397] = 37;
    exp_40_ram[3398] = 38;
    exp_40_ram[3399] = 38;
    exp_40_ram[3400] = 39;
    exp_40_ram[3401] = 39;
    exp_40_ram[3402] = 160;
    exp_40_ram[3403] = 162;
    exp_40_ram[3404] = 164;
    exp_40_ram[3405] = 166;
    exp_40_ram[3406] = 168;
    exp_40_ram[3407] = 170;
    exp_40_ram[3408] = 172;
    exp_40_ram[3409] = 174;
    exp_40_ram[3410] = 160;
    exp_40_ram[3411] = 37;
    exp_40_ram[3412] = 37;
    exp_40_ram[3413] = 224;
    exp_40_ram[3414] = 7;
    exp_40_ram[3415] = 71;
    exp_40_ram[3416] = 135;
    exp_40_ram[3417] = 160;
    exp_40_ram[3418] = 71;
    exp_40_ram[3419] = 135;
    exp_40_ram[3420] = 133;
    exp_40_ram[3421] = 32;
    exp_40_ram[3422] = 36;
    exp_40_ram[3423] = 36;
    exp_40_ram[3424] = 41;
    exp_40_ram[3425] = 41;
    exp_40_ram[3426] = 1;
    exp_40_ram[3427] = 128;
    exp_40_ram[3428] = 1;
    exp_40_ram[3429] = 38;
    exp_40_ram[3430] = 36;
    exp_40_ram[3431] = 4;
    exp_40_ram[3432] = 46;
    exp_40_ram[3433] = 38;
    exp_40_ram[3434] = 37;
    exp_40_ram[3435] = 208;
    exp_40_ram[3436] = 7;
    exp_40_ram[3437] = 5;
    exp_40_ram[3438] = 71;
    exp_40_ram[3439] = 135;
    exp_40_ram[3440] = 7;
    exp_40_ram[3441] = 234;
    exp_40_ram[3442] = 39;
    exp_40_ram[3443] = 7;
    exp_40_ram[3444] = 151;
    exp_40_ram[3445] = 135;
    exp_40_ram[3446] = 151;
    exp_40_ram[3447] = 38;
    exp_40_ram[3448] = 71;
    exp_40_ram[3449] = 39;
    exp_40_ram[3450] = 7;
    exp_40_ram[3451] = 135;
    exp_40_ram[3452] = 38;
    exp_40_ram[3453] = 240;
    exp_40_ram[3454] = 0;
    exp_40_ram[3455] = 39;
    exp_40_ram[3456] = 133;
    exp_40_ram[3457] = 32;
    exp_40_ram[3458] = 36;
    exp_40_ram[3459] = 1;
    exp_40_ram[3460] = 128;
    exp_40_ram[3461] = 1;
    exp_40_ram[3462] = 38;
    exp_40_ram[3463] = 36;
    exp_40_ram[3464] = 4;
    exp_40_ram[3465] = 71;
    exp_40_ram[3466] = 167;
    exp_40_ram[3467] = 133;
    exp_40_ram[3468] = 240;
    exp_40_ram[3469] = 7;
    exp_40_ram[3470] = 133;
    exp_40_ram[3471] = 32;
    exp_40_ram[3472] = 36;
    exp_40_ram[3473] = 1;
    exp_40_ram[3474] = 128;
    exp_40_ram[3475] = 1;
    exp_40_ram[3476] = 38;
    exp_40_ram[3477] = 36;
    exp_40_ram[3478] = 34;
    exp_40_ram[3479] = 32;
    exp_40_ram[3480] = 4;
    exp_40_ram[3481] = 46;
    exp_40_ram[3482] = 224;
    exp_40_ram[3483] = 36;
    exp_40_ram[3484] = 38;
    exp_40_ram[3485] = 0;
    exp_40_ram[3486] = 224;
    exp_40_ram[3487] = 6;
    exp_40_ram[3488] = 134;
    exp_40_ram[3489] = 37;
    exp_40_ram[3490] = 37;
    exp_40_ram[3491] = 7;
    exp_40_ram[3492] = 8;
    exp_40_ram[3493] = 56;
    exp_40_ram[3494] = 135;
    exp_40_ram[3495] = 134;
    exp_40_ram[3496] = 135;
    exp_40_ram[3497] = 38;
    exp_40_ram[3498] = 137;
    exp_40_ram[3499] = 9;
    exp_40_ram[3500] = 134;
    exp_40_ram[3501] = 134;
    exp_40_ram[3502] = 224;
    exp_40_ram[3503] = 134;
    exp_40_ram[3504] = 134;
    exp_40_ram[3505] = 24;
    exp_40_ram[3506] = 6;
    exp_40_ram[3507] = 7;
    exp_40_ram[3508] = 228;
    exp_40_ram[3509] = 0;
    exp_40_ram[3510] = 133;
    exp_40_ram[3511] = 32;
    exp_40_ram[3512] = 36;
    exp_40_ram[3513] = 41;
    exp_40_ram[3514] = 41;
    exp_40_ram[3515] = 1;
    exp_40_ram[3516] = 128;
    exp_40_ram[3517] = 1;
    exp_40_ram[3518] = 38;
    exp_40_ram[3519] = 36;
    exp_40_ram[3520] = 4;
    exp_40_ram[3521] = 23;
    exp_40_ram[3522] = 133;
    exp_40_ram[3523] = 224;
    exp_40_ram[3524] = 0;
    exp_40_ram[3525] = 32;
    exp_40_ram[3526] = 36;
    exp_40_ram[3527] = 1;
    exp_40_ram[3528] = 128;
    exp_40_ram[3529] = 1;
    exp_40_ram[3530] = 46;
    exp_40_ram[3531] = 44;
    exp_40_ram[3532] = 4;
    exp_40_ram[3533] = 23;
    exp_40_ram[3534] = 133;
    exp_40_ram[3535] = 224;
    exp_40_ram[3536] = 7;
    exp_40_ram[3537] = 38;
    exp_40_ram[3538] = 36;
    exp_40_ram[3539] = 0;
    exp_40_ram[3540] = 37;
    exp_40_ram[3541] = 23;
    exp_40_ram[3542] = 133;
    exp_40_ram[3543] = 224;
    exp_40_ram[3544] = 0;
    exp_40_ram[3545] = 39;
    exp_40_ram[3546] = 151;
    exp_40_ram[3547] = 38;
    exp_40_ram[3548] = 71;
    exp_40_ram[3549] = 167;
    exp_40_ram[3550] = 133;
    exp_40_ram[3551] = 37;
    exp_40_ram[3552] = 208;
    exp_40_ram[3553] = 71;
    exp_40_ram[3554] = 167;
    exp_40_ram[3555] = 7;
    exp_40_ram[3556] = 87;
    exp_40_ram[3557] = 133;
    exp_40_ram[3558] = 240;
    exp_40_ram[3559] = 39;
    exp_40_ram[3560] = 7;
    exp_40_ram[3561] = 208;
    exp_40_ram[3562] = 0;
    exp_40_ram[3563] = 39;
    exp_40_ram[3564] = 215;
    exp_40_ram[3565] = 38;
    exp_40_ram[3566] = 71;
    exp_40_ram[3567] = 167;
    exp_40_ram[3568] = 133;
    exp_40_ram[3569] = 37;
    exp_40_ram[3570] = 208;
    exp_40_ram[3571] = 71;
    exp_40_ram[3572] = 167;
    exp_40_ram[3573] = 7;
    exp_40_ram[3574] = 87;
    exp_40_ram[3575] = 133;
    exp_40_ram[3576] = 240;
    exp_40_ram[3577] = 39;
    exp_40_ram[3578] = 7;
    exp_40_ram[3579] = 192;
    exp_40_ram[3580] = 39;
    exp_40_ram[3581] = 135;
    exp_40_ram[3582] = 36;
    exp_40_ram[3583] = 39;
    exp_40_ram[3584] = 7;
    exp_40_ram[3585] = 214;
    exp_40_ram[3586] = 71;
    exp_40_ram[3587] = 167;
    exp_40_ram[3588] = 133;
    exp_40_ram[3589] = 5;
    exp_40_ram[3590] = 208;
    exp_40_ram[3591] = 0;
    exp_40_ram[3592] = 32;
    exp_40_ram[3593] = 36;
    exp_40_ram[3594] = 1;
    exp_40_ram[3595] = 128;
    exp_40_ram[3596] = 1;
    exp_40_ram[3597] = 38;
    exp_40_ram[3598] = 36;
    exp_40_ram[3599] = 34;
    exp_40_ram[3600] = 32;
    exp_40_ram[3601] = 46;
    exp_40_ram[3602] = 44;
    exp_40_ram[3603] = 42;
    exp_40_ram[3604] = 40;
    exp_40_ram[3605] = 38;
    exp_40_ram[3606] = 36;
    exp_40_ram[3607] = 34;
    exp_40_ram[3608] = 32;
    exp_40_ram[3609] = 4;
    exp_40_ram[3610] = 7;
    exp_40_ram[3611] = 46;
    exp_40_ram[3612] = 7;
    exp_40_ram[3613] = 7;
    exp_40_ram[3614] = 40;
    exp_40_ram[3615] = 42;
    exp_40_ram[3616] = 224;
    exp_40_ram[3617] = 32;
    exp_40_ram[3618] = 34;
    exp_40_ram[3619] = 38;
    exp_40_ram[3620] = 0;
    exp_40_ram[3621] = 39;
    exp_40_ram[3622] = 87;
    exp_40_ram[3623] = 135;
    exp_40_ram[3624] = 7;
    exp_40_ram[3625] = 46;
    exp_40_ram[3626] = 39;
    exp_40_ram[3627] = 87;
    exp_40_ram[3628] = 135;
    exp_40_ram[3629] = 7;
    exp_40_ram[3630] = 46;
    exp_40_ram[3631] = 39;
    exp_40_ram[3632] = 87;
    exp_40_ram[3633] = 135;
    exp_40_ram[3634] = 7;
    exp_40_ram[3635] = 46;
    exp_40_ram[3636] = 39;
    exp_40_ram[3637] = 87;
    exp_40_ram[3638] = 135;
    exp_40_ram[3639] = 7;
    exp_40_ram[3640] = 46;
    exp_40_ram[3641] = 39;
    exp_40_ram[3642] = 135;
    exp_40_ram[3643] = 38;
    exp_40_ram[3644] = 224;
    exp_40_ram[3645] = 6;
    exp_40_ram[3646] = 134;
    exp_40_ram[3647] = 37;
    exp_40_ram[3648] = 37;
    exp_40_ram[3649] = 7;
    exp_40_ram[3650] = 8;
    exp_40_ram[3651] = 56;
    exp_40_ram[3652] = 135;
    exp_40_ram[3653] = 134;
    exp_40_ram[3654] = 135;
    exp_40_ram[3655] = 70;
    exp_40_ram[3656] = 166;
    exp_40_ram[3657] = 36;
    exp_40_ram[3658] = 38;
    exp_40_ram[3659] = 37;
    exp_40_ram[3660] = 37;
    exp_40_ram[3661] = 134;
    exp_40_ram[3662] = 134;
    exp_40_ram[3663] = 236;
    exp_40_ram[3664] = 134;
    exp_40_ram[3665] = 134;
    exp_40_ram[3666] = 24;
    exp_40_ram[3667] = 6;
    exp_40_ram[3668] = 7;
    exp_40_ram[3669] = 224;
    exp_40_ram[3670] = 37;
    exp_40_ram[3671] = 23;
    exp_40_ram[3672] = 133;
    exp_40_ram[3673] = 224;
    exp_40_ram[3674] = 224;
    exp_40_ram[3675] = 32;
    exp_40_ram[3676] = 34;
    exp_40_ram[3677] = 38;
    exp_40_ram[3678] = 0;
    exp_40_ram[3679] = 39;
    exp_40_ram[3680] = 39;
    exp_40_ram[3681] = 86;
    exp_40_ram[3682] = 134;
    exp_40_ram[3683] = 134;
    exp_40_ram[3684] = 6;
    exp_40_ram[3685] = 6;
    exp_40_ram[3686] = 6;
    exp_40_ram[3687] = 86;
    exp_40_ram[3688] = 134;
    exp_40_ram[3689] = 5;
    exp_40_ram[3690] = 57;
    exp_40_ram[3691] = 137;
    exp_40_ram[3692] = 7;
    exp_40_ram[3693] = 137;
    exp_40_ram[3694] = 40;
    exp_40_ram[3695] = 42;
    exp_40_ram[3696] = 39;
    exp_40_ram[3697] = 39;
    exp_40_ram[3698] = 86;
    exp_40_ram[3699] = 134;
    exp_40_ram[3700] = 134;
    exp_40_ram[3701] = 6;
    exp_40_ram[3702] = 6;
    exp_40_ram[3703] = 6;
    exp_40_ram[3704] = 86;
    exp_40_ram[3705] = 134;
    exp_40_ram[3706] = 5;
    exp_40_ram[3707] = 58;
    exp_40_ram[3708] = 138;
    exp_40_ram[3709] = 7;
    exp_40_ram[3710] = 138;
    exp_40_ram[3711] = 40;
    exp_40_ram[3712] = 42;
    exp_40_ram[3713] = 39;
    exp_40_ram[3714] = 39;
    exp_40_ram[3715] = 86;
    exp_40_ram[3716] = 134;
    exp_40_ram[3717] = 134;
    exp_40_ram[3718] = 6;
    exp_40_ram[3719] = 6;
    exp_40_ram[3720] = 6;
    exp_40_ram[3721] = 86;
    exp_40_ram[3722] = 134;
    exp_40_ram[3723] = 5;
    exp_40_ram[3724] = 59;
    exp_40_ram[3725] = 139;
    exp_40_ram[3726] = 7;
    exp_40_ram[3727] = 139;
    exp_40_ram[3728] = 40;
    exp_40_ram[3729] = 42;
    exp_40_ram[3730] = 39;
    exp_40_ram[3731] = 39;
    exp_40_ram[3732] = 86;
    exp_40_ram[3733] = 134;
    exp_40_ram[3734] = 134;
    exp_40_ram[3735] = 6;
    exp_40_ram[3736] = 6;
    exp_40_ram[3737] = 6;
    exp_40_ram[3738] = 86;
    exp_40_ram[3739] = 134;
    exp_40_ram[3740] = 5;
    exp_40_ram[3741] = 60;
    exp_40_ram[3742] = 140;
    exp_40_ram[3743] = 7;
    exp_40_ram[3744] = 140;
    exp_40_ram[3745] = 40;
    exp_40_ram[3746] = 42;
    exp_40_ram[3747] = 39;
    exp_40_ram[3748] = 135;
    exp_40_ram[3749] = 38;
    exp_40_ram[3750] = 224;
    exp_40_ram[3751] = 6;
    exp_40_ram[3752] = 134;
    exp_40_ram[3753] = 37;
    exp_40_ram[3754] = 37;
    exp_40_ram[3755] = 7;
    exp_40_ram[3756] = 8;
    exp_40_ram[3757] = 56;
    exp_40_ram[3758] = 135;
    exp_40_ram[3759] = 134;
    exp_40_ram[3760] = 135;
    exp_40_ram[3761] = 70;
    exp_40_ram[3762] = 166;
    exp_40_ram[3763] = 32;
    exp_40_ram[3764] = 34;
    exp_40_ram[3765] = 37;
    exp_40_ram[3766] = 37;
    exp_40_ram[3767] = 134;
    exp_40_ram[3768] = 134;
    exp_40_ram[3769] = 236;
    exp_40_ram[3770] = 134;
    exp_40_ram[3771] = 134;
    exp_40_ram[3772] = 24;
    exp_40_ram[3773] = 6;
    exp_40_ram[3774] = 7;
    exp_40_ram[3775] = 224;
    exp_40_ram[3776] = 37;
    exp_40_ram[3777] = 23;
    exp_40_ram[3778] = 133;
    exp_40_ram[3779] = 224;
    exp_40_ram[3780] = 224;
    exp_40_ram[3781] = 32;
    exp_40_ram[3782] = 34;
    exp_40_ram[3783] = 38;
    exp_40_ram[3784] = 0;
    exp_40_ram[3785] = 39;
    exp_40_ram[3786] = 87;
    exp_40_ram[3787] = 135;
    exp_40_ram[3788] = 87;
    exp_40_ram[3789] = 46;
    exp_40_ram[3790] = 39;
    exp_40_ram[3791] = 87;
    exp_40_ram[3792] = 135;
    exp_40_ram[3793] = 87;
    exp_40_ram[3794] = 46;
    exp_40_ram[3795] = 39;
    exp_40_ram[3796] = 87;
    exp_40_ram[3797] = 135;
    exp_40_ram[3798] = 87;
    exp_40_ram[3799] = 46;
    exp_40_ram[3800] = 39;
    exp_40_ram[3801] = 87;
    exp_40_ram[3802] = 135;
    exp_40_ram[3803] = 87;
    exp_40_ram[3804] = 46;
    exp_40_ram[3805] = 39;
    exp_40_ram[3806] = 135;
    exp_40_ram[3807] = 38;
    exp_40_ram[3808] = 224;
    exp_40_ram[3809] = 6;
    exp_40_ram[3810] = 134;
    exp_40_ram[3811] = 37;
    exp_40_ram[3812] = 37;
    exp_40_ram[3813] = 7;
    exp_40_ram[3814] = 8;
    exp_40_ram[3815] = 56;
    exp_40_ram[3816] = 135;
    exp_40_ram[3817] = 134;
    exp_40_ram[3818] = 135;
    exp_40_ram[3819] = 70;
    exp_40_ram[3820] = 166;
    exp_40_ram[3821] = 44;
    exp_40_ram[3822] = 46;
    exp_40_ram[3823] = 37;
    exp_40_ram[3824] = 37;
    exp_40_ram[3825] = 134;
    exp_40_ram[3826] = 134;
    exp_40_ram[3827] = 236;
    exp_40_ram[3828] = 134;
    exp_40_ram[3829] = 134;
    exp_40_ram[3830] = 24;
    exp_40_ram[3831] = 6;
    exp_40_ram[3832] = 7;
    exp_40_ram[3833] = 224;
    exp_40_ram[3834] = 37;
    exp_40_ram[3835] = 23;
    exp_40_ram[3836] = 133;
    exp_40_ram[3837] = 224;
    exp_40_ram[3838] = 224;
    exp_40_ram[3839] = 32;
    exp_40_ram[3840] = 34;
    exp_40_ram[3841] = 38;
    exp_40_ram[3842] = 0;
    exp_40_ram[3843] = 39;
    exp_40_ram[3844] = 39;
    exp_40_ram[3845] = 86;
    exp_40_ram[3846] = 6;
    exp_40_ram[3847] = 6;
    exp_40_ram[3848] = 5;
    exp_40_ram[3849] = 133;
    exp_40_ram[3850] = 192;
    exp_40_ram[3851] = 7;
    exp_40_ram[3852] = 135;
    exp_40_ram[3853] = 40;
    exp_40_ram[3854] = 42;
    exp_40_ram[3855] = 39;
    exp_40_ram[3856] = 39;
    exp_40_ram[3857] = 86;
    exp_40_ram[3858] = 6;
    exp_40_ram[3859] = 6;
    exp_40_ram[3860] = 5;
    exp_40_ram[3861] = 133;
    exp_40_ram[3862] = 192;
    exp_40_ram[3863] = 7;
    exp_40_ram[3864] = 135;
    exp_40_ram[3865] = 40;
    exp_40_ram[3866] = 42;
    exp_40_ram[3867] = 39;
    exp_40_ram[3868] = 39;
    exp_40_ram[3869] = 86;
    exp_40_ram[3870] = 6;
    exp_40_ram[3871] = 6;
    exp_40_ram[3872] = 5;
    exp_40_ram[3873] = 133;
    exp_40_ram[3874] = 192;
    exp_40_ram[3875] = 7;
    exp_40_ram[3876] = 135;
    exp_40_ram[3877] = 40;
    exp_40_ram[3878] = 42;
    exp_40_ram[3879] = 39;
    exp_40_ram[3880] = 39;
    exp_40_ram[3881] = 86;
    exp_40_ram[3882] = 6;
    exp_40_ram[3883] = 6;
    exp_40_ram[3884] = 5;
    exp_40_ram[3885] = 133;
    exp_40_ram[3886] = 192;
    exp_40_ram[3887] = 7;
    exp_40_ram[3888] = 135;
    exp_40_ram[3889] = 40;
    exp_40_ram[3890] = 42;
    exp_40_ram[3891] = 39;
    exp_40_ram[3892] = 135;
    exp_40_ram[3893] = 38;
    exp_40_ram[3894] = 224;
    exp_40_ram[3895] = 6;
    exp_40_ram[3896] = 134;
    exp_40_ram[3897] = 37;
    exp_40_ram[3898] = 37;
    exp_40_ram[3899] = 7;
    exp_40_ram[3900] = 8;
    exp_40_ram[3901] = 56;
    exp_40_ram[3902] = 135;
    exp_40_ram[3903] = 134;
    exp_40_ram[3904] = 135;
    exp_40_ram[3905] = 70;
    exp_40_ram[3906] = 166;
    exp_40_ram[3907] = 141;
    exp_40_ram[3908] = 13;
    exp_40_ram[3909] = 134;
    exp_40_ram[3910] = 134;
    exp_40_ram[3911] = 232;
    exp_40_ram[3912] = 134;
    exp_40_ram[3913] = 134;
    exp_40_ram[3914] = 24;
    exp_40_ram[3915] = 6;
    exp_40_ram[3916] = 7;
    exp_40_ram[3917] = 236;
    exp_40_ram[3918] = 37;
    exp_40_ram[3919] = 23;
    exp_40_ram[3920] = 133;
    exp_40_ram[3921] = 224;
    exp_40_ram[3922] = 0;
    exp_40_ram[3923] = 32;
    exp_40_ram[3924] = 36;
    exp_40_ram[3925] = 41;
    exp_40_ram[3926] = 41;
    exp_40_ram[3927] = 42;
    exp_40_ram[3928] = 42;
    exp_40_ram[3929] = 43;
    exp_40_ram[3930] = 43;
    exp_40_ram[3931] = 44;
    exp_40_ram[3932] = 44;
    exp_40_ram[3933] = 45;
    exp_40_ram[3934] = 45;
    exp_40_ram[3935] = 1;
    exp_40_ram[3936] = 128;
    exp_40_ram[3937] = 1;
    exp_40_ram[3938] = 46;
    exp_40_ram[3939] = 44;
    exp_40_ram[3940] = 42;
    exp_40_ram[3941] = 40;
    exp_40_ram[3942] = 38;
    exp_40_ram[3943] = 36;
    exp_40_ram[3944] = 4;
    exp_40_ram[3945] = 23;
    exp_40_ram[3946] = 133;
    exp_40_ram[3947] = 224;
    exp_40_ram[3948] = 240;
    exp_40_ram[3949] = 7;
    exp_40_ram[3950] = 135;
    exp_40_ram[3951] = 34;
    exp_40_ram[3952] = 23;
    exp_40_ram[3953] = 133;
    exp_40_ram[3954] = 224;
    exp_40_ram[3955] = 240;
    exp_40_ram[3956] = 7;
    exp_40_ram[3957] = 135;
    exp_40_ram[3958] = 32;
    exp_40_ram[3959] = 23;
    exp_40_ram[3960] = 133;
    exp_40_ram[3961] = 224;
    exp_40_ram[3962] = 240;
    exp_40_ram[3963] = 7;
    exp_40_ram[3964] = 46;
    exp_40_ram[3965] = 23;
    exp_40_ram[3966] = 133;
    exp_40_ram[3967] = 224;
    exp_40_ram[3968] = 240;
    exp_40_ram[3969] = 7;
    exp_40_ram[3970] = 44;
    exp_40_ram[3971] = 23;
    exp_40_ram[3972] = 133;
    exp_40_ram[3973] = 224;
    exp_40_ram[3974] = 240;
    exp_40_ram[3975] = 7;
    exp_40_ram[3976] = 42;
    exp_40_ram[3977] = 7;
    exp_40_ram[3978] = 40;
    exp_40_ram[3979] = 7;
    exp_40_ram[3980] = 40;
    exp_40_ram[3981] = 7;
    exp_40_ram[3982] = 133;
    exp_40_ram[3983] = 224;
    exp_40_ram[3984] = 7;
    exp_40_ram[3985] = 135;
    exp_40_ram[3986] = 36;
    exp_40_ram[3987] = 38;
    exp_40_ram[3988] = 7;
    exp_40_ram[3989] = 133;
    exp_40_ram[3990] = 224;
    exp_40_ram[3991] = 7;
    exp_40_ram[3992] = 133;
    exp_40_ram[3993] = 192;
    exp_40_ram[3994] = 7;
    exp_40_ram[3995] = 133;
    exp_40_ram[3996] = 240;
    exp_40_ram[3997] = 7;
    exp_40_ram[3998] = 133;
    exp_40_ram[3999] = 192;
    exp_40_ram[4000] = 39;
    exp_40_ram[4001] = 39;
    exp_40_ram[4002] = 5;
    exp_40_ram[4003] = 133;
    exp_40_ram[4004] = 224;
    exp_40_ram[4005] = 5;
    exp_40_ram[4006] = 224;
    exp_40_ram[4007] = 7;
    exp_40_ram[4008] = 135;
    exp_40_ram[4009] = 36;
    exp_40_ram[4010] = 38;
    exp_40_ram[4011] = 7;
    exp_40_ram[4012] = 133;
    exp_40_ram[4013] = 240;
    exp_40_ram[4014] = 7;
    exp_40_ram[4015] = 133;
    exp_40_ram[4016] = 192;
    exp_40_ram[4017] = 224;
    exp_40_ram[4018] = 44;
    exp_40_ram[4019] = 46;
    exp_40_ram[4020] = 42;
    exp_40_ram[4021] = 0;
    exp_40_ram[4022] = 0;
    exp_40_ram[4023] = 224;
    exp_40_ram[4024] = 7;
    exp_40_ram[4025] = 135;
    exp_40_ram[4026] = 38;
    exp_40_ram[4027] = 38;
    exp_40_ram[4028] = 5;
    exp_40_ram[4029] = 133;
    exp_40_ram[4030] = 224;
    exp_40_ram[4031] = 10;
    exp_40_ram[4032] = 138;
    exp_40_ram[4033] = 71;
    exp_40_ram[4034] = 167;
    exp_40_ram[4035] = 133;
    exp_40_ram[4036] = 192;
    exp_40_ram[4037] = 7;
    exp_40_ram[4038] = 135;
    exp_40_ram[4039] = 6;
    exp_40_ram[4040] = 134;
    exp_40_ram[4041] = 5;
    exp_40_ram[4042] = 133;
    exp_40_ram[4043] = 192;
    exp_40_ram[4044] = 7;
    exp_40_ram[4045] = 196;
    exp_40_ram[4046] = 71;
    exp_40_ram[4047] = 167;
    exp_40_ram[4048] = 137;
    exp_40_ram[4049] = 9;
    exp_40_ram[4050] = 38;
    exp_40_ram[4051] = 38;
    exp_40_ram[4052] = 7;
    exp_40_ram[4053] = 5;
    exp_40_ram[4054] = 181;
    exp_40_ram[4055] = 135;
    exp_40_ram[4056] = 134;
    exp_40_ram[4057] = 135;
    exp_40_ram[4058] = 44;
    exp_40_ram[4059] = 46;
    exp_40_ram[4060] = 5;
    exp_40_ram[4061] = 224;
    exp_40_ram[4062] = 7;
    exp_40_ram[4063] = 135;
    exp_40_ram[4064] = 36;
    exp_40_ram[4065] = 38;
    exp_40_ram[4066] = 7;
    exp_40_ram[4067] = 133;
    exp_40_ram[4068] = 240;
    exp_40_ram[4069] = 7;
    exp_40_ram[4070] = 133;
    exp_40_ram[4071] = 192;
    exp_40_ram[4072] = 39;
    exp_40_ram[4073] = 135;
    exp_40_ram[4074] = 42;
    exp_40_ram[4075] = 39;
    exp_40_ram[4076] = 7;
    exp_40_ram[4077] = 210;
    exp_40_ram[4078] = 0;
    exp_40_ram[4079] = 0;
    exp_40_ram[4080] = 32;
    exp_40_ram[4081] = 36;
    exp_40_ram[4082] = 41;
    exp_40_ram[4083] = 41;
    exp_40_ram[4084] = 42;
    exp_40_ram[4085] = 42;
    exp_40_ram[4086] = 1;
    exp_40_ram[4087] = 128;
    exp_40_ram[4088] = 1;
    exp_40_ram[4089] = 46;
    exp_40_ram[4090] = 44;
    exp_40_ram[4091] = 4;
    exp_40_ram[4092] = 23;
    exp_40_ram[4093] = 133;
    exp_40_ram[4094] = 208;
    exp_40_ram[4095] = 23;
    exp_40_ram[4096] = 133;
    exp_40_ram[4097] = 208;
    exp_40_ram[4098] = 23;
    exp_40_ram[4099] = 133;
    exp_40_ram[4100] = 208;
    exp_40_ram[4101] = 23;
    exp_40_ram[4102] = 133;
    exp_40_ram[4103] = 208;
    exp_40_ram[4104] = 23;
    exp_40_ram[4105] = 133;
    exp_40_ram[4106] = 208;
    exp_40_ram[4107] = 192;
    exp_40_ram[4108] = 7;
    exp_40_ram[4109] = 7;
    exp_40_ram[4110] = 71;
    exp_40_ram[4111] = 7;
    exp_40_ram[4112] = 132;
    exp_40_ram[4113] = 7;
    exp_40_ram[4114] = 68;
    exp_40_ram[4115] = 7;
    exp_40_ram[4116] = 136;
    exp_40_ram[4117] = 7;
    exp_40_ram[4118] = 76;
    exp_40_ram[4119] = 7;
    exp_40_ram[4120] = 136;
    exp_40_ram[4121] = 7;
    exp_40_ram[4122] = 136;
    exp_40_ram[4123] = 0;
    exp_40_ram[4124] = 240;
    exp_40_ram[4125] = 0;
    exp_40_ram[4126] = 240;
    exp_40_ram[4127] = 0;
    exp_40_ram[4128] = 240;
    exp_40_ram[4129] = 0;
    exp_40_ram[4130] = 240;
    exp_40_ram[4131] = 0;
    exp_40_ram[4132] = 240;
    exp_40_ram[4133] = 7;
    exp_40_ram[4134] = 135;
    exp_40_ram[4135] = 69;
    exp_40_ram[4136] = 1;
    exp_40_ram[4137] = 101;
    exp_40_ram[4138] = 76;
    exp_40_ram[4139] = 214;
    exp_40_ram[4140] = 5;
    exp_40_ram[4141] = 133;
    exp_40_ram[4142] = 1;
    exp_40_ram[4143] = 128;
    exp_40_ram[4144] = 92;
    exp_40_ram[4145] = 5;
    exp_40_ram[4146] = 133;
    exp_40_ram[4147] = 240;
    exp_40_ram[4148] = 240;
    exp_40_ram[4149] = 0;
    exp_40_ram[4150] = 0;
    exp_40_ram[4151] = 0;
    exp_40_ram[4152] = 21;
    exp_40_ram[4153] = 21;
    exp_40_ram[4154] = 21;
    exp_40_ram[4155] = 21;
    exp_40_ram[4156] = 21;
    exp_40_ram[4157] = 21;
    exp_40_ram[4158] = 21;
    exp_40_ram[4159] = 21;
    exp_40_ram[4160] = 21;
    exp_40_ram[4161] = 21;
    exp_40_ram[4162] = 21;
    exp_40_ram[4163] = 21;
    exp_40_ram[4164] = 21;
    exp_40_ram[4165] = 20;
    exp_40_ram[4166] = 21;
    exp_40_ram[4167] = 21;
    exp_40_ram[4168] = 20;
    exp_40_ram[4169] = 23;
    exp_40_ram[4170] = 23;
    exp_40_ram[4171] = 23;
    exp_40_ram[4172] = 23;
    exp_40_ram[4173] = 22;
    exp_40_ram[4174] = 23;
    exp_40_ram[4175] = 23;
    exp_40_ram[4176] = 23;
    exp_40_ram[4177] = 23;
    exp_40_ram[4178] = 23;
    exp_40_ram[4179] = 23;
    exp_40_ram[4180] = 23;
    exp_40_ram[4181] = 23;
    exp_40_ram[4182] = 23;
    exp_40_ram[4183] = 23;
    exp_40_ram[4184] = 23;
    exp_40_ram[4185] = 23;
    exp_40_ram[4186] = 23;
    exp_40_ram[4187] = 23;
    exp_40_ram[4188] = 29;
    exp_40_ram[4189] = 30;
    exp_40_ram[4190] = 30;
    exp_40_ram[4191] = 30;
    exp_40_ram[4192] = 30;
    exp_40_ram[4193] = 30;
    exp_40_ram[4194] = 30;
    exp_40_ram[4195] = 30;
    exp_40_ram[4196] = 30;
    exp_40_ram[4197] = 30;
    exp_40_ram[4198] = 30;
    exp_40_ram[4199] = 30;
    exp_40_ram[4200] = 30;
    exp_40_ram[4201] = 30;
    exp_40_ram[4202] = 30;
    exp_40_ram[4203] = 30;
    exp_40_ram[4204] = 30;
    exp_40_ram[4205] = 30;
    exp_40_ram[4206] = 30;
    exp_40_ram[4207] = 30;
    exp_40_ram[4208] = 30;
    exp_40_ram[4209] = 30;
    exp_40_ram[4210] = 30;
    exp_40_ram[4211] = 30;
    exp_40_ram[4212] = 30;
    exp_40_ram[4213] = 30;
    exp_40_ram[4214] = 30;
    exp_40_ram[4215] = 30;
    exp_40_ram[4216] = 30;
    exp_40_ram[4217] = 30;
    exp_40_ram[4218] = 30;
    exp_40_ram[4219] = 30;
    exp_40_ram[4220] = 30;
    exp_40_ram[4221] = 30;
    exp_40_ram[4222] = 30;
    exp_40_ram[4223] = 30;
    exp_40_ram[4224] = 30;
    exp_40_ram[4225] = 30;
    exp_40_ram[4226] = 30;
    exp_40_ram[4227] = 30;
    exp_40_ram[4228] = 30;
    exp_40_ram[4229] = 30;
    exp_40_ram[4230] = 30;
    exp_40_ram[4231] = 30;
    exp_40_ram[4232] = 30;
    exp_40_ram[4233] = 30;
    exp_40_ram[4234] = 30;
    exp_40_ram[4235] = 30;
    exp_40_ram[4236] = 30;
    exp_40_ram[4237] = 30;
    exp_40_ram[4238] = 30;
    exp_40_ram[4239] = 23;
    exp_40_ram[4240] = 30;
    exp_40_ram[4241] = 30;
    exp_40_ram[4242] = 30;
    exp_40_ram[4243] = 30;
    exp_40_ram[4244] = 30;
    exp_40_ram[4245] = 30;
    exp_40_ram[4246] = 30;
    exp_40_ram[4247] = 30;
    exp_40_ram[4248] = 30;
    exp_40_ram[4249] = 23;
    exp_40_ram[4250] = 27;
    exp_40_ram[4251] = 23;
    exp_40_ram[4252] = 30;
    exp_40_ram[4253] = 30;
    exp_40_ram[4254] = 30;
    exp_40_ram[4255] = 30;
    exp_40_ram[4256] = 23;
    exp_40_ram[4257] = 30;
    exp_40_ram[4258] = 30;
    exp_40_ram[4259] = 30;
    exp_40_ram[4260] = 30;
    exp_40_ram[4261] = 30;
    exp_40_ram[4262] = 23;
    exp_40_ram[4263] = 29;
    exp_40_ram[4264] = 30;
    exp_40_ram[4265] = 30;
    exp_40_ram[4266] = 28;
    exp_40_ram[4267] = 30;
    exp_40_ram[4268] = 23;
    exp_40_ram[4269] = 30;
    exp_40_ram[4270] = 30;
    exp_40_ram[4271] = 23;
    exp_40_ram[4272] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 55;
    exp_33_ram[32] = 19;
    exp_33_ram[33] = 239;
    exp_33_ram[34] = 111;
    exp_33_ram[35] = 147;
    exp_33_ram[36] = 147;
    exp_33_ram[37] = 19;
    exp_33_ram[38] = 19;
    exp_33_ram[39] = 19;
    exp_33_ram[40] = 99;
    exp_33_ram[41] = 183;
    exp_33_ram[42] = 147;
    exp_33_ram[43] = 99;
    exp_33_ram[44] = 55;
    exp_33_ram[45] = 99;
    exp_33_ram[46] = 19;
    exp_33_ram[47] = 51;
    exp_33_ram[48] = 19;
    exp_33_ram[49] = 51;
    exp_33_ram[50] = 179;
    exp_33_ram[51] = 131;
    exp_33_ram[52] = 19;
    exp_33_ram[53] = 51;
    exp_33_ram[54] = 179;
    exp_33_ram[55] = 99;
    exp_33_ram[56] = 179;
    exp_33_ram[57] = 51;
    exp_33_ram[58] = 51;
    exp_33_ram[59] = 179;
    exp_33_ram[60] = 51;
    exp_33_ram[61] = 147;
    exp_33_ram[62] = 179;
    exp_33_ram[63] = 19;
    exp_33_ram[64] = 19;
    exp_33_ram[65] = 147;
    exp_33_ram[66] = 51;
    exp_33_ram[67] = 19;
    exp_33_ram[68] = 179;
    exp_33_ram[69] = 19;
    exp_33_ram[70] = 179;
    exp_33_ram[71] = 99;
    exp_33_ram[72] = 179;
    exp_33_ram[73] = 19;
    exp_33_ram[74] = 99;
    exp_33_ram[75] = 99;
    exp_33_ram[76] = 19;
    exp_33_ram[77] = 179;
    exp_33_ram[78] = 179;
    exp_33_ram[79] = 51;
    exp_33_ram[80] = 19;
    exp_33_ram[81] = 19;
    exp_33_ram[82] = 179;
    exp_33_ram[83] = 19;
    exp_33_ram[84] = 51;
    exp_33_ram[85] = 179;
    exp_33_ram[86] = 19;
    exp_33_ram[87] = 99;
    exp_33_ram[88] = 51;
    exp_33_ram[89] = 19;
    exp_33_ram[90] = 99;
    exp_33_ram[91] = 99;
    exp_33_ram[92] = 19;
    exp_33_ram[93] = 19;
    exp_33_ram[94] = 51;
    exp_33_ram[95] = 147;
    exp_33_ram[96] = 111;
    exp_33_ram[97] = 55;
    exp_33_ram[98] = 19;
    exp_33_ram[99] = 227;
    exp_33_ram[100] = 19;
    exp_33_ram[101] = 111;
    exp_33_ram[102] = 99;
    exp_33_ram[103] = 19;
    exp_33_ram[104] = 51;
    exp_33_ram[105] = 55;
    exp_33_ram[106] = 99;
    exp_33_ram[107] = 19;
    exp_33_ram[108] = 99;
    exp_33_ram[109] = 19;
    exp_33_ram[110] = 51;
    exp_33_ram[111] = 179;
    exp_33_ram[112] = 3;
    exp_33_ram[113] = 19;
    exp_33_ram[114] = 51;
    exp_33_ram[115] = 179;
    exp_33_ram[116] = 99;
    exp_33_ram[117] = 179;
    exp_33_ram[118] = 147;
    exp_33_ram[119] = 147;
    exp_33_ram[120] = 19;
    exp_33_ram[121] = 19;
    exp_33_ram[122] = 19;
    exp_33_ram[123] = 179;
    exp_33_ram[124] = 179;
    exp_33_ram[125] = 147;
    exp_33_ram[126] = 51;
    exp_33_ram[127] = 51;
    exp_33_ram[128] = 19;
    exp_33_ram[129] = 99;
    exp_33_ram[130] = 51;
    exp_33_ram[131] = 19;
    exp_33_ram[132] = 99;
    exp_33_ram[133] = 99;
    exp_33_ram[134] = 19;
    exp_33_ram[135] = 51;
    exp_33_ram[136] = 51;
    exp_33_ram[137] = 179;
    exp_33_ram[138] = 19;
    exp_33_ram[139] = 19;
    exp_33_ram[140] = 51;
    exp_33_ram[141] = 147;
    exp_33_ram[142] = 51;
    exp_33_ram[143] = 179;
    exp_33_ram[144] = 19;
    exp_33_ram[145] = 99;
    exp_33_ram[146] = 51;
    exp_33_ram[147] = 19;
    exp_33_ram[148] = 99;
    exp_33_ram[149] = 99;
    exp_33_ram[150] = 19;
    exp_33_ram[151] = 19;
    exp_33_ram[152] = 51;
    exp_33_ram[153] = 103;
    exp_33_ram[154] = 55;
    exp_33_ram[155] = 19;
    exp_33_ram[156] = 227;
    exp_33_ram[157] = 19;
    exp_33_ram[158] = 111;
    exp_33_ram[159] = 51;
    exp_33_ram[160] = 51;
    exp_33_ram[161] = 51;
    exp_33_ram[162] = 179;
    exp_33_ram[163] = 51;
    exp_33_ram[164] = 147;
    exp_33_ram[165] = 51;
    exp_33_ram[166] = 51;
    exp_33_ram[167] = 147;
    exp_33_ram[168] = 147;
    exp_33_ram[169] = 147;
    exp_33_ram[170] = 51;
    exp_33_ram[171] = 19;
    exp_33_ram[172] = 51;
    exp_33_ram[173] = 179;
    exp_33_ram[174] = 147;
    exp_33_ram[175] = 99;
    exp_33_ram[176] = 51;
    exp_33_ram[177] = 147;
    exp_33_ram[178] = 99;
    exp_33_ram[179] = 99;
    exp_33_ram[180] = 147;
    exp_33_ram[181] = 51;
    exp_33_ram[182] = 179;
    exp_33_ram[183] = 51;
    exp_33_ram[184] = 19;
    exp_33_ram[185] = 19;
    exp_33_ram[186] = 179;
    exp_33_ram[187] = 19;
    exp_33_ram[188] = 51;
    exp_33_ram[189] = 179;
    exp_33_ram[190] = 19;
    exp_33_ram[191] = 99;
    exp_33_ram[192] = 179;
    exp_33_ram[193] = 19;
    exp_33_ram[194] = 99;
    exp_33_ram[195] = 99;
    exp_33_ram[196] = 19;
    exp_33_ram[197] = 179;
    exp_33_ram[198] = 147;
    exp_33_ram[199] = 179;
    exp_33_ram[200] = 179;
    exp_33_ram[201] = 111;
    exp_33_ram[202] = 99;
    exp_33_ram[203] = 55;
    exp_33_ram[204] = 99;
    exp_33_ram[205] = 19;
    exp_33_ram[206] = 179;
    exp_33_ram[207] = 147;
    exp_33_ram[208] = 55;
    exp_33_ram[209] = 51;
    exp_33_ram[210] = 19;
    exp_33_ram[211] = 51;
    exp_33_ram[212] = 3;
    exp_33_ram[213] = 19;
    exp_33_ram[214] = 51;
    exp_33_ram[215] = 179;
    exp_33_ram[216] = 99;
    exp_33_ram[217] = 19;
    exp_33_ram[218] = 227;
    exp_33_ram[219] = 51;
    exp_33_ram[220] = 19;
    exp_33_ram[221] = 111;
    exp_33_ram[222] = 55;
    exp_33_ram[223] = 147;
    exp_33_ram[224] = 227;
    exp_33_ram[225] = 147;
    exp_33_ram[226] = 111;
    exp_33_ram[227] = 51;
    exp_33_ram[228] = 179;
    exp_33_ram[229] = 51;
    exp_33_ram[230] = 51;
    exp_33_ram[231] = 147;
    exp_33_ram[232] = 179;
    exp_33_ram[233] = 179;
    exp_33_ram[234] = 51;
    exp_33_ram[235] = 51;
    exp_33_ram[236] = 51;
    exp_33_ram[237] = 147;
    exp_33_ram[238] = 147;
    exp_33_ram[239] = 19;
    exp_33_ram[240] = 51;
    exp_33_ram[241] = 147;
    exp_33_ram[242] = 51;
    exp_33_ram[243] = 51;
    exp_33_ram[244] = 19;
    exp_33_ram[245] = 99;
    exp_33_ram[246] = 51;
    exp_33_ram[247] = 19;
    exp_33_ram[248] = 99;
    exp_33_ram[249] = 99;
    exp_33_ram[250] = 19;
    exp_33_ram[251] = 51;
    exp_33_ram[252] = 51;
    exp_33_ram[253] = 179;
    exp_33_ram[254] = 51;
    exp_33_ram[255] = 147;
    exp_33_ram[256] = 51;
    exp_33_ram[257] = 147;
    exp_33_ram[258] = 147;
    exp_33_ram[259] = 179;
    exp_33_ram[260] = 19;
    exp_33_ram[261] = 99;
    exp_33_ram[262] = 179;
    exp_33_ram[263] = 19;
    exp_33_ram[264] = 99;
    exp_33_ram[265] = 99;
    exp_33_ram[266] = 19;
    exp_33_ram[267] = 179;
    exp_33_ram[268] = 19;
    exp_33_ram[269] = 183;
    exp_33_ram[270] = 51;
    exp_33_ram[271] = 147;
    exp_33_ram[272] = 51;
    exp_33_ram[273] = 19;
    exp_33_ram[274] = 179;
    exp_33_ram[275] = 19;
    exp_33_ram[276] = 179;
    exp_33_ram[277] = 51;
    exp_33_ram[278] = 179;
    exp_33_ram[279] = 19;
    exp_33_ram[280] = 51;
    exp_33_ram[281] = 51;
    exp_33_ram[282] = 51;
    exp_33_ram[283] = 51;
    exp_33_ram[284] = 99;
    exp_33_ram[285] = 51;
    exp_33_ram[286] = 147;
    exp_33_ram[287] = 51;
    exp_33_ram[288] = 99;
    exp_33_ram[289] = 227;
    exp_33_ram[290] = 183;
    exp_33_ram[291] = 147;
    exp_33_ram[292] = 51;
    exp_33_ram[293] = 19;
    exp_33_ram[294] = 51;
    exp_33_ram[295] = 179;
    exp_33_ram[296] = 51;
    exp_33_ram[297] = 147;
    exp_33_ram[298] = 227;
    exp_33_ram[299] = 19;
    exp_33_ram[300] = 111;
    exp_33_ram[301] = 147;
    exp_33_ram[302] = 19;
    exp_33_ram[303] = 111;
    exp_33_ram[304] = 55;
    exp_33_ram[305] = 19;
    exp_33_ram[306] = 19;
    exp_33_ram[307] = 179;
    exp_33_ram[308] = 147;
    exp_33_ram[309] = 19;
    exp_33_ram[310] = 19;
    exp_33_ram[311] = 19;
    exp_33_ram[312] = 147;
    exp_33_ram[313] = 147;
    exp_33_ram[314] = 51;
    exp_33_ram[315] = 19;
    exp_33_ram[316] = 147;
    exp_33_ram[317] = 147;
    exp_33_ram[318] = 99;
    exp_33_ram[319] = 179;
    exp_33_ram[320] = 99;
    exp_33_ram[321] = 19;
    exp_33_ram[322] = 103;
    exp_33_ram[323] = 99;
    exp_33_ram[324] = 179;
    exp_33_ram[325] = 227;
    exp_33_ram[326] = 99;
    exp_33_ram[327] = 179;
    exp_33_ram[328] = 147;
    exp_33_ram[329] = 99;
    exp_33_ram[330] = 51;
    exp_33_ram[331] = 99;
    exp_33_ram[332] = 99;
    exp_33_ram[333] = 99;
    exp_33_ram[334] = 99;
    exp_33_ram[335] = 99;
    exp_33_ram[336] = 19;
    exp_33_ram[337] = 103;
    exp_33_ram[338] = 19;
    exp_33_ram[339] = 99;
    exp_33_ram[340] = 19;
    exp_33_ram[341] = 103;
    exp_33_ram[342] = 99;
    exp_33_ram[343] = 227;
    exp_33_ram[344] = 103;
    exp_33_ram[345] = 227;
    exp_33_ram[346] = 99;
    exp_33_ram[347] = 227;
    exp_33_ram[348] = 227;
    exp_33_ram[349] = 19;
    exp_33_ram[350] = 103;
    exp_33_ram[351] = 19;
    exp_33_ram[352] = 103;
    exp_33_ram[353] = 227;
    exp_33_ram[354] = 111;
    exp_33_ram[355] = 227;
    exp_33_ram[356] = 111;
    exp_33_ram[357] = 227;
    exp_33_ram[358] = 227;
    exp_33_ram[359] = 147;
    exp_33_ram[360] = 111;
    exp_33_ram[361] = 19;
    exp_33_ram[362] = 35;
    exp_33_ram[363] = 35;
    exp_33_ram[364] = 19;
    exp_33_ram[365] = 99;
    exp_33_ram[366] = 239;
    exp_33_ram[367] = 19;
    exp_33_ram[368] = 147;
    exp_33_ram[369] = 51;
    exp_33_ram[370] = 99;
    exp_33_ram[371] = 147;
    exp_33_ram[372] = 179;
    exp_33_ram[373] = 19;
    exp_33_ram[374] = 179;
    exp_33_ram[375] = 51;
    exp_33_ram[376] = 131;
    exp_33_ram[377] = 19;
    exp_33_ram[378] = 147;
    exp_33_ram[379] = 3;
    exp_33_ram[380] = 19;
    exp_33_ram[381] = 147;
    exp_33_ram[382] = 179;
    exp_33_ram[383] = 147;
    exp_33_ram[384] = 19;
    exp_33_ram[385] = 103;
    exp_33_ram[386] = 147;
    exp_33_ram[387] = 179;
    exp_33_ram[388] = 19;
    exp_33_ram[389] = 111;
    exp_33_ram[390] = 147;
    exp_33_ram[391] = 19;
    exp_33_ram[392] = 111;
    exp_33_ram[393] = 19;
    exp_33_ram[394] = 35;
    exp_33_ram[395] = 35;
    exp_33_ram[396] = 35;
    exp_33_ram[397] = 35;
    exp_33_ram[398] = 35;
    exp_33_ram[399] = 35;
    exp_33_ram[400] = 179;
    exp_33_ram[401] = 99;
    exp_33_ram[402] = 19;
    exp_33_ram[403] = 19;
    exp_33_ram[404] = 147;
    exp_33_ram[405] = 99;
    exp_33_ram[406] = 19;
    exp_33_ram[407] = 239;
    exp_33_ram[408] = 147;
    exp_33_ram[409] = 19;
    exp_33_ram[410] = 51;
    exp_33_ram[411] = 147;
    exp_33_ram[412] = 99;
    exp_33_ram[413] = 19;
    exp_33_ram[414] = 147;
    exp_33_ram[415] = 99;
    exp_33_ram[416] = 19;
    exp_33_ram[417] = 99;
    exp_33_ram[418] = 147;
    exp_33_ram[419] = 19;
    exp_33_ram[420] = 179;
    exp_33_ram[421] = 179;
    exp_33_ram[422] = 179;
    exp_33_ram[423] = 179;
    exp_33_ram[424] = 179;
    exp_33_ram[425] = 131;
    exp_33_ram[426] = 3;
    exp_33_ram[427] = 147;
    exp_33_ram[428] = 19;
    exp_33_ram[429] = 147;
    exp_33_ram[430] = 51;
    exp_33_ram[431] = 131;
    exp_33_ram[432] = 3;
    exp_33_ram[433] = 131;
    exp_33_ram[434] = 3;
    exp_33_ram[435] = 19;
    exp_33_ram[436] = 147;
    exp_33_ram[437] = 19;
    exp_33_ram[438] = 103;
    exp_33_ram[439] = 239;
    exp_33_ram[440] = 147;
    exp_33_ram[441] = 111;
    exp_33_ram[442] = 147;
    exp_33_ram[443] = 179;
    exp_33_ram[444] = 147;
    exp_33_ram[445] = 111;
    exp_33_ram[446] = 147;
    exp_33_ram[447] = 99;
    exp_33_ram[448] = 19;
    exp_33_ram[449] = 19;
    exp_33_ram[450] = 147;
    exp_33_ram[451] = 239;
    exp_33_ram[452] = 51;
    exp_33_ram[453] = 19;
    exp_33_ram[454] = 179;
    exp_33_ram[455] = 147;
    exp_33_ram[456] = 19;
    exp_33_ram[457] = 51;
    exp_33_ram[458] = 239;
    exp_33_ram[459] = 51;
    exp_33_ram[460] = 19;
    exp_33_ram[461] = 19;
    exp_33_ram[462] = 147;
    exp_33_ram[463] = 147;
    exp_33_ram[464] = 99;
    exp_33_ram[465] = 19;
    exp_33_ram[466] = 99;
    exp_33_ram[467] = 19;
    exp_33_ram[468] = 179;
    exp_33_ram[469] = 19;
    exp_33_ram[470] = 51;
    exp_33_ram[471] = 51;
    exp_33_ram[472] = 179;
    exp_33_ram[473] = 179;
    exp_33_ram[474] = 55;
    exp_33_ram[475] = 19;
    exp_33_ram[476] = 179;
    exp_33_ram[477] = 19;
    exp_33_ram[478] = 99;
    exp_33_ram[479] = 19;
    exp_33_ram[480] = 147;
    exp_33_ram[481] = 99;
    exp_33_ram[482] = 19;
    exp_33_ram[483] = 179;
    exp_33_ram[484] = 179;
    exp_33_ram[485] = 147;
    exp_33_ram[486] = 55;
    exp_33_ram[487] = 51;
    exp_33_ram[488] = 99;
    exp_33_ram[489] = 55;
    exp_33_ram[490] = 19;
    exp_33_ram[491] = 19;
    exp_33_ram[492] = 179;
    exp_33_ram[493] = 51;
    exp_33_ram[494] = 147;
    exp_33_ram[495] = 19;
    exp_33_ram[496] = 179;
    exp_33_ram[497] = 147;
    exp_33_ram[498] = 111;
    exp_33_ram[499] = 147;
    exp_33_ram[500] = 179;
    exp_33_ram[501] = 147;
    exp_33_ram[502] = 111;
    exp_33_ram[503] = 147;
    exp_33_ram[504] = 147;
    exp_33_ram[505] = 19;
    exp_33_ram[506] = 111;
    exp_33_ram[507] = 99;
    exp_33_ram[508] = 147;
    exp_33_ram[509] = 179;
    exp_33_ram[510] = 99;
    exp_33_ram[511] = 19;
    exp_33_ram[512] = 19;
    exp_33_ram[513] = 51;
    exp_33_ram[514] = 147;
    exp_33_ram[515] = 103;
    exp_33_ram[516] = 51;
    exp_33_ram[517] = 51;
    exp_33_ram[518] = 179;
    exp_33_ram[519] = 51;
    exp_33_ram[520] = 111;
    exp_33_ram[521] = 99;
    exp_33_ram[522] = 147;
    exp_33_ram[523] = 179;
    exp_33_ram[524] = 99;
    exp_33_ram[525] = 147;
    exp_33_ram[526] = 19;
    exp_33_ram[527] = 179;
    exp_33_ram[528] = 19;
    exp_33_ram[529] = 103;
    exp_33_ram[530] = 51;
    exp_33_ram[531] = 179;
    exp_33_ram[532] = 51;
    exp_33_ram[533] = 179;
    exp_33_ram[534] = 111;
    exp_33_ram[535] = 183;
    exp_33_ram[536] = 99;
    exp_33_ram[537] = 147;
    exp_33_ram[538] = 179;
    exp_33_ram[539] = 147;
    exp_33_ram[540] = 55;
    exp_33_ram[541] = 147;
    exp_33_ram[542] = 179;
    exp_33_ram[543] = 51;
    exp_33_ram[544] = 147;
    exp_33_ram[545] = 51;
    exp_33_ram[546] = 3;
    exp_33_ram[547] = 51;
    exp_33_ram[548] = 103;
    exp_33_ram[549] = 55;
    exp_33_ram[550] = 147;
    exp_33_ram[551] = 227;
    exp_33_ram[552] = 147;
    exp_33_ram[553] = 111;
    exp_33_ram[554] = 83;
    exp_33_ram[555] = 111;
    exp_33_ram[556] = 101;
    exp_33_ram[557] = 84;
    exp_33_ram[558] = 114;
    exp_33_ram[559] = 116;
    exp_33_ram[560] = 74;
    exp_33_ram[561] = 101;
    exp_33_ram[562] = 114;
    exp_33_ram[563] = 77;
    exp_33_ram[564] = 117;
    exp_33_ram[565] = 108;
    exp_33_ram[566] = 83;
    exp_33_ram[567] = 99;
    exp_33_ram[568] = 118;
    exp_33_ram[569] = 0;
    exp_33_ram[570] = 72;
    exp_33_ram[571] = 111;
    exp_33_ram[572] = 114;
    exp_33_ram[573] = 10;
    exp_33_ram[574] = 114;
    exp_33_ram[575] = 105;
    exp_33_ram[576] = 107;
    exp_33_ram[577] = 104;
    exp_33_ram[578] = 105;
    exp_33_ram[579] = 32;
    exp_33_ram[580] = 111;
    exp_33_ram[581] = 10;
    exp_33_ram[582] = 37;
    exp_33_ram[583] = 37;
    exp_33_ram[584] = 50;
    exp_33_ram[585] = 116;
    exp_33_ram[586] = 116;
    exp_33_ram[587] = 114;
    exp_33_ram[588] = 108;
    exp_33_ram[589] = 108;
    exp_33_ram[590] = 32;
    exp_33_ram[591] = 49;
    exp_33_ram[592] = 99;
    exp_33_ram[593] = 10;
    exp_33_ram[594] = 37;
    exp_33_ram[595] = 52;
    exp_33_ram[596] = 116;
    exp_33_ram[597] = 116;
    exp_33_ram[598] = 114;
    exp_33_ram[599] = 108;
    exp_33_ram[600] = 108;
    exp_33_ram[601] = 32;
    exp_33_ram[602] = 49;
    exp_33_ram[603] = 99;
    exp_33_ram[604] = 10;
    exp_33_ram[605] = 37;
    exp_33_ram[606] = 50;
    exp_33_ram[607] = 116;
    exp_33_ram[608] = 116;
    exp_33_ram[609] = 114;
    exp_33_ram[610] = 118;
    exp_33_ram[611] = 115;
    exp_33_ram[612] = 32;
    exp_33_ram[613] = 101;
    exp_33_ram[614] = 100;
    exp_33_ram[615] = 37;
    exp_33_ram[616] = 52;
    exp_33_ram[617] = 116;
    exp_33_ram[618] = 116;
    exp_33_ram[619] = 114;
    exp_33_ram[620] = 118;
    exp_33_ram[621] = 115;
    exp_33_ram[622] = 32;
    exp_33_ram[623] = 101;
    exp_33_ram[624] = 100;
    exp_33_ram[625] = 89;
    exp_33_ram[626] = 58;
    exp_33_ram[627] = 77;
    exp_33_ram[628] = 104;
    exp_33_ram[629] = 68;
    exp_33_ram[630] = 10;
    exp_33_ram[631] = 72;
    exp_33_ram[632] = 58;
    exp_33_ram[633] = 77;
    exp_33_ram[634] = 116;
    exp_33_ram[635] = 0;
    exp_33_ram[636] = 10;
    exp_33_ram[637] = 112;
    exp_33_ram[638] = 32;
    exp_33_ram[639] = 111;
    exp_33_ram[640] = 10;
    exp_33_ram[641] = 72;
    exp_33_ram[642] = 111;
    exp_33_ram[643] = 114;
    exp_33_ram[644] = 0;
    exp_33_ram[645] = 98;
    exp_33_ram[646] = 110;
    exp_33_ram[647] = 116;
    exp_33_ram[648] = 100;
    exp_33_ram[649] = 0;
    exp_33_ram[650] = 99;
    exp_33_ram[651] = 101;
    exp_33_ram[652] = 77;
    exp_33_ram[653] = 105;
    exp_33_ram[654] = 99;
    exp_33_ram[655] = 111;
    exp_33_ram[656] = 100;
    exp_33_ram[657] = 97;
    exp_33_ram[658] = 67;
    exp_33_ram[659] = 107;
    exp_33_ram[660] = 0;
    exp_33_ram[661] = 3;
    exp_33_ram[662] = 4;
    exp_33_ram[663] = 4;
    exp_33_ram[664] = 5;
    exp_33_ram[665] = 5;
    exp_33_ram[666] = 5;
    exp_33_ram[667] = 5;
    exp_33_ram[668] = 6;
    exp_33_ram[669] = 6;
    exp_33_ram[670] = 6;
    exp_33_ram[671] = 6;
    exp_33_ram[672] = 6;
    exp_33_ram[673] = 6;
    exp_33_ram[674] = 6;
    exp_33_ram[675] = 6;
    exp_33_ram[676] = 7;
    exp_33_ram[677] = 7;
    exp_33_ram[678] = 7;
    exp_33_ram[679] = 7;
    exp_33_ram[680] = 7;
    exp_33_ram[681] = 7;
    exp_33_ram[682] = 7;
    exp_33_ram[683] = 7;
    exp_33_ram[684] = 7;
    exp_33_ram[685] = 7;
    exp_33_ram[686] = 7;
    exp_33_ram[687] = 7;
    exp_33_ram[688] = 7;
    exp_33_ram[689] = 7;
    exp_33_ram[690] = 7;
    exp_33_ram[691] = 7;
    exp_33_ram[692] = 8;
    exp_33_ram[693] = 8;
    exp_33_ram[694] = 8;
    exp_33_ram[695] = 8;
    exp_33_ram[696] = 8;
    exp_33_ram[697] = 8;
    exp_33_ram[698] = 8;
    exp_33_ram[699] = 8;
    exp_33_ram[700] = 8;
    exp_33_ram[701] = 8;
    exp_33_ram[702] = 8;
    exp_33_ram[703] = 8;
    exp_33_ram[704] = 8;
    exp_33_ram[705] = 8;
    exp_33_ram[706] = 8;
    exp_33_ram[707] = 8;
    exp_33_ram[708] = 8;
    exp_33_ram[709] = 8;
    exp_33_ram[710] = 8;
    exp_33_ram[711] = 8;
    exp_33_ram[712] = 8;
    exp_33_ram[713] = 8;
    exp_33_ram[714] = 8;
    exp_33_ram[715] = 8;
    exp_33_ram[716] = 8;
    exp_33_ram[717] = 8;
    exp_33_ram[718] = 8;
    exp_33_ram[719] = 8;
    exp_33_ram[720] = 8;
    exp_33_ram[721] = 8;
    exp_33_ram[722] = 8;
    exp_33_ram[723] = 8;
    exp_33_ram[724] = 19;
    exp_33_ram[725] = 35;
    exp_33_ram[726] = 19;
    exp_33_ram[727] = 35;
    exp_33_ram[728] = 131;
    exp_33_ram[729] = 35;
    exp_33_ram[730] = 131;
    exp_33_ram[731] = 131;
    exp_33_ram[732] = 19;
    exp_33_ram[733] = 3;
    exp_33_ram[734] = 19;
    exp_33_ram[735] = 103;
    exp_33_ram[736] = 19;
    exp_33_ram[737] = 35;
    exp_33_ram[738] = 19;
    exp_33_ram[739] = 35;
    exp_33_ram[740] = 35;
    exp_33_ram[741] = 131;
    exp_33_ram[742] = 35;
    exp_33_ram[743] = 3;
    exp_33_ram[744] = 131;
    exp_33_ram[745] = 35;
    exp_33_ram[746] = 131;
    exp_33_ram[747] = 19;
    exp_33_ram[748] = 3;
    exp_33_ram[749] = 19;
    exp_33_ram[750] = 103;
    exp_33_ram[751] = 19;
    exp_33_ram[752] = 35;
    exp_33_ram[753] = 35;
    exp_33_ram[754] = 19;
    exp_33_ram[755] = 183;
    exp_33_ram[756] = 131;
    exp_33_ram[757] = 19;
    exp_33_ram[758] = 239;
    exp_33_ram[759] = 147;
    exp_33_ram[760] = 19;
    exp_33_ram[761] = 131;
    exp_33_ram[762] = 3;
    exp_33_ram[763] = 19;
    exp_33_ram[764] = 103;
    exp_33_ram[765] = 19;
    exp_33_ram[766] = 35;
    exp_33_ram[767] = 35;
    exp_33_ram[768] = 19;
    exp_33_ram[769] = 35;
    exp_33_ram[770] = 35;
    exp_33_ram[771] = 35;
    exp_33_ram[772] = 111;
    exp_33_ram[773] = 131;
    exp_33_ram[774] = 19;
    exp_33_ram[775] = 35;
    exp_33_ram[776] = 3;
    exp_33_ram[777] = 179;
    exp_33_ram[778] = 131;
    exp_33_ram[779] = 131;
    exp_33_ram[780] = 19;
    exp_33_ram[781] = 239;
    exp_33_ram[782] = 3;
    exp_33_ram[783] = 131;
    exp_33_ram[784] = 179;
    exp_33_ram[785] = 131;
    exp_33_ram[786] = 227;
    exp_33_ram[787] = 131;
    exp_33_ram[788] = 19;
    exp_33_ram[789] = 131;
    exp_33_ram[790] = 3;
    exp_33_ram[791] = 19;
    exp_33_ram[792] = 103;
    exp_33_ram[793] = 19;
    exp_33_ram[794] = 35;
    exp_33_ram[795] = 35;
    exp_33_ram[796] = 19;
    exp_33_ram[797] = 35;
    exp_33_ram[798] = 183;
    exp_33_ram[799] = 131;
    exp_33_ram[800] = 147;
    exp_33_ram[801] = 3;
    exp_33_ram[802] = 239;
    exp_33_ram[803] = 183;
    exp_33_ram[804] = 131;
    exp_33_ram[805] = 147;
    exp_33_ram[806] = 19;
    exp_33_ram[807] = 239;
    exp_33_ram[808] = 147;
    exp_33_ram[809] = 19;
    exp_33_ram[810] = 131;
    exp_33_ram[811] = 3;
    exp_33_ram[812] = 19;
    exp_33_ram[813] = 103;
    exp_33_ram[814] = 19;
    exp_33_ram[815] = 35;
    exp_33_ram[816] = 19;
    exp_33_ram[817] = 147;
    exp_33_ram[818] = 35;
    exp_33_ram[819] = 35;
    exp_33_ram[820] = 35;
    exp_33_ram[821] = 163;
    exp_33_ram[822] = 19;
    exp_33_ram[823] = 3;
    exp_33_ram[824] = 19;
    exp_33_ram[825] = 103;
    exp_33_ram[826] = 19;
    exp_33_ram[827] = 35;
    exp_33_ram[828] = 35;
    exp_33_ram[829] = 19;
    exp_33_ram[830] = 147;
    exp_33_ram[831] = 35;
    exp_33_ram[832] = 35;
    exp_33_ram[833] = 35;
    exp_33_ram[834] = 163;
    exp_33_ram[835] = 131;
    exp_33_ram[836] = 99;
    exp_33_ram[837] = 131;
    exp_33_ram[838] = 19;
    exp_33_ram[839] = 239;
    exp_33_ram[840] = 19;
    exp_33_ram[841] = 131;
    exp_33_ram[842] = 3;
    exp_33_ram[843] = 19;
    exp_33_ram[844] = 103;
    exp_33_ram[845] = 19;
    exp_33_ram[846] = 35;
    exp_33_ram[847] = 19;
    exp_33_ram[848] = 35;
    exp_33_ram[849] = 35;
    exp_33_ram[850] = 131;
    exp_33_ram[851] = 35;
    exp_33_ram[852] = 111;
    exp_33_ram[853] = 131;
    exp_33_ram[854] = 147;
    exp_33_ram[855] = 35;
    exp_33_ram[856] = 131;
    exp_33_ram[857] = 131;
    exp_33_ram[858] = 99;
    exp_33_ram[859] = 131;
    exp_33_ram[860] = 19;
    exp_33_ram[861] = 35;
    exp_33_ram[862] = 227;
    exp_33_ram[863] = 3;
    exp_33_ram[864] = 131;
    exp_33_ram[865] = 179;
    exp_33_ram[866] = 19;
    exp_33_ram[867] = 3;
    exp_33_ram[868] = 19;
    exp_33_ram[869] = 103;
    exp_33_ram[870] = 19;
    exp_33_ram[871] = 35;
    exp_33_ram[872] = 19;
    exp_33_ram[873] = 147;
    exp_33_ram[874] = 163;
    exp_33_ram[875] = 3;
    exp_33_ram[876] = 147;
    exp_33_ram[877] = 99;
    exp_33_ram[878] = 3;
    exp_33_ram[879] = 147;
    exp_33_ram[880] = 99;
    exp_33_ram[881] = 147;
    exp_33_ram[882] = 111;
    exp_33_ram[883] = 147;
    exp_33_ram[884] = 147;
    exp_33_ram[885] = 147;
    exp_33_ram[886] = 19;
    exp_33_ram[887] = 3;
    exp_33_ram[888] = 19;
    exp_33_ram[889] = 103;
    exp_33_ram[890] = 19;
    exp_33_ram[891] = 35;
    exp_33_ram[892] = 35;
    exp_33_ram[893] = 19;
    exp_33_ram[894] = 35;
    exp_33_ram[895] = 35;
    exp_33_ram[896] = 111;
    exp_33_ram[897] = 3;
    exp_33_ram[898] = 147;
    exp_33_ram[899] = 147;
    exp_33_ram[900] = 179;
    exp_33_ram[901] = 147;
    exp_33_ram[902] = 19;
    exp_33_ram[903] = 131;
    exp_33_ram[904] = 131;
    exp_33_ram[905] = 147;
    exp_33_ram[906] = 3;
    exp_33_ram[907] = 35;
    exp_33_ram[908] = 131;
    exp_33_ram[909] = 179;
    exp_33_ram[910] = 147;
    exp_33_ram[911] = 35;
    exp_33_ram[912] = 131;
    exp_33_ram[913] = 131;
    exp_33_ram[914] = 131;
    exp_33_ram[915] = 19;
    exp_33_ram[916] = 239;
    exp_33_ram[917] = 147;
    exp_33_ram[918] = 227;
    exp_33_ram[919] = 131;
    exp_33_ram[920] = 19;
    exp_33_ram[921] = 131;
    exp_33_ram[922] = 3;
    exp_33_ram[923] = 19;
    exp_33_ram[924] = 103;
    exp_33_ram[925] = 19;
    exp_33_ram[926] = 35;
    exp_33_ram[927] = 35;
    exp_33_ram[928] = 19;
    exp_33_ram[929] = 35;
    exp_33_ram[930] = 35;
    exp_33_ram[931] = 35;
    exp_33_ram[932] = 35;
    exp_33_ram[933] = 35;
    exp_33_ram[934] = 35;
    exp_33_ram[935] = 35;
    exp_33_ram[936] = 35;
    exp_33_ram[937] = 131;
    exp_33_ram[938] = 35;
    exp_33_ram[939] = 131;
    exp_33_ram[940] = 147;
    exp_33_ram[941] = 99;
    exp_33_ram[942] = 131;
    exp_33_ram[943] = 147;
    exp_33_ram[944] = 99;
    exp_33_ram[945] = 131;
    exp_33_ram[946] = 35;
    exp_33_ram[947] = 111;
    exp_33_ram[948] = 131;
    exp_33_ram[949] = 19;
    exp_33_ram[950] = 35;
    exp_33_ram[951] = 3;
    exp_33_ram[952] = 131;
    exp_33_ram[953] = 19;
    exp_33_ram[954] = 131;
    exp_33_ram[955] = 19;
    exp_33_ram[956] = 231;
    exp_33_ram[957] = 131;
    exp_33_ram[958] = 147;
    exp_33_ram[959] = 35;
    exp_33_ram[960] = 3;
    exp_33_ram[961] = 131;
    exp_33_ram[962] = 227;
    exp_33_ram[963] = 111;
    exp_33_ram[964] = 131;
    exp_33_ram[965] = 147;
    exp_33_ram[966] = 35;
    exp_33_ram[967] = 3;
    exp_33_ram[968] = 131;
    exp_33_ram[969] = 179;
    exp_33_ram[970] = 3;
    exp_33_ram[971] = 131;
    exp_33_ram[972] = 19;
    exp_33_ram[973] = 35;
    exp_33_ram[974] = 3;
    exp_33_ram[975] = 131;
    exp_33_ram[976] = 19;
    exp_33_ram[977] = 131;
    exp_33_ram[978] = 231;
    exp_33_ram[979] = 131;
    exp_33_ram[980] = 227;
    exp_33_ram[981] = 131;
    exp_33_ram[982] = 147;
    exp_33_ram[983] = 99;
    exp_33_ram[984] = 111;
    exp_33_ram[985] = 131;
    exp_33_ram[986] = 19;
    exp_33_ram[987] = 35;
    exp_33_ram[988] = 3;
    exp_33_ram[989] = 131;
    exp_33_ram[990] = 19;
    exp_33_ram[991] = 131;
    exp_33_ram[992] = 19;
    exp_33_ram[993] = 231;
    exp_33_ram[994] = 3;
    exp_33_ram[995] = 131;
    exp_33_ram[996] = 179;
    exp_33_ram[997] = 3;
    exp_33_ram[998] = 227;
    exp_33_ram[999] = 131;
    exp_33_ram[1000] = 19;
    exp_33_ram[1001] = 131;
    exp_33_ram[1002] = 3;
    exp_33_ram[1003] = 19;
    exp_33_ram[1004] = 103;
    exp_33_ram[1005] = 19;
    exp_33_ram[1006] = 35;
    exp_33_ram[1007] = 35;
    exp_33_ram[1008] = 19;
    exp_33_ram[1009] = 35;
    exp_33_ram[1010] = 35;
    exp_33_ram[1011] = 35;
    exp_33_ram[1012] = 35;
    exp_33_ram[1013] = 35;
    exp_33_ram[1014] = 35;
    exp_33_ram[1015] = 147;
    exp_33_ram[1016] = 35;
    exp_33_ram[1017] = 163;
    exp_33_ram[1018] = 131;
    exp_33_ram[1019] = 147;
    exp_33_ram[1020] = 99;
    exp_33_ram[1021] = 131;
    exp_33_ram[1022] = 99;
    exp_33_ram[1023] = 131;
    exp_33_ram[1024] = 147;
    exp_33_ram[1025] = 99;
    exp_33_ram[1026] = 131;
    exp_33_ram[1027] = 99;
    exp_33_ram[1028] = 131;
    exp_33_ram[1029] = 147;
    exp_33_ram[1030] = 99;
    exp_33_ram[1031] = 131;
    exp_33_ram[1032] = 147;
    exp_33_ram[1033] = 35;
    exp_33_ram[1034] = 111;
    exp_33_ram[1035] = 131;
    exp_33_ram[1036] = 19;
    exp_33_ram[1037] = 35;
    exp_33_ram[1038] = 3;
    exp_33_ram[1039] = 179;
    exp_33_ram[1040] = 19;
    exp_33_ram[1041] = 35;
    exp_33_ram[1042] = 3;
    exp_33_ram[1043] = 131;
    exp_33_ram[1044] = 99;
    exp_33_ram[1045] = 3;
    exp_33_ram[1046] = 147;
    exp_33_ram[1047] = 227;
    exp_33_ram[1048] = 111;
    exp_33_ram[1049] = 131;
    exp_33_ram[1050] = 19;
    exp_33_ram[1051] = 35;
    exp_33_ram[1052] = 3;
    exp_33_ram[1053] = 179;
    exp_33_ram[1054] = 19;
    exp_33_ram[1055] = 35;
    exp_33_ram[1056] = 131;
    exp_33_ram[1057] = 147;
    exp_33_ram[1058] = 99;
    exp_33_ram[1059] = 3;
    exp_33_ram[1060] = 131;
    exp_33_ram[1061] = 99;
    exp_33_ram[1062] = 3;
    exp_33_ram[1063] = 147;
    exp_33_ram[1064] = 227;
    exp_33_ram[1065] = 131;
    exp_33_ram[1066] = 147;
    exp_33_ram[1067] = 99;
    exp_33_ram[1068] = 131;
    exp_33_ram[1069] = 147;
    exp_33_ram[1070] = 99;
    exp_33_ram[1071] = 131;
    exp_33_ram[1072] = 99;
    exp_33_ram[1073] = 3;
    exp_33_ram[1074] = 131;
    exp_33_ram[1075] = 99;
    exp_33_ram[1076] = 3;
    exp_33_ram[1077] = 131;
    exp_33_ram[1078] = 99;
    exp_33_ram[1079] = 131;
    exp_33_ram[1080] = 147;
    exp_33_ram[1081] = 35;
    exp_33_ram[1082] = 131;
    exp_33_ram[1083] = 99;
    exp_33_ram[1084] = 3;
    exp_33_ram[1085] = 147;
    exp_33_ram[1086] = 99;
    exp_33_ram[1087] = 131;
    exp_33_ram[1088] = 147;
    exp_33_ram[1089] = 35;
    exp_33_ram[1090] = 3;
    exp_33_ram[1091] = 147;
    exp_33_ram[1092] = 99;
    exp_33_ram[1093] = 131;
    exp_33_ram[1094] = 147;
    exp_33_ram[1095] = 99;
    exp_33_ram[1096] = 3;
    exp_33_ram[1097] = 147;
    exp_33_ram[1098] = 99;
    exp_33_ram[1099] = 131;
    exp_33_ram[1100] = 19;
    exp_33_ram[1101] = 35;
    exp_33_ram[1102] = 3;
    exp_33_ram[1103] = 179;
    exp_33_ram[1104] = 19;
    exp_33_ram[1105] = 35;
    exp_33_ram[1106] = 111;
    exp_33_ram[1107] = 3;
    exp_33_ram[1108] = 147;
    exp_33_ram[1109] = 99;
    exp_33_ram[1110] = 131;
    exp_33_ram[1111] = 147;
    exp_33_ram[1112] = 99;
    exp_33_ram[1113] = 3;
    exp_33_ram[1114] = 147;
    exp_33_ram[1115] = 99;
    exp_33_ram[1116] = 131;
    exp_33_ram[1117] = 19;
    exp_33_ram[1118] = 35;
    exp_33_ram[1119] = 3;
    exp_33_ram[1120] = 179;
    exp_33_ram[1121] = 19;
    exp_33_ram[1122] = 35;
    exp_33_ram[1123] = 111;
    exp_33_ram[1124] = 3;
    exp_33_ram[1125] = 147;
    exp_33_ram[1126] = 99;
    exp_33_ram[1127] = 3;
    exp_33_ram[1128] = 147;
    exp_33_ram[1129] = 99;
    exp_33_ram[1130] = 131;
    exp_33_ram[1131] = 19;
    exp_33_ram[1132] = 35;
    exp_33_ram[1133] = 3;
    exp_33_ram[1134] = 179;
    exp_33_ram[1135] = 19;
    exp_33_ram[1136] = 35;
    exp_33_ram[1137] = 3;
    exp_33_ram[1138] = 147;
    exp_33_ram[1139] = 99;
    exp_33_ram[1140] = 131;
    exp_33_ram[1141] = 19;
    exp_33_ram[1142] = 35;
    exp_33_ram[1143] = 3;
    exp_33_ram[1144] = 179;
    exp_33_ram[1145] = 19;
    exp_33_ram[1146] = 35;
    exp_33_ram[1147] = 3;
    exp_33_ram[1148] = 147;
    exp_33_ram[1149] = 99;
    exp_33_ram[1150] = 131;
    exp_33_ram[1151] = 99;
    exp_33_ram[1152] = 131;
    exp_33_ram[1153] = 19;
    exp_33_ram[1154] = 35;
    exp_33_ram[1155] = 3;
    exp_33_ram[1156] = 179;
    exp_33_ram[1157] = 19;
    exp_33_ram[1158] = 35;
    exp_33_ram[1159] = 111;
    exp_33_ram[1160] = 131;
    exp_33_ram[1161] = 147;
    exp_33_ram[1162] = 99;
    exp_33_ram[1163] = 131;
    exp_33_ram[1164] = 19;
    exp_33_ram[1165] = 35;
    exp_33_ram[1166] = 3;
    exp_33_ram[1167] = 179;
    exp_33_ram[1168] = 19;
    exp_33_ram[1169] = 35;
    exp_33_ram[1170] = 111;
    exp_33_ram[1171] = 131;
    exp_33_ram[1172] = 147;
    exp_33_ram[1173] = 99;
    exp_33_ram[1174] = 131;
    exp_33_ram[1175] = 19;
    exp_33_ram[1176] = 35;
    exp_33_ram[1177] = 3;
    exp_33_ram[1178] = 179;
    exp_33_ram[1179] = 19;
    exp_33_ram[1180] = 35;
    exp_33_ram[1181] = 131;
    exp_33_ram[1182] = 3;
    exp_33_ram[1183] = 131;
    exp_33_ram[1184] = 3;
    exp_33_ram[1185] = 131;
    exp_33_ram[1186] = 3;
    exp_33_ram[1187] = 131;
    exp_33_ram[1188] = 3;
    exp_33_ram[1189] = 239;
    exp_33_ram[1190] = 147;
    exp_33_ram[1191] = 19;
    exp_33_ram[1192] = 131;
    exp_33_ram[1193] = 3;
    exp_33_ram[1194] = 19;
    exp_33_ram[1195] = 103;
    exp_33_ram[1196] = 19;
    exp_33_ram[1197] = 35;
    exp_33_ram[1198] = 35;
    exp_33_ram[1199] = 19;
    exp_33_ram[1200] = 35;
    exp_33_ram[1201] = 35;
    exp_33_ram[1202] = 35;
    exp_33_ram[1203] = 35;
    exp_33_ram[1204] = 35;
    exp_33_ram[1205] = 35;
    exp_33_ram[1206] = 35;
    exp_33_ram[1207] = 163;
    exp_33_ram[1208] = 35;
    exp_33_ram[1209] = 131;
    exp_33_ram[1210] = 99;
    exp_33_ram[1211] = 131;
    exp_33_ram[1212] = 147;
    exp_33_ram[1213] = 35;
    exp_33_ram[1214] = 131;
    exp_33_ram[1215] = 147;
    exp_33_ram[1216] = 99;
    exp_33_ram[1217] = 131;
    exp_33_ram[1218] = 99;
    exp_33_ram[1219] = 3;
    exp_33_ram[1220] = 131;
    exp_33_ram[1221] = 179;
    exp_33_ram[1222] = 163;
    exp_33_ram[1223] = 3;
    exp_33_ram[1224] = 147;
    exp_33_ram[1225] = 99;
    exp_33_ram[1226] = 131;
    exp_33_ram[1227] = 147;
    exp_33_ram[1228] = 147;
    exp_33_ram[1229] = 111;
    exp_33_ram[1230] = 131;
    exp_33_ram[1231] = 147;
    exp_33_ram[1232] = 99;
    exp_33_ram[1233] = 147;
    exp_33_ram[1234] = 111;
    exp_33_ram[1235] = 147;
    exp_33_ram[1236] = 3;
    exp_33_ram[1237] = 179;
    exp_33_ram[1238] = 147;
    exp_33_ram[1239] = 147;
    exp_33_ram[1240] = 147;
    exp_33_ram[1241] = 3;
    exp_33_ram[1242] = 147;
    exp_33_ram[1243] = 35;
    exp_33_ram[1244] = 147;
    exp_33_ram[1245] = 51;
    exp_33_ram[1246] = 35;
    exp_33_ram[1247] = 3;
    exp_33_ram[1248] = 131;
    exp_33_ram[1249] = 179;
    exp_33_ram[1250] = 35;
    exp_33_ram[1251] = 131;
    exp_33_ram[1252] = 99;
    exp_33_ram[1253] = 3;
    exp_33_ram[1254] = 147;
    exp_33_ram[1255] = 227;
    exp_33_ram[1256] = 131;
    exp_33_ram[1257] = 19;
    exp_33_ram[1258] = 131;
    exp_33_ram[1259] = 35;
    exp_33_ram[1260] = 131;
    exp_33_ram[1261] = 35;
    exp_33_ram[1262] = 131;
    exp_33_ram[1263] = 35;
    exp_33_ram[1264] = 131;
    exp_33_ram[1265] = 19;
    exp_33_ram[1266] = 131;
    exp_33_ram[1267] = 131;
    exp_33_ram[1268] = 3;
    exp_33_ram[1269] = 131;
    exp_33_ram[1270] = 3;
    exp_33_ram[1271] = 239;
    exp_33_ram[1272] = 147;
    exp_33_ram[1273] = 19;
    exp_33_ram[1274] = 131;
    exp_33_ram[1275] = 3;
    exp_33_ram[1276] = 19;
    exp_33_ram[1277] = 103;
    exp_33_ram[1278] = 19;
    exp_33_ram[1279] = 35;
    exp_33_ram[1280] = 35;
    exp_33_ram[1281] = 19;
    exp_33_ram[1282] = 35;
    exp_33_ram[1283] = 35;
    exp_33_ram[1284] = 35;
    exp_33_ram[1285] = 35;
    exp_33_ram[1286] = 35;
    exp_33_ram[1287] = 35;
    exp_33_ram[1288] = 131;
    exp_33_ram[1289] = 227;
    exp_33_ram[1290] = 183;
    exp_33_ram[1291] = 147;
    exp_33_ram[1292] = 35;
    exp_33_ram[1293] = 111;
    exp_33_ram[1294] = 131;
    exp_33_ram[1295] = 3;
    exp_33_ram[1296] = 147;
    exp_33_ram[1297] = 99;
    exp_33_ram[1298] = 131;
    exp_33_ram[1299] = 3;
    exp_33_ram[1300] = 131;
    exp_33_ram[1301] = 19;
    exp_33_ram[1302] = 35;
    exp_33_ram[1303] = 3;
    exp_33_ram[1304] = 131;
    exp_33_ram[1305] = 19;
    exp_33_ram[1306] = 131;
    exp_33_ram[1307] = 231;
    exp_33_ram[1308] = 131;
    exp_33_ram[1309] = 147;
    exp_33_ram[1310] = 35;
    exp_33_ram[1311] = 111;
    exp_33_ram[1312] = 131;
    exp_33_ram[1313] = 147;
    exp_33_ram[1314] = 35;
    exp_33_ram[1315] = 35;
    exp_33_ram[1316] = 131;
    exp_33_ram[1317] = 131;
    exp_33_ram[1318] = 147;
    exp_33_ram[1319] = 19;
    exp_33_ram[1320] = 99;
    exp_33_ram[1321] = 19;
    exp_33_ram[1322] = 183;
    exp_33_ram[1323] = 147;
    exp_33_ram[1324] = 179;
    exp_33_ram[1325] = 131;
    exp_33_ram[1326] = 103;
    exp_33_ram[1327] = 131;
    exp_33_ram[1328] = 147;
    exp_33_ram[1329] = 35;
    exp_33_ram[1330] = 131;
    exp_33_ram[1331] = 147;
    exp_33_ram[1332] = 35;
    exp_33_ram[1333] = 147;
    exp_33_ram[1334] = 35;
    exp_33_ram[1335] = 111;
    exp_33_ram[1336] = 131;
    exp_33_ram[1337] = 147;
    exp_33_ram[1338] = 35;
    exp_33_ram[1339] = 131;
    exp_33_ram[1340] = 147;
    exp_33_ram[1341] = 35;
    exp_33_ram[1342] = 147;
    exp_33_ram[1343] = 35;
    exp_33_ram[1344] = 111;
    exp_33_ram[1345] = 131;
    exp_33_ram[1346] = 147;
    exp_33_ram[1347] = 35;
    exp_33_ram[1348] = 131;
    exp_33_ram[1349] = 147;
    exp_33_ram[1350] = 35;
    exp_33_ram[1351] = 147;
    exp_33_ram[1352] = 35;
    exp_33_ram[1353] = 111;
    exp_33_ram[1354] = 131;
    exp_33_ram[1355] = 147;
    exp_33_ram[1356] = 35;
    exp_33_ram[1357] = 131;
    exp_33_ram[1358] = 147;
    exp_33_ram[1359] = 35;
    exp_33_ram[1360] = 147;
    exp_33_ram[1361] = 35;
    exp_33_ram[1362] = 111;
    exp_33_ram[1363] = 131;
    exp_33_ram[1364] = 147;
    exp_33_ram[1365] = 35;
    exp_33_ram[1366] = 131;
    exp_33_ram[1367] = 147;
    exp_33_ram[1368] = 35;
    exp_33_ram[1369] = 147;
    exp_33_ram[1370] = 35;
    exp_33_ram[1371] = 111;
    exp_33_ram[1372] = 35;
    exp_33_ram[1373] = 19;
    exp_33_ram[1374] = 131;
    exp_33_ram[1375] = 227;
    exp_33_ram[1376] = 35;
    exp_33_ram[1377] = 131;
    exp_33_ram[1378] = 131;
    exp_33_ram[1379] = 19;
    exp_33_ram[1380] = 239;
    exp_33_ram[1381] = 147;
    exp_33_ram[1382] = 99;
    exp_33_ram[1383] = 147;
    exp_33_ram[1384] = 19;
    exp_33_ram[1385] = 239;
    exp_33_ram[1386] = 35;
    exp_33_ram[1387] = 111;
    exp_33_ram[1388] = 131;
    exp_33_ram[1389] = 3;
    exp_33_ram[1390] = 147;
    exp_33_ram[1391] = 99;
    exp_33_ram[1392] = 131;
    exp_33_ram[1393] = 19;
    exp_33_ram[1394] = 35;
    exp_33_ram[1395] = 131;
    exp_33_ram[1396] = 35;
    exp_33_ram[1397] = 131;
    exp_33_ram[1398] = 99;
    exp_33_ram[1399] = 131;
    exp_33_ram[1400] = 147;
    exp_33_ram[1401] = 35;
    exp_33_ram[1402] = 131;
    exp_33_ram[1403] = 179;
    exp_33_ram[1404] = 35;
    exp_33_ram[1405] = 111;
    exp_33_ram[1406] = 131;
    exp_33_ram[1407] = 35;
    exp_33_ram[1408] = 131;
    exp_33_ram[1409] = 147;
    exp_33_ram[1410] = 35;
    exp_33_ram[1411] = 35;
    exp_33_ram[1412] = 131;
    exp_33_ram[1413] = 3;
    exp_33_ram[1414] = 147;
    exp_33_ram[1415] = 99;
    exp_33_ram[1416] = 131;
    exp_33_ram[1417] = 147;
    exp_33_ram[1418] = 35;
    exp_33_ram[1419] = 131;
    exp_33_ram[1420] = 147;
    exp_33_ram[1421] = 35;
    exp_33_ram[1422] = 131;
    exp_33_ram[1423] = 131;
    exp_33_ram[1424] = 19;
    exp_33_ram[1425] = 239;
    exp_33_ram[1426] = 147;
    exp_33_ram[1427] = 99;
    exp_33_ram[1428] = 147;
    exp_33_ram[1429] = 19;
    exp_33_ram[1430] = 239;
    exp_33_ram[1431] = 35;
    exp_33_ram[1432] = 111;
    exp_33_ram[1433] = 131;
    exp_33_ram[1434] = 3;
    exp_33_ram[1435] = 147;
    exp_33_ram[1436] = 99;
    exp_33_ram[1437] = 131;
    exp_33_ram[1438] = 19;
    exp_33_ram[1439] = 35;
    exp_33_ram[1440] = 131;
    exp_33_ram[1441] = 35;
    exp_33_ram[1442] = 131;
    exp_33_ram[1443] = 99;
    exp_33_ram[1444] = 147;
    exp_33_ram[1445] = 35;
    exp_33_ram[1446] = 131;
    exp_33_ram[1447] = 147;
    exp_33_ram[1448] = 35;
    exp_33_ram[1449] = 131;
    exp_33_ram[1450] = 131;
    exp_33_ram[1451] = 147;
    exp_33_ram[1452] = 19;
    exp_33_ram[1453] = 99;
    exp_33_ram[1454] = 19;
    exp_33_ram[1455] = 183;
    exp_33_ram[1456] = 147;
    exp_33_ram[1457] = 179;
    exp_33_ram[1458] = 131;
    exp_33_ram[1459] = 103;
    exp_33_ram[1460] = 131;
    exp_33_ram[1461] = 147;
    exp_33_ram[1462] = 35;
    exp_33_ram[1463] = 131;
    exp_33_ram[1464] = 147;
    exp_33_ram[1465] = 35;
    exp_33_ram[1466] = 131;
    exp_33_ram[1467] = 3;
    exp_33_ram[1468] = 147;
    exp_33_ram[1469] = 99;
    exp_33_ram[1470] = 131;
    exp_33_ram[1471] = 147;
    exp_33_ram[1472] = 35;
    exp_33_ram[1473] = 131;
    exp_33_ram[1474] = 147;
    exp_33_ram[1475] = 35;
    exp_33_ram[1476] = 111;
    exp_33_ram[1477] = 131;
    exp_33_ram[1478] = 147;
    exp_33_ram[1479] = 35;
    exp_33_ram[1480] = 131;
    exp_33_ram[1481] = 147;
    exp_33_ram[1482] = 35;
    exp_33_ram[1483] = 131;
    exp_33_ram[1484] = 3;
    exp_33_ram[1485] = 147;
    exp_33_ram[1486] = 99;
    exp_33_ram[1487] = 131;
    exp_33_ram[1488] = 147;
    exp_33_ram[1489] = 35;
    exp_33_ram[1490] = 131;
    exp_33_ram[1491] = 147;
    exp_33_ram[1492] = 35;
    exp_33_ram[1493] = 111;
    exp_33_ram[1494] = 131;
    exp_33_ram[1495] = 147;
    exp_33_ram[1496] = 35;
    exp_33_ram[1497] = 131;
    exp_33_ram[1498] = 147;
    exp_33_ram[1499] = 35;
    exp_33_ram[1500] = 111;
    exp_33_ram[1501] = 131;
    exp_33_ram[1502] = 147;
    exp_33_ram[1503] = 35;
    exp_33_ram[1504] = 131;
    exp_33_ram[1505] = 147;
    exp_33_ram[1506] = 35;
    exp_33_ram[1507] = 111;
    exp_33_ram[1508] = 131;
    exp_33_ram[1509] = 147;
    exp_33_ram[1510] = 35;
    exp_33_ram[1511] = 131;
    exp_33_ram[1512] = 147;
    exp_33_ram[1513] = 35;
    exp_33_ram[1514] = 111;
    exp_33_ram[1515] = 19;
    exp_33_ram[1516] = 111;
    exp_33_ram[1517] = 19;
    exp_33_ram[1518] = 111;
    exp_33_ram[1519] = 19;
    exp_33_ram[1520] = 131;
    exp_33_ram[1521] = 131;
    exp_33_ram[1522] = 147;
    exp_33_ram[1523] = 19;
    exp_33_ram[1524] = 99;
    exp_33_ram[1525] = 19;
    exp_33_ram[1526] = 183;
    exp_33_ram[1527] = 147;
    exp_33_ram[1528] = 179;
    exp_33_ram[1529] = 131;
    exp_33_ram[1530] = 103;
    exp_33_ram[1531] = 131;
    exp_33_ram[1532] = 3;
    exp_33_ram[1533] = 147;
    exp_33_ram[1534] = 99;
    exp_33_ram[1535] = 131;
    exp_33_ram[1536] = 3;
    exp_33_ram[1537] = 147;
    exp_33_ram[1538] = 99;
    exp_33_ram[1539] = 147;
    exp_33_ram[1540] = 35;
    exp_33_ram[1541] = 111;
    exp_33_ram[1542] = 131;
    exp_33_ram[1543] = 3;
    exp_33_ram[1544] = 147;
    exp_33_ram[1545] = 99;
    exp_33_ram[1546] = 147;
    exp_33_ram[1547] = 35;
    exp_33_ram[1548] = 111;
    exp_33_ram[1549] = 131;
    exp_33_ram[1550] = 3;
    exp_33_ram[1551] = 147;
    exp_33_ram[1552] = 99;
    exp_33_ram[1553] = 147;
    exp_33_ram[1554] = 35;
    exp_33_ram[1555] = 111;
    exp_33_ram[1556] = 147;
    exp_33_ram[1557] = 35;
    exp_33_ram[1558] = 131;
    exp_33_ram[1559] = 147;
    exp_33_ram[1560] = 35;
    exp_33_ram[1561] = 131;
    exp_33_ram[1562] = 3;
    exp_33_ram[1563] = 147;
    exp_33_ram[1564] = 99;
    exp_33_ram[1565] = 131;
    exp_33_ram[1566] = 147;
    exp_33_ram[1567] = 35;
    exp_33_ram[1568] = 131;
    exp_33_ram[1569] = 3;
    exp_33_ram[1570] = 147;
    exp_33_ram[1571] = 99;
    exp_33_ram[1572] = 131;
    exp_33_ram[1573] = 3;
    exp_33_ram[1574] = 147;
    exp_33_ram[1575] = 99;
    exp_33_ram[1576] = 131;
    exp_33_ram[1577] = 147;
    exp_33_ram[1578] = 35;
    exp_33_ram[1579] = 131;
    exp_33_ram[1580] = 147;
    exp_33_ram[1581] = 99;
    exp_33_ram[1582] = 131;
    exp_33_ram[1583] = 147;
    exp_33_ram[1584] = 35;
    exp_33_ram[1585] = 131;
    exp_33_ram[1586] = 3;
    exp_33_ram[1587] = 147;
    exp_33_ram[1588] = 99;
    exp_33_ram[1589] = 131;
    exp_33_ram[1590] = 3;
    exp_33_ram[1591] = 147;
    exp_33_ram[1592] = 99;
    exp_33_ram[1593] = 131;
    exp_33_ram[1594] = 147;
    exp_33_ram[1595] = 99;
    exp_33_ram[1596] = 131;
    exp_33_ram[1597] = 147;
    exp_33_ram[1598] = 99;
    exp_33_ram[1599] = 131;
    exp_33_ram[1600] = 19;
    exp_33_ram[1601] = 35;
    exp_33_ram[1602] = 131;
    exp_33_ram[1603] = 35;
    exp_33_ram[1604] = 131;
    exp_33_ram[1605] = 19;
    exp_33_ram[1606] = 131;
    exp_33_ram[1607] = 179;
    exp_33_ram[1608] = 179;
    exp_33_ram[1609] = 147;
    exp_33_ram[1610] = 131;
    exp_33_ram[1611] = 147;
    exp_33_ram[1612] = 19;
    exp_33_ram[1613] = 131;
    exp_33_ram[1614] = 35;
    exp_33_ram[1615] = 131;
    exp_33_ram[1616] = 35;
    exp_33_ram[1617] = 131;
    exp_33_ram[1618] = 3;
    exp_33_ram[1619] = 147;
    exp_33_ram[1620] = 19;
    exp_33_ram[1621] = 131;
    exp_33_ram[1622] = 3;
    exp_33_ram[1623] = 131;
    exp_33_ram[1624] = 3;
    exp_33_ram[1625] = 239;
    exp_33_ram[1626] = 35;
    exp_33_ram[1627] = 111;
    exp_33_ram[1628] = 131;
    exp_33_ram[1629] = 147;
    exp_33_ram[1630] = 99;
    exp_33_ram[1631] = 131;
    exp_33_ram[1632] = 19;
    exp_33_ram[1633] = 35;
    exp_33_ram[1634] = 131;
    exp_33_ram[1635] = 147;
    exp_33_ram[1636] = 111;
    exp_33_ram[1637] = 131;
    exp_33_ram[1638] = 147;
    exp_33_ram[1639] = 99;
    exp_33_ram[1640] = 131;
    exp_33_ram[1641] = 19;
    exp_33_ram[1642] = 35;
    exp_33_ram[1643] = 131;
    exp_33_ram[1644] = 147;
    exp_33_ram[1645] = 147;
    exp_33_ram[1646] = 111;
    exp_33_ram[1647] = 131;
    exp_33_ram[1648] = 19;
    exp_33_ram[1649] = 35;
    exp_33_ram[1650] = 131;
    exp_33_ram[1651] = 35;
    exp_33_ram[1652] = 131;
    exp_33_ram[1653] = 19;
    exp_33_ram[1654] = 131;
    exp_33_ram[1655] = 179;
    exp_33_ram[1656] = 179;
    exp_33_ram[1657] = 147;
    exp_33_ram[1658] = 131;
    exp_33_ram[1659] = 147;
    exp_33_ram[1660] = 19;
    exp_33_ram[1661] = 131;
    exp_33_ram[1662] = 35;
    exp_33_ram[1663] = 131;
    exp_33_ram[1664] = 35;
    exp_33_ram[1665] = 131;
    exp_33_ram[1666] = 3;
    exp_33_ram[1667] = 147;
    exp_33_ram[1668] = 19;
    exp_33_ram[1669] = 131;
    exp_33_ram[1670] = 3;
    exp_33_ram[1671] = 131;
    exp_33_ram[1672] = 3;
    exp_33_ram[1673] = 239;
    exp_33_ram[1674] = 35;
    exp_33_ram[1675] = 111;
    exp_33_ram[1676] = 131;
    exp_33_ram[1677] = 147;
    exp_33_ram[1678] = 99;
    exp_33_ram[1679] = 131;
    exp_33_ram[1680] = 147;
    exp_33_ram[1681] = 99;
    exp_33_ram[1682] = 131;
    exp_33_ram[1683] = 19;
    exp_33_ram[1684] = 35;
    exp_33_ram[1685] = 3;
    exp_33_ram[1686] = 131;
    exp_33_ram[1687] = 35;
    exp_33_ram[1688] = 131;
    exp_33_ram[1689] = 35;
    exp_33_ram[1690] = 131;
    exp_33_ram[1691] = 3;
    exp_33_ram[1692] = 147;
    exp_33_ram[1693] = 131;
    exp_33_ram[1694] = 3;
    exp_33_ram[1695] = 131;
    exp_33_ram[1696] = 3;
    exp_33_ram[1697] = 239;
    exp_33_ram[1698] = 35;
    exp_33_ram[1699] = 111;
    exp_33_ram[1700] = 131;
    exp_33_ram[1701] = 147;
    exp_33_ram[1702] = 99;
    exp_33_ram[1703] = 131;
    exp_33_ram[1704] = 19;
    exp_33_ram[1705] = 35;
    exp_33_ram[1706] = 131;
    exp_33_ram[1707] = 147;
    exp_33_ram[1708] = 111;
    exp_33_ram[1709] = 131;
    exp_33_ram[1710] = 147;
    exp_33_ram[1711] = 99;
    exp_33_ram[1712] = 131;
    exp_33_ram[1713] = 19;
    exp_33_ram[1714] = 35;
    exp_33_ram[1715] = 131;
    exp_33_ram[1716] = 147;
    exp_33_ram[1717] = 147;
    exp_33_ram[1718] = 111;
    exp_33_ram[1719] = 131;
    exp_33_ram[1720] = 19;
    exp_33_ram[1721] = 35;
    exp_33_ram[1722] = 131;
    exp_33_ram[1723] = 35;
    exp_33_ram[1724] = 131;
    exp_33_ram[1725] = 35;
    exp_33_ram[1726] = 131;
    exp_33_ram[1727] = 35;
    exp_33_ram[1728] = 131;
    exp_33_ram[1729] = 3;
    exp_33_ram[1730] = 147;
    exp_33_ram[1731] = 3;
    exp_33_ram[1732] = 131;
    exp_33_ram[1733] = 3;
    exp_33_ram[1734] = 131;
    exp_33_ram[1735] = 3;
    exp_33_ram[1736] = 239;
    exp_33_ram[1737] = 35;
    exp_33_ram[1738] = 131;
    exp_33_ram[1739] = 147;
    exp_33_ram[1740] = 35;
    exp_33_ram[1741] = 111;
    exp_33_ram[1742] = 147;
    exp_33_ram[1743] = 35;
    exp_33_ram[1744] = 131;
    exp_33_ram[1745] = 147;
    exp_33_ram[1746] = 99;
    exp_33_ram[1747] = 111;
    exp_33_ram[1748] = 131;
    exp_33_ram[1749] = 19;
    exp_33_ram[1750] = 35;
    exp_33_ram[1751] = 3;
    exp_33_ram[1752] = 131;
    exp_33_ram[1753] = 19;
    exp_33_ram[1754] = 131;
    exp_33_ram[1755] = 19;
    exp_33_ram[1756] = 231;
    exp_33_ram[1757] = 131;
    exp_33_ram[1758] = 19;
    exp_33_ram[1759] = 35;
    exp_33_ram[1760] = 3;
    exp_33_ram[1761] = 227;
    exp_33_ram[1762] = 131;
    exp_33_ram[1763] = 19;
    exp_33_ram[1764] = 35;
    exp_33_ram[1765] = 131;
    exp_33_ram[1766] = 19;
    exp_33_ram[1767] = 131;
    exp_33_ram[1768] = 19;
    exp_33_ram[1769] = 35;
    exp_33_ram[1770] = 3;
    exp_33_ram[1771] = 131;
    exp_33_ram[1772] = 19;
    exp_33_ram[1773] = 131;
    exp_33_ram[1774] = 231;
    exp_33_ram[1775] = 131;
    exp_33_ram[1776] = 147;
    exp_33_ram[1777] = 99;
    exp_33_ram[1778] = 111;
    exp_33_ram[1779] = 131;
    exp_33_ram[1780] = 19;
    exp_33_ram[1781] = 35;
    exp_33_ram[1782] = 3;
    exp_33_ram[1783] = 131;
    exp_33_ram[1784] = 19;
    exp_33_ram[1785] = 131;
    exp_33_ram[1786] = 19;
    exp_33_ram[1787] = 231;
    exp_33_ram[1788] = 131;
    exp_33_ram[1789] = 19;
    exp_33_ram[1790] = 35;
    exp_33_ram[1791] = 3;
    exp_33_ram[1792] = 227;
    exp_33_ram[1793] = 131;
    exp_33_ram[1794] = 147;
    exp_33_ram[1795] = 35;
    exp_33_ram[1796] = 111;
    exp_33_ram[1797] = 131;
    exp_33_ram[1798] = 19;
    exp_33_ram[1799] = 35;
    exp_33_ram[1800] = 131;
    exp_33_ram[1801] = 35;
    exp_33_ram[1802] = 131;
    exp_33_ram[1803] = 99;
    exp_33_ram[1804] = 131;
    exp_33_ram[1805] = 111;
    exp_33_ram[1806] = 147;
    exp_33_ram[1807] = 147;
    exp_33_ram[1808] = 3;
    exp_33_ram[1809] = 239;
    exp_33_ram[1810] = 35;
    exp_33_ram[1811] = 131;
    exp_33_ram[1812] = 147;
    exp_33_ram[1813] = 99;
    exp_33_ram[1814] = 3;
    exp_33_ram[1815] = 131;
    exp_33_ram[1816] = 99;
    exp_33_ram[1817] = 147;
    exp_33_ram[1818] = 35;
    exp_33_ram[1819] = 131;
    exp_33_ram[1820] = 147;
    exp_33_ram[1821] = 99;
    exp_33_ram[1822] = 111;
    exp_33_ram[1823] = 131;
    exp_33_ram[1824] = 19;
    exp_33_ram[1825] = 35;
    exp_33_ram[1826] = 3;
    exp_33_ram[1827] = 131;
    exp_33_ram[1828] = 19;
    exp_33_ram[1829] = 131;
    exp_33_ram[1830] = 19;
    exp_33_ram[1831] = 231;
    exp_33_ram[1832] = 131;
    exp_33_ram[1833] = 19;
    exp_33_ram[1834] = 35;
    exp_33_ram[1835] = 3;
    exp_33_ram[1836] = 227;
    exp_33_ram[1837] = 111;
    exp_33_ram[1838] = 131;
    exp_33_ram[1839] = 19;
    exp_33_ram[1840] = 35;
    exp_33_ram[1841] = 3;
    exp_33_ram[1842] = 131;
    exp_33_ram[1843] = 19;
    exp_33_ram[1844] = 35;
    exp_33_ram[1845] = 3;
    exp_33_ram[1846] = 131;
    exp_33_ram[1847] = 19;
    exp_33_ram[1848] = 131;
    exp_33_ram[1849] = 231;
    exp_33_ram[1850] = 131;
    exp_33_ram[1851] = 131;
    exp_33_ram[1852] = 99;
    exp_33_ram[1853] = 131;
    exp_33_ram[1854] = 147;
    exp_33_ram[1855] = 227;
    exp_33_ram[1856] = 131;
    exp_33_ram[1857] = 19;
    exp_33_ram[1858] = 35;
    exp_33_ram[1859] = 227;
    exp_33_ram[1860] = 131;
    exp_33_ram[1861] = 147;
    exp_33_ram[1862] = 99;
    exp_33_ram[1863] = 111;
    exp_33_ram[1864] = 131;
    exp_33_ram[1865] = 19;
    exp_33_ram[1866] = 35;
    exp_33_ram[1867] = 3;
    exp_33_ram[1868] = 131;
    exp_33_ram[1869] = 19;
    exp_33_ram[1870] = 131;
    exp_33_ram[1871] = 19;
    exp_33_ram[1872] = 231;
    exp_33_ram[1873] = 131;
    exp_33_ram[1874] = 19;
    exp_33_ram[1875] = 35;
    exp_33_ram[1876] = 3;
    exp_33_ram[1877] = 227;
    exp_33_ram[1878] = 131;
    exp_33_ram[1879] = 147;
    exp_33_ram[1880] = 35;
    exp_33_ram[1881] = 111;
    exp_33_ram[1882] = 147;
    exp_33_ram[1883] = 35;
    exp_33_ram[1884] = 131;
    exp_33_ram[1885] = 147;
    exp_33_ram[1886] = 35;
    exp_33_ram[1887] = 131;
    exp_33_ram[1888] = 19;
    exp_33_ram[1889] = 35;
    exp_33_ram[1890] = 131;
    exp_33_ram[1891] = 19;
    exp_33_ram[1892] = 131;
    exp_33_ram[1893] = 35;
    exp_33_ram[1894] = 131;
    exp_33_ram[1895] = 35;
    exp_33_ram[1896] = 131;
    exp_33_ram[1897] = 19;
    exp_33_ram[1898] = 147;
    exp_33_ram[1899] = 131;
    exp_33_ram[1900] = 3;
    exp_33_ram[1901] = 131;
    exp_33_ram[1902] = 3;
    exp_33_ram[1903] = 239;
    exp_33_ram[1904] = 35;
    exp_33_ram[1905] = 131;
    exp_33_ram[1906] = 147;
    exp_33_ram[1907] = 35;
    exp_33_ram[1908] = 111;
    exp_33_ram[1909] = 131;
    exp_33_ram[1910] = 19;
    exp_33_ram[1911] = 35;
    exp_33_ram[1912] = 3;
    exp_33_ram[1913] = 131;
    exp_33_ram[1914] = 19;
    exp_33_ram[1915] = 131;
    exp_33_ram[1916] = 19;
    exp_33_ram[1917] = 231;
    exp_33_ram[1918] = 131;
    exp_33_ram[1919] = 147;
    exp_33_ram[1920] = 35;
    exp_33_ram[1921] = 111;
    exp_33_ram[1922] = 131;
    exp_33_ram[1923] = 3;
    exp_33_ram[1924] = 131;
    exp_33_ram[1925] = 19;
    exp_33_ram[1926] = 35;
    exp_33_ram[1927] = 3;
    exp_33_ram[1928] = 131;
    exp_33_ram[1929] = 19;
    exp_33_ram[1930] = 131;
    exp_33_ram[1931] = 231;
    exp_33_ram[1932] = 131;
    exp_33_ram[1933] = 147;
    exp_33_ram[1934] = 35;
    exp_33_ram[1935] = 19;
    exp_33_ram[1936] = 131;
    exp_33_ram[1937] = 131;
    exp_33_ram[1938] = 99;
    exp_33_ram[1939] = 3;
    exp_33_ram[1940] = 131;
    exp_33_ram[1941] = 99;
    exp_33_ram[1942] = 131;
    exp_33_ram[1943] = 147;
    exp_33_ram[1944] = 111;
    exp_33_ram[1945] = 131;
    exp_33_ram[1946] = 3;
    exp_33_ram[1947] = 131;
    exp_33_ram[1948] = 19;
    exp_33_ram[1949] = 131;
    exp_33_ram[1950] = 19;
    exp_33_ram[1951] = 231;
    exp_33_ram[1952] = 131;
    exp_33_ram[1953] = 19;
    exp_33_ram[1954] = 131;
    exp_33_ram[1955] = 3;
    exp_33_ram[1956] = 19;
    exp_33_ram[1957] = 103;
    exp_33_ram[1958] = 19;
    exp_33_ram[1959] = 35;
    exp_33_ram[1960] = 35;
    exp_33_ram[1961] = 19;
    exp_33_ram[1962] = 35;
    exp_33_ram[1963] = 35;
    exp_33_ram[1964] = 35;
    exp_33_ram[1965] = 35;
    exp_33_ram[1966] = 35;
    exp_33_ram[1967] = 35;
    exp_33_ram[1968] = 35;
    exp_33_ram[1969] = 35;
    exp_33_ram[1970] = 147;
    exp_33_ram[1971] = 35;
    exp_33_ram[1972] = 131;
    exp_33_ram[1973] = 147;
    exp_33_ram[1974] = 35;
    exp_33_ram[1975] = 3;
    exp_33_ram[1976] = 147;
    exp_33_ram[1977] = 131;
    exp_33_ram[1978] = 19;
    exp_33_ram[1979] = 147;
    exp_33_ram[1980] = 183;
    exp_33_ram[1981] = 19;
    exp_33_ram[1982] = 239;
    exp_33_ram[1983] = 35;
    exp_33_ram[1984] = 131;
    exp_33_ram[1985] = 19;
    exp_33_ram[1986] = 131;
    exp_33_ram[1987] = 3;
    exp_33_ram[1988] = 19;
    exp_33_ram[1989] = 103;
    exp_33_ram[1990] = 19;
    exp_33_ram[1991] = 35;
    exp_33_ram[1992] = 35;
    exp_33_ram[1993] = 19;
    exp_33_ram[1994] = 147;
    exp_33_ram[1995] = 163;
    exp_33_ram[1996] = 3;
    exp_33_ram[1997] = 183;
    exp_33_ram[1998] = 131;
    exp_33_ram[1999] = 147;
    exp_33_ram[2000] = 19;
    exp_33_ram[2001] = 239;
    exp_33_ram[2002] = 19;
    exp_33_ram[2003] = 131;
    exp_33_ram[2004] = 3;
    exp_33_ram[2005] = 19;
    exp_33_ram[2006] = 103;
    exp_33_ram[2007] = 19;
    exp_33_ram[2008] = 35;
    exp_33_ram[2009] = 35;
    exp_33_ram[2010] = 35;
    exp_33_ram[2011] = 19;
    exp_33_ram[2012] = 147;
    exp_33_ram[2013] = 131;
    exp_33_ram[2014] = 35;
    exp_33_ram[2015] = 147;
    exp_33_ram[2016] = 35;
    exp_33_ram[2017] = 147;
    exp_33_ram[2018] = 35;
    exp_33_ram[2019] = 147;
    exp_33_ram[2020] = 35;
    exp_33_ram[2021] = 35;
    exp_33_ram[2022] = 35;
    exp_33_ram[2023] = 35;
    exp_33_ram[2024] = 3;
    exp_33_ram[2025] = 131;
    exp_33_ram[2026] = 3;
    exp_33_ram[2027] = 3;
    exp_33_ram[2028] = 131;
    exp_33_ram[2029] = 3;
    exp_33_ram[2030] = 131;
    exp_33_ram[2031] = 3;
    exp_33_ram[2032] = 131;
    exp_33_ram[2033] = 35;
    exp_33_ram[2034] = 35;
    exp_33_ram[2035] = 35;
    exp_33_ram[2036] = 35;
    exp_33_ram[2037] = 35;
    exp_33_ram[2038] = 35;
    exp_33_ram[2039] = 35;
    exp_33_ram[2040] = 35;
    exp_33_ram[2041] = 35;
    exp_33_ram[2042] = 147;
    exp_33_ram[2043] = 19;
    exp_33_ram[2044] = 239;
    exp_33_ram[2045] = 35;
    exp_33_ram[2046] = 35;
    exp_33_ram[2047] = 147;
    exp_33_ram[2048] = 131;
    exp_33_ram[2049] = 3;
    exp_33_ram[2050] = 19;
    exp_33_ram[2051] = 239;
    exp_33_ram[2052] = 3;
    exp_33_ram[2053] = 131;
    exp_33_ram[2054] = 179;
    exp_33_ram[2055] = 35;
    exp_33_ram[2056] = 3;
    exp_33_ram[2057] = 131;
    exp_33_ram[2058] = 3;
    exp_33_ram[2059] = 3;
    exp_33_ram[2060] = 131;
    exp_33_ram[2061] = 3;
    exp_33_ram[2062] = 131;
    exp_33_ram[2063] = 3;
    exp_33_ram[2064] = 131;
    exp_33_ram[2065] = 35;
    exp_33_ram[2066] = 35;
    exp_33_ram[2067] = 35;
    exp_33_ram[2068] = 35;
    exp_33_ram[2069] = 35;
    exp_33_ram[2070] = 35;
    exp_33_ram[2071] = 35;
    exp_33_ram[2072] = 35;
    exp_33_ram[2073] = 35;
    exp_33_ram[2074] = 147;
    exp_33_ram[2075] = 19;
    exp_33_ram[2076] = 239;
    exp_33_ram[2077] = 35;
    exp_33_ram[2078] = 35;
    exp_33_ram[2079] = 131;
    exp_33_ram[2080] = 35;
    exp_33_ram[2081] = 147;
    exp_33_ram[2082] = 35;
    exp_33_ram[2083] = 147;
    exp_33_ram[2084] = 35;
    exp_33_ram[2085] = 147;
    exp_33_ram[2086] = 35;
    exp_33_ram[2087] = 35;
    exp_33_ram[2088] = 35;
    exp_33_ram[2089] = 35;
    exp_33_ram[2090] = 3;
    exp_33_ram[2091] = 131;
    exp_33_ram[2092] = 3;
    exp_33_ram[2093] = 3;
    exp_33_ram[2094] = 131;
    exp_33_ram[2095] = 3;
    exp_33_ram[2096] = 131;
    exp_33_ram[2097] = 3;
    exp_33_ram[2098] = 131;
    exp_33_ram[2099] = 35;
    exp_33_ram[2100] = 35;
    exp_33_ram[2101] = 35;
    exp_33_ram[2102] = 35;
    exp_33_ram[2103] = 35;
    exp_33_ram[2104] = 35;
    exp_33_ram[2105] = 35;
    exp_33_ram[2106] = 35;
    exp_33_ram[2107] = 35;
    exp_33_ram[2108] = 147;
    exp_33_ram[2109] = 19;
    exp_33_ram[2110] = 239;
    exp_33_ram[2111] = 35;
    exp_33_ram[2112] = 35;
    exp_33_ram[2113] = 147;
    exp_33_ram[2114] = 131;
    exp_33_ram[2115] = 3;
    exp_33_ram[2116] = 19;
    exp_33_ram[2117] = 239;
    exp_33_ram[2118] = 3;
    exp_33_ram[2119] = 131;
    exp_33_ram[2120] = 179;
    exp_33_ram[2121] = 35;
    exp_33_ram[2122] = 3;
    exp_33_ram[2123] = 131;
    exp_33_ram[2124] = 3;
    exp_33_ram[2125] = 3;
    exp_33_ram[2126] = 131;
    exp_33_ram[2127] = 3;
    exp_33_ram[2128] = 131;
    exp_33_ram[2129] = 3;
    exp_33_ram[2130] = 131;
    exp_33_ram[2131] = 35;
    exp_33_ram[2132] = 35;
    exp_33_ram[2133] = 35;
    exp_33_ram[2134] = 35;
    exp_33_ram[2135] = 35;
    exp_33_ram[2136] = 35;
    exp_33_ram[2137] = 35;
    exp_33_ram[2138] = 35;
    exp_33_ram[2139] = 35;
    exp_33_ram[2140] = 147;
    exp_33_ram[2141] = 19;
    exp_33_ram[2142] = 239;
    exp_33_ram[2143] = 35;
    exp_33_ram[2144] = 35;
    exp_33_ram[2145] = 3;
    exp_33_ram[2146] = 131;
    exp_33_ram[2147] = 3;
    exp_33_ram[2148] = 3;
    exp_33_ram[2149] = 131;
    exp_33_ram[2150] = 3;
    exp_33_ram[2151] = 131;
    exp_33_ram[2152] = 3;
    exp_33_ram[2153] = 131;
    exp_33_ram[2154] = 35;
    exp_33_ram[2155] = 35;
    exp_33_ram[2156] = 35;
    exp_33_ram[2157] = 35;
    exp_33_ram[2158] = 35;
    exp_33_ram[2159] = 35;
    exp_33_ram[2160] = 35;
    exp_33_ram[2161] = 35;
    exp_33_ram[2162] = 35;
    exp_33_ram[2163] = 147;
    exp_33_ram[2164] = 19;
    exp_33_ram[2165] = 239;
    exp_33_ram[2166] = 35;
    exp_33_ram[2167] = 35;
    exp_33_ram[2168] = 3;
    exp_33_ram[2169] = 131;
    exp_33_ram[2170] = 99;
    exp_33_ram[2171] = 3;
    exp_33_ram[2172] = 131;
    exp_33_ram[2173] = 99;
    exp_33_ram[2174] = 3;
    exp_33_ram[2175] = 131;
    exp_33_ram[2176] = 99;
    exp_33_ram[2177] = 3;
    exp_33_ram[2178] = 131;
    exp_33_ram[2179] = 99;
    exp_33_ram[2180] = 3;
    exp_33_ram[2181] = 131;
    exp_33_ram[2182] = 99;
    exp_33_ram[2183] = 3;
    exp_33_ram[2184] = 131;
    exp_33_ram[2185] = 99;
    exp_33_ram[2186] = 147;
    exp_33_ram[2187] = 111;
    exp_33_ram[2188] = 147;
    exp_33_ram[2189] = 19;
    exp_33_ram[2190] = 131;
    exp_33_ram[2191] = 3;
    exp_33_ram[2192] = 131;
    exp_33_ram[2193] = 19;
    exp_33_ram[2194] = 103;
    exp_33_ram[2195] = 19;
    exp_33_ram[2196] = 35;
    exp_33_ram[2197] = 35;
    exp_33_ram[2198] = 19;
    exp_33_ram[2199] = 35;
    exp_33_ram[2200] = 35;
    exp_33_ram[2201] = 147;
    exp_33_ram[2202] = 131;
    exp_33_ram[2203] = 3;
    exp_33_ram[2204] = 19;
    exp_33_ram[2205] = 239;
    exp_33_ram[2206] = 3;
    exp_33_ram[2207] = 131;
    exp_33_ram[2208] = 3;
    exp_33_ram[2209] = 3;
    exp_33_ram[2210] = 131;
    exp_33_ram[2211] = 3;
    exp_33_ram[2212] = 131;
    exp_33_ram[2213] = 3;
    exp_33_ram[2214] = 131;
    exp_33_ram[2215] = 35;
    exp_33_ram[2216] = 35;
    exp_33_ram[2217] = 35;
    exp_33_ram[2218] = 35;
    exp_33_ram[2219] = 35;
    exp_33_ram[2220] = 35;
    exp_33_ram[2221] = 35;
    exp_33_ram[2222] = 35;
    exp_33_ram[2223] = 35;
    exp_33_ram[2224] = 147;
    exp_33_ram[2225] = 19;
    exp_33_ram[2226] = 239;
    exp_33_ram[2227] = 147;
    exp_33_ram[2228] = 19;
    exp_33_ram[2229] = 131;
    exp_33_ram[2230] = 3;
    exp_33_ram[2231] = 19;
    exp_33_ram[2232] = 103;
    exp_33_ram[2233] = 19;
    exp_33_ram[2234] = 35;
    exp_33_ram[2235] = 19;
    exp_33_ram[2236] = 183;
    exp_33_ram[2237] = 35;
    exp_33_ram[2238] = 183;
    exp_33_ram[2239] = 147;
    exp_33_ram[2240] = 35;
    exp_33_ram[2241] = 131;
    exp_33_ram[2242] = 3;
    exp_33_ram[2243] = 131;
    exp_33_ram[2244] = 3;
    exp_33_ram[2245] = 131;
    exp_33_ram[2246] = 3;
    exp_33_ram[2247] = 147;
    exp_33_ram[2248] = 19;
    exp_33_ram[2249] = 51;
    exp_33_ram[2250] = 179;
    exp_33_ram[2251] = 19;
    exp_33_ram[2252] = 147;
    exp_33_ram[2253] = 19;
    exp_33_ram[2254] = 147;
    exp_33_ram[2255] = 3;
    exp_33_ram[2256] = 19;
    exp_33_ram[2257] = 103;
    exp_33_ram[2258] = 19;
    exp_33_ram[2259] = 35;
    exp_33_ram[2260] = 35;
    exp_33_ram[2261] = 19;
    exp_33_ram[2262] = 35;
    exp_33_ram[2263] = 35;
    exp_33_ram[2264] = 35;
    exp_33_ram[2265] = 35;
    exp_33_ram[2266] = 3;
    exp_33_ram[2267] = 131;
    exp_33_ram[2268] = 3;
    exp_33_ram[2269] = 131;
    exp_33_ram[2270] = 51;
    exp_33_ram[2271] = 19;
    exp_33_ram[2272] = 51;
    exp_33_ram[2273] = 179;
    exp_33_ram[2274] = 179;
    exp_33_ram[2275] = 147;
    exp_33_ram[2276] = 19;
    exp_33_ram[2277] = 147;
    exp_33_ram[2278] = 19;
    exp_33_ram[2279] = 147;
    exp_33_ram[2280] = 239;
    exp_33_ram[2281] = 19;
    exp_33_ram[2282] = 147;
    exp_33_ram[2283] = 19;
    exp_33_ram[2284] = 147;
    exp_33_ram[2285] = 131;
    exp_33_ram[2286] = 3;
    exp_33_ram[2287] = 19;
    exp_33_ram[2288] = 103;
    exp_33_ram[2289] = 19;
    exp_33_ram[2290] = 35;
    exp_33_ram[2291] = 19;
    exp_33_ram[2292] = 35;
    exp_33_ram[2293] = 131;
    exp_33_ram[2294] = 147;
    exp_33_ram[2295] = 99;
    exp_33_ram[2296] = 3;
    exp_33_ram[2297] = 147;
    exp_33_ram[2298] = 179;
    exp_33_ram[2299] = 99;
    exp_33_ram[2300] = 3;
    exp_33_ram[2301] = 147;
    exp_33_ram[2302] = 179;
    exp_33_ram[2303] = 99;
    exp_33_ram[2304] = 147;
    exp_33_ram[2305] = 111;
    exp_33_ram[2306] = 147;
    exp_33_ram[2307] = 19;
    exp_33_ram[2308] = 3;
    exp_33_ram[2309] = 19;
    exp_33_ram[2310] = 103;
    exp_33_ram[2311] = 19;
    exp_33_ram[2312] = 35;
    exp_33_ram[2313] = 35;
    exp_33_ram[2314] = 19;
    exp_33_ram[2315] = 35;
    exp_33_ram[2316] = 3;
    exp_33_ram[2317] = 239;
    exp_33_ram[2318] = 147;
    exp_33_ram[2319] = 99;
    exp_33_ram[2320] = 147;
    exp_33_ram[2321] = 111;
    exp_33_ram[2322] = 147;
    exp_33_ram[2323] = 19;
    exp_33_ram[2324] = 131;
    exp_33_ram[2325] = 3;
    exp_33_ram[2326] = 19;
    exp_33_ram[2327] = 103;
    exp_33_ram[2328] = 19;
    exp_33_ram[2329] = 35;
    exp_33_ram[2330] = 35;
    exp_33_ram[2331] = 19;
    exp_33_ram[2332] = 35;
    exp_33_ram[2333] = 35;
    exp_33_ram[2334] = 3;
    exp_33_ram[2335] = 147;
    exp_33_ram[2336] = 99;
    exp_33_ram[2337] = 3;
    exp_33_ram[2338] = 147;
    exp_33_ram[2339] = 99;
    exp_33_ram[2340] = 3;
    exp_33_ram[2341] = 147;
    exp_33_ram[2342] = 99;
    exp_33_ram[2343] = 3;
    exp_33_ram[2344] = 147;
    exp_33_ram[2345] = 99;
    exp_33_ram[2346] = 147;
    exp_33_ram[2347] = 111;
    exp_33_ram[2348] = 3;
    exp_33_ram[2349] = 147;
    exp_33_ram[2350] = 99;
    exp_33_ram[2351] = 3;
    exp_33_ram[2352] = 239;
    exp_33_ram[2353] = 147;
    exp_33_ram[2354] = 99;
    exp_33_ram[2355] = 147;
    exp_33_ram[2356] = 111;
    exp_33_ram[2357] = 147;
    exp_33_ram[2358] = 111;
    exp_33_ram[2359] = 147;
    exp_33_ram[2360] = 19;
    exp_33_ram[2361] = 131;
    exp_33_ram[2362] = 3;
    exp_33_ram[2363] = 19;
    exp_33_ram[2364] = 103;
    exp_33_ram[2365] = 19;
    exp_33_ram[2366] = 35;
    exp_33_ram[2367] = 35;
    exp_33_ram[2368] = 35;
    exp_33_ram[2369] = 35;
    exp_33_ram[2370] = 35;
    exp_33_ram[2371] = 35;
    exp_33_ram[2372] = 35;
    exp_33_ram[2373] = 35;
    exp_33_ram[2374] = 35;
    exp_33_ram[2375] = 35;
    exp_33_ram[2376] = 35;
    exp_33_ram[2377] = 35;
    exp_33_ram[2378] = 35;
    exp_33_ram[2379] = 19;
    exp_33_ram[2380] = 147;
    exp_33_ram[2381] = 147;
    exp_33_ram[2382] = 19;
    exp_33_ram[2383] = 35;
    exp_33_ram[2384] = 35;
    exp_33_ram[2385] = 147;
    exp_33_ram[2386] = 35;
    exp_33_ram[2387] = 131;
    exp_33_ram[2388] = 35;
    exp_33_ram[2389] = 131;
    exp_33_ram[2390] = 147;
    exp_33_ram[2391] = 3;
    exp_33_ram[2392] = 99;
    exp_33_ram[2393] = 3;
    exp_33_ram[2394] = 239;
    exp_33_ram[2395] = 19;
    exp_33_ram[2396] = 183;
    exp_33_ram[2397] = 147;
    exp_33_ram[2398] = 179;
    exp_33_ram[2399] = 35;
    exp_33_ram[2400] = 35;
    exp_33_ram[2401] = 3;
    exp_33_ram[2402] = 131;
    exp_33_ram[2403] = 3;
    exp_33_ram[2404] = 131;
    exp_33_ram[2405] = 147;
    exp_33_ram[2406] = 51;
    exp_33_ram[2407] = 147;
    exp_33_ram[2408] = 179;
    exp_33_ram[2409] = 19;
    exp_33_ram[2410] = 179;
    exp_33_ram[2411] = 179;
    exp_33_ram[2412] = 147;
    exp_33_ram[2413] = 35;
    exp_33_ram[2414] = 35;
    exp_33_ram[2415] = 131;
    exp_33_ram[2416] = 147;
    exp_33_ram[2417] = 35;
    exp_33_ram[2418] = 111;
    exp_33_ram[2419] = 19;
    exp_33_ram[2420] = 35;
    exp_33_ram[2421] = 131;
    exp_33_ram[2422] = 19;
    exp_33_ram[2423] = 131;
    exp_33_ram[2424] = 99;
    exp_33_ram[2425] = 131;
    exp_33_ram[2426] = 3;
    exp_33_ram[2427] = 239;
    exp_33_ram[2428] = 19;
    exp_33_ram[2429] = 183;
    exp_33_ram[2430] = 147;
    exp_33_ram[2431] = 179;
    exp_33_ram[2432] = 19;
    exp_33_ram[2433] = 147;
    exp_33_ram[2434] = 3;
    exp_33_ram[2435] = 131;
    exp_33_ram[2436] = 51;
    exp_33_ram[2437] = 147;
    exp_33_ram[2438] = 179;
    exp_33_ram[2439] = 179;
    exp_33_ram[2440] = 179;
    exp_33_ram[2441] = 147;
    exp_33_ram[2442] = 35;
    exp_33_ram[2443] = 35;
    exp_33_ram[2444] = 131;
    exp_33_ram[2445] = 147;
    exp_33_ram[2446] = 35;
    exp_33_ram[2447] = 111;
    exp_33_ram[2448] = 19;
    exp_33_ram[2449] = 131;
    exp_33_ram[2450] = 19;
    exp_33_ram[2451] = 183;
    exp_33_ram[2452] = 147;
    exp_33_ram[2453] = 179;
    exp_33_ram[2454] = 19;
    exp_33_ram[2455] = 147;
    exp_33_ram[2456] = 147;
    exp_33_ram[2457] = 3;
    exp_33_ram[2458] = 131;
    exp_33_ram[2459] = 51;
    exp_33_ram[2460] = 147;
    exp_33_ram[2461] = 179;
    exp_33_ram[2462] = 179;
    exp_33_ram[2463] = 179;
    exp_33_ram[2464] = 147;
    exp_33_ram[2465] = 35;
    exp_33_ram[2466] = 35;
    exp_33_ram[2467] = 3;
    exp_33_ram[2468] = 183;
    exp_33_ram[2469] = 147;
    exp_33_ram[2470] = 179;
    exp_33_ram[2471] = 19;
    exp_33_ram[2472] = 147;
    exp_33_ram[2473] = 147;
    exp_33_ram[2474] = 3;
    exp_33_ram[2475] = 131;
    exp_33_ram[2476] = 51;
    exp_33_ram[2477] = 147;
    exp_33_ram[2478] = 179;
    exp_33_ram[2479] = 179;
    exp_33_ram[2480] = 179;
    exp_33_ram[2481] = 147;
    exp_33_ram[2482] = 35;
    exp_33_ram[2483] = 35;
    exp_33_ram[2484] = 3;
    exp_33_ram[2485] = 147;
    exp_33_ram[2486] = 147;
    exp_33_ram[2487] = 179;
    exp_33_ram[2488] = 147;
    exp_33_ram[2489] = 19;
    exp_33_ram[2490] = 147;
    exp_33_ram[2491] = 147;
    exp_33_ram[2492] = 3;
    exp_33_ram[2493] = 131;
    exp_33_ram[2494] = 51;
    exp_33_ram[2495] = 147;
    exp_33_ram[2496] = 179;
    exp_33_ram[2497] = 179;
    exp_33_ram[2498] = 179;
    exp_33_ram[2499] = 147;
    exp_33_ram[2500] = 35;
    exp_33_ram[2501] = 35;
    exp_33_ram[2502] = 131;
    exp_33_ram[2503] = 19;
    exp_33_ram[2504] = 147;
    exp_33_ram[2505] = 147;
    exp_33_ram[2506] = 3;
    exp_33_ram[2507] = 131;
    exp_33_ram[2508] = 51;
    exp_33_ram[2509] = 147;
    exp_33_ram[2510] = 179;
    exp_33_ram[2511] = 179;
    exp_33_ram[2512] = 179;
    exp_33_ram[2513] = 147;
    exp_33_ram[2514] = 35;
    exp_33_ram[2515] = 35;
    exp_33_ram[2516] = 3;
    exp_33_ram[2517] = 131;
    exp_33_ram[2518] = 19;
    exp_33_ram[2519] = 147;
    exp_33_ram[2520] = 131;
    exp_33_ram[2521] = 3;
    exp_33_ram[2522] = 131;
    exp_33_ram[2523] = 3;
    exp_33_ram[2524] = 131;
    exp_33_ram[2525] = 3;
    exp_33_ram[2526] = 131;
    exp_33_ram[2527] = 3;
    exp_33_ram[2528] = 131;
    exp_33_ram[2529] = 3;
    exp_33_ram[2530] = 131;
    exp_33_ram[2531] = 3;
    exp_33_ram[2532] = 131;
    exp_33_ram[2533] = 19;
    exp_33_ram[2534] = 103;
    exp_33_ram[2535] = 19;
    exp_33_ram[2536] = 35;
    exp_33_ram[2537] = 35;
    exp_33_ram[2538] = 35;
    exp_33_ram[2539] = 35;
    exp_33_ram[2540] = 35;
    exp_33_ram[2541] = 19;
    exp_33_ram[2542] = 35;
    exp_33_ram[2543] = 131;
    exp_33_ram[2544] = 3;
    exp_33_ram[2545] = 131;
    exp_33_ram[2546] = 3;
    exp_33_ram[2547] = 3;
    exp_33_ram[2548] = 131;
    exp_33_ram[2549] = 3;
    exp_33_ram[2550] = 131;
    exp_33_ram[2551] = 3;
    exp_33_ram[2552] = 131;
    exp_33_ram[2553] = 35;
    exp_33_ram[2554] = 35;
    exp_33_ram[2555] = 35;
    exp_33_ram[2556] = 35;
    exp_33_ram[2557] = 35;
    exp_33_ram[2558] = 35;
    exp_33_ram[2559] = 35;
    exp_33_ram[2560] = 35;
    exp_33_ram[2561] = 35;
    exp_33_ram[2562] = 3;
    exp_33_ram[2563] = 131;
    exp_33_ram[2564] = 3;
    exp_33_ram[2565] = 3;
    exp_33_ram[2566] = 131;
    exp_33_ram[2567] = 3;
    exp_33_ram[2568] = 131;
    exp_33_ram[2569] = 3;
    exp_33_ram[2570] = 131;
    exp_33_ram[2571] = 35;
    exp_33_ram[2572] = 35;
    exp_33_ram[2573] = 35;
    exp_33_ram[2574] = 35;
    exp_33_ram[2575] = 35;
    exp_33_ram[2576] = 35;
    exp_33_ram[2577] = 35;
    exp_33_ram[2578] = 35;
    exp_33_ram[2579] = 35;
    exp_33_ram[2580] = 147;
    exp_33_ram[2581] = 19;
    exp_33_ram[2582] = 239;
    exp_33_ram[2583] = 35;
    exp_33_ram[2584] = 35;
    exp_33_ram[2585] = 131;
    exp_33_ram[2586] = 99;
    exp_33_ram[2587] = 3;
    exp_33_ram[2588] = 131;
    exp_33_ram[2589] = 55;
    exp_33_ram[2590] = 19;
    exp_33_ram[2591] = 147;
    exp_33_ram[2592] = 51;
    exp_33_ram[2593] = 19;
    exp_33_ram[2594] = 51;
    exp_33_ram[2595] = 179;
    exp_33_ram[2596] = 179;
    exp_33_ram[2597] = 147;
    exp_33_ram[2598] = 35;
    exp_33_ram[2599] = 35;
    exp_33_ram[2600] = 111;
    exp_33_ram[2601] = 131;
    exp_33_ram[2602] = 99;
    exp_33_ram[2603] = 3;
    exp_33_ram[2604] = 131;
    exp_33_ram[2605] = 3;
    exp_33_ram[2606] = 3;
    exp_33_ram[2607] = 131;
    exp_33_ram[2608] = 3;
    exp_33_ram[2609] = 131;
    exp_33_ram[2610] = 3;
    exp_33_ram[2611] = 131;
    exp_33_ram[2612] = 35;
    exp_33_ram[2613] = 35;
    exp_33_ram[2614] = 35;
    exp_33_ram[2615] = 35;
    exp_33_ram[2616] = 35;
    exp_33_ram[2617] = 35;
    exp_33_ram[2618] = 35;
    exp_33_ram[2619] = 35;
    exp_33_ram[2620] = 35;
    exp_33_ram[2621] = 147;
    exp_33_ram[2622] = 19;
    exp_33_ram[2623] = 239;
    exp_33_ram[2624] = 147;
    exp_33_ram[2625] = 99;
    exp_33_ram[2626] = 55;
    exp_33_ram[2627] = 19;
    exp_33_ram[2628] = 147;
    exp_33_ram[2629] = 111;
    exp_33_ram[2630] = 19;
    exp_33_ram[2631] = 147;
    exp_33_ram[2632] = 3;
    exp_33_ram[2633] = 131;
    exp_33_ram[2634] = 51;
    exp_33_ram[2635] = 19;
    exp_33_ram[2636] = 51;
    exp_33_ram[2637] = 179;
    exp_33_ram[2638] = 179;
    exp_33_ram[2639] = 147;
    exp_33_ram[2640] = 35;
    exp_33_ram[2641] = 35;
    exp_33_ram[2642] = 111;
    exp_33_ram[2643] = 3;
    exp_33_ram[2644] = 131;
    exp_33_ram[2645] = 35;
    exp_33_ram[2646] = 35;
    exp_33_ram[2647] = 183;
    exp_33_ram[2648] = 131;
    exp_33_ram[2649] = 19;
    exp_33_ram[2650] = 147;
    exp_33_ram[2651] = 147;
    exp_33_ram[2652] = 3;
    exp_33_ram[2653] = 131;
    exp_33_ram[2654] = 51;
    exp_33_ram[2655] = 147;
    exp_33_ram[2656] = 179;
    exp_33_ram[2657] = 179;
    exp_33_ram[2658] = 179;
    exp_33_ram[2659] = 147;
    exp_33_ram[2660] = 35;
    exp_33_ram[2661] = 35;
    exp_33_ram[2662] = 131;
    exp_33_ram[2663] = 147;
    exp_33_ram[2664] = 131;
    exp_33_ram[2665] = 3;
    exp_33_ram[2666] = 19;
    exp_33_ram[2667] = 239;
    exp_33_ram[2668] = 3;
    exp_33_ram[2669] = 131;
    exp_33_ram[2670] = 3;
    exp_33_ram[2671] = 3;
    exp_33_ram[2672] = 131;
    exp_33_ram[2673] = 3;
    exp_33_ram[2674] = 131;
    exp_33_ram[2675] = 3;
    exp_33_ram[2676] = 131;
    exp_33_ram[2677] = 35;
    exp_33_ram[2678] = 35;
    exp_33_ram[2679] = 35;
    exp_33_ram[2680] = 35;
    exp_33_ram[2681] = 35;
    exp_33_ram[2682] = 35;
    exp_33_ram[2683] = 35;
    exp_33_ram[2684] = 35;
    exp_33_ram[2685] = 35;
    exp_33_ram[2686] = 131;
    exp_33_ram[2687] = 99;
    exp_33_ram[2688] = 131;
    exp_33_ram[2689] = 19;
    exp_33_ram[2690] = 35;
    exp_33_ram[2691] = 111;
    exp_33_ram[2692] = 131;
    exp_33_ram[2693] = 99;
    exp_33_ram[2694] = 3;
    exp_33_ram[2695] = 131;
    exp_33_ram[2696] = 3;
    exp_33_ram[2697] = 3;
    exp_33_ram[2698] = 131;
    exp_33_ram[2699] = 3;
    exp_33_ram[2700] = 131;
    exp_33_ram[2701] = 3;
    exp_33_ram[2702] = 131;
    exp_33_ram[2703] = 35;
    exp_33_ram[2704] = 35;
    exp_33_ram[2705] = 35;
    exp_33_ram[2706] = 35;
    exp_33_ram[2707] = 35;
    exp_33_ram[2708] = 35;
    exp_33_ram[2709] = 35;
    exp_33_ram[2710] = 35;
    exp_33_ram[2711] = 35;
    exp_33_ram[2712] = 147;
    exp_33_ram[2713] = 19;
    exp_33_ram[2714] = 239;
    exp_33_ram[2715] = 19;
    exp_33_ram[2716] = 131;
    exp_33_ram[2717] = 35;
    exp_33_ram[2718] = 111;
    exp_33_ram[2719] = 131;
    exp_33_ram[2720] = 35;
    exp_33_ram[2721] = 3;
    exp_33_ram[2722] = 131;
    exp_33_ram[2723] = 19;
    exp_33_ram[2724] = 147;
    exp_33_ram[2725] = 131;
    exp_33_ram[2726] = 3;
    exp_33_ram[2727] = 131;
    exp_33_ram[2728] = 3;
    exp_33_ram[2729] = 131;
    exp_33_ram[2730] = 19;
    exp_33_ram[2731] = 103;
    exp_33_ram[2732] = 19;
    exp_33_ram[2733] = 35;
    exp_33_ram[2734] = 35;
    exp_33_ram[2735] = 35;
    exp_33_ram[2736] = 35;
    exp_33_ram[2737] = 35;
    exp_33_ram[2738] = 35;
    exp_33_ram[2739] = 35;
    exp_33_ram[2740] = 35;
    exp_33_ram[2741] = 19;
    exp_33_ram[2742] = 35;
    exp_33_ram[2743] = 239;
    exp_33_ram[2744] = 19;
    exp_33_ram[2745] = 147;
    exp_33_ram[2746] = 183;
    exp_33_ram[2747] = 131;
    exp_33_ram[2748] = 19;
    exp_33_ram[2749] = 147;
    exp_33_ram[2750] = 19;
    exp_33_ram[2751] = 147;
    exp_33_ram[2752] = 19;
    exp_33_ram[2753] = 147;
    exp_33_ram[2754] = 239;
    exp_33_ram[2755] = 19;
    exp_33_ram[2756] = 147;
    exp_33_ram[2757] = 35;
    exp_33_ram[2758] = 183;
    exp_33_ram[2759] = 3;
    exp_33_ram[2760] = 131;
    exp_33_ram[2761] = 131;
    exp_33_ram[2762] = 179;
    exp_33_ram[2763] = 35;
    exp_33_ram[2764] = 131;
    exp_33_ram[2765] = 99;
    exp_33_ram[2766] = 131;
    exp_33_ram[2767] = 19;
    exp_33_ram[2768] = 147;
    exp_33_ram[2769] = 131;
    exp_33_ram[2770] = 35;
    exp_33_ram[2771] = 35;
    exp_33_ram[2772] = 131;
    exp_33_ram[2773] = 19;
    exp_33_ram[2774] = 147;
    exp_33_ram[2775] = 19;
    exp_33_ram[2776] = 147;
    exp_33_ram[2777] = 19;
    exp_33_ram[2778] = 147;
    exp_33_ram[2779] = 131;
    exp_33_ram[2780] = 3;
    exp_33_ram[2781] = 3;
    exp_33_ram[2782] = 131;
    exp_33_ram[2783] = 3;
    exp_33_ram[2784] = 131;
    exp_33_ram[2785] = 3;
    exp_33_ram[2786] = 131;
    exp_33_ram[2787] = 19;
    exp_33_ram[2788] = 103;
    exp_33_ram[2789] = 19;
    exp_33_ram[2790] = 35;
    exp_33_ram[2791] = 35;
    exp_33_ram[2792] = 35;
    exp_33_ram[2793] = 35;
    exp_33_ram[2794] = 19;
    exp_33_ram[2795] = 35;
    exp_33_ram[2796] = 35;
    exp_33_ram[2797] = 239;
    exp_33_ram[2798] = 19;
    exp_33_ram[2799] = 147;
    exp_33_ram[2800] = 183;
    exp_33_ram[2801] = 131;
    exp_33_ram[2802] = 19;
    exp_33_ram[2803] = 147;
    exp_33_ram[2804] = 19;
    exp_33_ram[2805] = 147;
    exp_33_ram[2806] = 19;
    exp_33_ram[2807] = 147;
    exp_33_ram[2808] = 239;
    exp_33_ram[2809] = 19;
    exp_33_ram[2810] = 147;
    exp_33_ram[2811] = 35;
    exp_33_ram[2812] = 35;
    exp_33_ram[2813] = 3;
    exp_33_ram[2814] = 131;
    exp_33_ram[2815] = 3;
    exp_33_ram[2816] = 131;
    exp_33_ram[2817] = 51;
    exp_33_ram[2818] = 19;
    exp_33_ram[2819] = 51;
    exp_33_ram[2820] = 179;
    exp_33_ram[2821] = 179;
    exp_33_ram[2822] = 147;
    exp_33_ram[2823] = 19;
    exp_33_ram[2824] = 147;
    exp_33_ram[2825] = 183;
    exp_33_ram[2826] = 35;
    exp_33_ram[2827] = 35;
    exp_33_ram[2828] = 19;
    exp_33_ram[2829] = 131;
    exp_33_ram[2830] = 3;
    exp_33_ram[2831] = 3;
    exp_33_ram[2832] = 131;
    exp_33_ram[2833] = 19;
    exp_33_ram[2834] = 103;
    exp_33_ram[2835] = 19;
    exp_33_ram[2836] = 35;
    exp_33_ram[2837] = 35;
    exp_33_ram[2838] = 19;
    exp_33_ram[2839] = 35;
    exp_33_ram[2840] = 183;
    exp_33_ram[2841] = 147;
    exp_33_ram[2842] = 3;
    exp_33_ram[2843] = 131;
    exp_33_ram[2844] = 3;
    exp_33_ram[2845] = 131;
    exp_33_ram[2846] = 3;
    exp_33_ram[2847] = 35;
    exp_33_ram[2848] = 35;
    exp_33_ram[2849] = 35;
    exp_33_ram[2850] = 35;
    exp_33_ram[2851] = 35;
    exp_33_ram[2852] = 131;
    exp_33_ram[2853] = 35;
    exp_33_ram[2854] = 183;
    exp_33_ram[2855] = 147;
    exp_33_ram[2856] = 3;
    exp_33_ram[2857] = 3;
    exp_33_ram[2858] = 131;
    exp_33_ram[2859] = 3;
    exp_33_ram[2860] = 3;
    exp_33_ram[2861] = 131;
    exp_33_ram[2862] = 3;
    exp_33_ram[2863] = 131;
    exp_33_ram[2864] = 3;
    exp_33_ram[2865] = 35;
    exp_33_ram[2866] = 35;
    exp_33_ram[2867] = 35;
    exp_33_ram[2868] = 35;
    exp_33_ram[2869] = 35;
    exp_33_ram[2870] = 35;
    exp_33_ram[2871] = 35;
    exp_33_ram[2872] = 35;
    exp_33_ram[2873] = 35;
    exp_33_ram[2874] = 131;
    exp_33_ram[2875] = 35;
    exp_33_ram[2876] = 35;
    exp_33_ram[2877] = 111;
    exp_33_ram[2878] = 131;
    exp_33_ram[2879] = 3;
    exp_33_ram[2880] = 147;
    exp_33_ram[2881] = 147;
    exp_33_ram[2882] = 51;
    exp_33_ram[2883] = 131;
    exp_33_ram[2884] = 179;
    exp_33_ram[2885] = 19;
    exp_33_ram[2886] = 179;
    exp_33_ram[2887] = 3;
    exp_33_ram[2888] = 183;
    exp_33_ram[2889] = 147;
    exp_33_ram[2890] = 131;
    exp_33_ram[2891] = 179;
    exp_33_ram[2892] = 35;
    exp_33_ram[2893] = 131;
    exp_33_ram[2894] = 147;
    exp_33_ram[2895] = 35;
    exp_33_ram[2896] = 3;
    exp_33_ram[2897] = 147;
    exp_33_ram[2898] = 227;
    exp_33_ram[2899] = 183;
    exp_33_ram[2900] = 147;
    exp_33_ram[2901] = 19;
    exp_33_ram[2902] = 163;
    exp_33_ram[2903] = 35;
    exp_33_ram[2904] = 111;
    exp_33_ram[2905] = 131;
    exp_33_ram[2906] = 3;
    exp_33_ram[2907] = 147;
    exp_33_ram[2908] = 147;
    exp_33_ram[2909] = 51;
    exp_33_ram[2910] = 131;
    exp_33_ram[2911] = 51;
    exp_33_ram[2912] = 131;
    exp_33_ram[2913] = 147;
    exp_33_ram[2914] = 147;
    exp_33_ram[2915] = 51;
    exp_33_ram[2916] = 3;
    exp_33_ram[2917] = 183;
    exp_33_ram[2918] = 147;
    exp_33_ram[2919] = 179;
    exp_33_ram[2920] = 35;
    exp_33_ram[2921] = 131;
    exp_33_ram[2922] = 147;
    exp_33_ram[2923] = 35;
    exp_33_ram[2924] = 3;
    exp_33_ram[2925] = 147;
    exp_33_ram[2926] = 227;
    exp_33_ram[2927] = 183;
    exp_33_ram[2928] = 147;
    exp_33_ram[2929] = 19;
    exp_33_ram[2930] = 163;
    exp_33_ram[2931] = 131;
    exp_33_ram[2932] = 131;
    exp_33_ram[2933] = 147;
    exp_33_ram[2934] = 19;
    exp_33_ram[2935] = 239;
    exp_33_ram[2936] = 19;
    exp_33_ram[2937] = 147;
    exp_33_ram[2938] = 35;
    exp_33_ram[2939] = 35;
    exp_33_ram[2940] = 131;
    exp_33_ram[2941] = 147;
    exp_33_ram[2942] = 147;
    exp_33_ram[2943] = 19;
    exp_33_ram[2944] = 183;
    exp_33_ram[2945] = 147;
    exp_33_ram[2946] = 35;
    exp_33_ram[2947] = 131;
    exp_33_ram[2948] = 147;
    exp_33_ram[2949] = 147;
    exp_33_ram[2950] = 19;
    exp_33_ram[2951] = 183;
    exp_33_ram[2952] = 147;
    exp_33_ram[2953] = 163;
    exp_33_ram[2954] = 183;
    exp_33_ram[2955] = 147;
    exp_33_ram[2956] = 19;
    exp_33_ram[2957] = 35;
    exp_33_ram[2958] = 131;
    exp_33_ram[2959] = 131;
    exp_33_ram[2960] = 147;
    exp_33_ram[2961] = 19;
    exp_33_ram[2962] = 239;
    exp_33_ram[2963] = 19;
    exp_33_ram[2964] = 147;
    exp_33_ram[2965] = 35;
    exp_33_ram[2966] = 35;
    exp_33_ram[2967] = 131;
    exp_33_ram[2968] = 147;
    exp_33_ram[2969] = 147;
    exp_33_ram[2970] = 19;
    exp_33_ram[2971] = 183;
    exp_33_ram[2972] = 147;
    exp_33_ram[2973] = 163;
    exp_33_ram[2974] = 131;
    exp_33_ram[2975] = 147;
    exp_33_ram[2976] = 147;
    exp_33_ram[2977] = 19;
    exp_33_ram[2978] = 183;
    exp_33_ram[2979] = 147;
    exp_33_ram[2980] = 35;
    exp_33_ram[2981] = 183;
    exp_33_ram[2982] = 147;
    exp_33_ram[2983] = 19;
    exp_33_ram[2984] = 163;
    exp_33_ram[2985] = 131;
    exp_33_ram[2986] = 131;
    exp_33_ram[2987] = 147;
    exp_33_ram[2988] = 19;
    exp_33_ram[2989] = 239;
    exp_33_ram[2990] = 19;
    exp_33_ram[2991] = 147;
    exp_33_ram[2992] = 35;
    exp_33_ram[2993] = 35;
    exp_33_ram[2994] = 131;
    exp_33_ram[2995] = 147;
    exp_33_ram[2996] = 147;
    exp_33_ram[2997] = 19;
    exp_33_ram[2998] = 183;
    exp_33_ram[2999] = 147;
    exp_33_ram[3000] = 35;
    exp_33_ram[3001] = 131;
    exp_33_ram[3002] = 147;
    exp_33_ram[3003] = 147;
    exp_33_ram[3004] = 19;
    exp_33_ram[3005] = 183;
    exp_33_ram[3006] = 147;
    exp_33_ram[3007] = 163;
    exp_33_ram[3008] = 183;
    exp_33_ram[3009] = 147;
    exp_33_ram[3010] = 19;
    exp_33_ram[3011] = 35;
    exp_33_ram[3012] = 131;
    exp_33_ram[3013] = 131;
    exp_33_ram[3014] = 147;
    exp_33_ram[3015] = 19;
    exp_33_ram[3016] = 239;
    exp_33_ram[3017] = 19;
    exp_33_ram[3018] = 147;
    exp_33_ram[3019] = 35;
    exp_33_ram[3020] = 35;
    exp_33_ram[3021] = 131;
    exp_33_ram[3022] = 147;
    exp_33_ram[3023] = 147;
    exp_33_ram[3024] = 19;
    exp_33_ram[3025] = 183;
    exp_33_ram[3026] = 147;
    exp_33_ram[3027] = 163;
    exp_33_ram[3028] = 131;
    exp_33_ram[3029] = 147;
    exp_33_ram[3030] = 147;
    exp_33_ram[3031] = 19;
    exp_33_ram[3032] = 183;
    exp_33_ram[3033] = 147;
    exp_33_ram[3034] = 35;
    exp_33_ram[3035] = 183;
    exp_33_ram[3036] = 147;
    exp_33_ram[3037] = 19;
    exp_33_ram[3038] = 163;
    exp_33_ram[3039] = 131;
    exp_33_ram[3040] = 131;
    exp_33_ram[3041] = 147;
    exp_33_ram[3042] = 147;
    exp_33_ram[3043] = 19;
    exp_33_ram[3044] = 239;
    exp_33_ram[3045] = 19;
    exp_33_ram[3046] = 147;
    exp_33_ram[3047] = 35;
    exp_33_ram[3048] = 35;
    exp_33_ram[3049] = 131;
    exp_33_ram[3050] = 147;
    exp_33_ram[3051] = 147;
    exp_33_ram[3052] = 19;
    exp_33_ram[3053] = 183;
    exp_33_ram[3054] = 147;
    exp_33_ram[3055] = 35;
    exp_33_ram[3056] = 131;
    exp_33_ram[3057] = 147;
    exp_33_ram[3058] = 19;
    exp_33_ram[3059] = 239;
    exp_33_ram[3060] = 19;
    exp_33_ram[3061] = 147;
    exp_33_ram[3062] = 35;
    exp_33_ram[3063] = 35;
    exp_33_ram[3064] = 131;
    exp_33_ram[3065] = 147;
    exp_33_ram[3066] = 147;
    exp_33_ram[3067] = 19;
    exp_33_ram[3068] = 183;
    exp_33_ram[3069] = 147;
    exp_33_ram[3070] = 163;
    exp_33_ram[3071] = 131;
    exp_33_ram[3072] = 147;
    exp_33_ram[3073] = 19;
    exp_33_ram[3074] = 239;
    exp_33_ram[3075] = 19;
    exp_33_ram[3076] = 147;
    exp_33_ram[3077] = 35;
    exp_33_ram[3078] = 35;
    exp_33_ram[3079] = 131;
    exp_33_ram[3080] = 147;
    exp_33_ram[3081] = 147;
    exp_33_ram[3082] = 19;
    exp_33_ram[3083] = 183;
    exp_33_ram[3084] = 147;
    exp_33_ram[3085] = 35;
    exp_33_ram[3086] = 131;
    exp_33_ram[3087] = 147;
    exp_33_ram[3088] = 147;
    exp_33_ram[3089] = 19;
    exp_33_ram[3090] = 183;
    exp_33_ram[3091] = 147;
    exp_33_ram[3092] = 163;
    exp_33_ram[3093] = 183;
    exp_33_ram[3094] = 147;
    exp_33_ram[3095] = 19;
    exp_33_ram[3096] = 35;
    exp_33_ram[3097] = 183;
    exp_33_ram[3098] = 147;
    exp_33_ram[3099] = 163;
    exp_33_ram[3100] = 183;
    exp_33_ram[3101] = 147;
    exp_33_ram[3102] = 19;
    exp_33_ram[3103] = 131;
    exp_33_ram[3104] = 3;
    exp_33_ram[3105] = 19;
    exp_33_ram[3106] = 103;
    exp_33_ram[3107] = 19;
    exp_33_ram[3108] = 35;
    exp_33_ram[3109] = 35;
    exp_33_ram[3110] = 19;
    exp_33_ram[3111] = 35;
    exp_33_ram[3112] = 3;
    exp_33_ram[3113] = 239;
    exp_33_ram[3114] = 147;
    exp_33_ram[3115] = 19;
    exp_33_ram[3116] = 239;
    exp_33_ram[3117] = 147;
    exp_33_ram[3118] = 19;
    exp_33_ram[3119] = 131;
    exp_33_ram[3120] = 3;
    exp_33_ram[3121] = 19;
    exp_33_ram[3122] = 103;
    exp_33_ram[3123] = 19;
    exp_33_ram[3124] = 35;
    exp_33_ram[3125] = 35;
    exp_33_ram[3126] = 35;
    exp_33_ram[3127] = 35;
    exp_33_ram[3128] = 35;
    exp_33_ram[3129] = 35;
    exp_33_ram[3130] = 35;
    exp_33_ram[3131] = 35;
    exp_33_ram[3132] = 35;
    exp_33_ram[3133] = 35;
    exp_33_ram[3134] = 19;
    exp_33_ram[3135] = 35;
    exp_33_ram[3136] = 35;
    exp_33_ram[3137] = 35;
    exp_33_ram[3138] = 147;
    exp_33_ram[3139] = 35;
    exp_33_ram[3140] = 147;
    exp_33_ram[3141] = 35;
    exp_33_ram[3142] = 131;
    exp_33_ram[3143] = 19;
    exp_33_ram[3144] = 239;
    exp_33_ram[3145] = 35;
    exp_33_ram[3146] = 3;
    exp_33_ram[3147] = 183;
    exp_33_ram[3148] = 147;
    exp_33_ram[3149] = 179;
    exp_33_ram[3150] = 35;
    exp_33_ram[3151] = 131;
    exp_33_ram[3152] = 19;
    exp_33_ram[3153] = 147;
    exp_33_ram[3154] = 131;
    exp_33_ram[3155] = 19;
    exp_33_ram[3156] = 99;
    exp_33_ram[3157] = 131;
    exp_33_ram[3158] = 19;
    exp_33_ram[3159] = 99;
    exp_33_ram[3160] = 131;
    exp_33_ram[3161] = 19;
    exp_33_ram[3162] = 99;
    exp_33_ram[3163] = 131;
    exp_33_ram[3164] = 147;
    exp_33_ram[3165] = 35;
    exp_33_ram[3166] = 131;
    exp_33_ram[3167] = 19;
    exp_33_ram[3168] = 131;
    exp_33_ram[3169] = 179;
    exp_33_ram[3170] = 35;
    exp_33_ram[3171] = 131;
    exp_33_ram[3172] = 19;
    exp_33_ram[3173] = 147;
    exp_33_ram[3174] = 3;
    exp_33_ram[3175] = 131;
    exp_33_ram[3176] = 51;
    exp_33_ram[3177] = 147;
    exp_33_ram[3178] = 179;
    exp_33_ram[3179] = 179;
    exp_33_ram[3180] = 179;
    exp_33_ram[3181] = 147;
    exp_33_ram[3182] = 35;
    exp_33_ram[3183] = 35;
    exp_33_ram[3184] = 111;
    exp_33_ram[3185] = 19;
    exp_33_ram[3186] = 35;
    exp_33_ram[3187] = 35;
    exp_33_ram[3188] = 131;
    exp_33_ram[3189] = 19;
    exp_33_ram[3190] = 131;
    exp_33_ram[3191] = 147;
    exp_33_ram[3192] = 19;
    exp_33_ram[3193] = 239;
    exp_33_ram[3194] = 35;
    exp_33_ram[3195] = 3;
    exp_33_ram[3196] = 183;
    exp_33_ram[3197] = 147;
    exp_33_ram[3198] = 179;
    exp_33_ram[3199] = 35;
    exp_33_ram[3200] = 131;
    exp_33_ram[3201] = 19;
    exp_33_ram[3202] = 147;
    exp_33_ram[3203] = 131;
    exp_33_ram[3204] = 19;
    exp_33_ram[3205] = 99;
    exp_33_ram[3206] = 131;
    exp_33_ram[3207] = 19;
    exp_33_ram[3208] = 99;
    exp_33_ram[3209] = 131;
    exp_33_ram[3210] = 19;
    exp_33_ram[3211] = 99;
    exp_33_ram[3212] = 131;
    exp_33_ram[3213] = 147;
    exp_33_ram[3214] = 35;
    exp_33_ram[3215] = 131;
    exp_33_ram[3216] = 19;
    exp_33_ram[3217] = 131;
    exp_33_ram[3218] = 179;
    exp_33_ram[3219] = 35;
    exp_33_ram[3220] = 131;
    exp_33_ram[3221] = 19;
    exp_33_ram[3222] = 131;
    exp_33_ram[3223] = 179;
    exp_33_ram[3224] = 35;
    exp_33_ram[3225] = 131;
    exp_33_ram[3226] = 19;
    exp_33_ram[3227] = 147;
    exp_33_ram[3228] = 3;
    exp_33_ram[3229] = 131;
    exp_33_ram[3230] = 51;
    exp_33_ram[3231] = 147;
    exp_33_ram[3232] = 179;
    exp_33_ram[3233] = 179;
    exp_33_ram[3234] = 179;
    exp_33_ram[3235] = 147;
    exp_33_ram[3236] = 35;
    exp_33_ram[3237] = 35;
    exp_33_ram[3238] = 111;
    exp_33_ram[3239] = 19;
    exp_33_ram[3240] = 131;
    exp_33_ram[3241] = 147;
    exp_33_ram[3242] = 35;
    exp_33_ram[3243] = 3;
    exp_33_ram[3244] = 183;
    exp_33_ram[3245] = 147;
    exp_33_ram[3246] = 19;
    exp_33_ram[3247] = 239;
    exp_33_ram[3248] = 19;
    exp_33_ram[3249] = 147;
    exp_33_ram[3250] = 35;
    exp_33_ram[3251] = 35;
    exp_33_ram[3252] = 131;
    exp_33_ram[3253] = 147;
    exp_33_ram[3254] = 35;
    exp_33_ram[3255] = 3;
    exp_33_ram[3256] = 131;
    exp_33_ram[3257] = 179;
    exp_33_ram[3258] = 35;
    exp_33_ram[3259] = 3;
    exp_33_ram[3260] = 147;
    exp_33_ram[3261] = 179;
    exp_33_ram[3262] = 35;
    exp_33_ram[3263] = 3;
    exp_33_ram[3264] = 131;
    exp_33_ram[3265] = 179;
    exp_33_ram[3266] = 35;
    exp_33_ram[3267] = 131;
    exp_33_ram[3268] = 35;
    exp_33_ram[3269] = 147;
    exp_33_ram[3270] = 35;
    exp_33_ram[3271] = 3;
    exp_33_ram[3272] = 183;
    exp_33_ram[3273] = 147;
    exp_33_ram[3274] = 19;
    exp_33_ram[3275] = 239;
    exp_33_ram[3276] = 19;
    exp_33_ram[3277] = 147;
    exp_33_ram[3278] = 35;
    exp_33_ram[3279] = 35;
    exp_33_ram[3280] = 131;
    exp_33_ram[3281] = 35;
    exp_33_ram[3282] = 131;
    exp_33_ram[3283] = 35;
    exp_33_ram[3284] = 147;
    exp_33_ram[3285] = 35;
    exp_33_ram[3286] = 131;
    exp_33_ram[3287] = 147;
    exp_33_ram[3288] = 19;
    exp_33_ram[3289] = 239;
    exp_33_ram[3290] = 19;
    exp_33_ram[3291] = 147;
    exp_33_ram[3292] = 35;
    exp_33_ram[3293] = 35;
    exp_33_ram[3294] = 131;
    exp_33_ram[3295] = 35;
    exp_33_ram[3296] = 131;
    exp_33_ram[3297] = 35;
    exp_33_ram[3298] = 147;
    exp_33_ram[3299] = 35;
    exp_33_ram[3300] = 131;
    exp_33_ram[3301] = 35;
    exp_33_ram[3302] = 131;
    exp_33_ram[3303] = 3;
    exp_33_ram[3304] = 3;
    exp_33_ram[3305] = 131;
    exp_33_ram[3306] = 3;
    exp_33_ram[3307] = 3;
    exp_33_ram[3308] = 131;
    exp_33_ram[3309] = 3;
    exp_33_ram[3310] = 131;
    exp_33_ram[3311] = 3;
    exp_33_ram[3312] = 35;
    exp_33_ram[3313] = 35;
    exp_33_ram[3314] = 35;
    exp_33_ram[3315] = 35;
    exp_33_ram[3316] = 35;
    exp_33_ram[3317] = 35;
    exp_33_ram[3318] = 35;
    exp_33_ram[3319] = 35;
    exp_33_ram[3320] = 35;
    exp_33_ram[3321] = 3;
    exp_33_ram[3322] = 131;
    exp_33_ram[3323] = 3;
    exp_33_ram[3324] = 3;
    exp_33_ram[3325] = 131;
    exp_33_ram[3326] = 3;
    exp_33_ram[3327] = 131;
    exp_33_ram[3328] = 3;
    exp_33_ram[3329] = 131;
    exp_33_ram[3330] = 3;
    exp_33_ram[3331] = 131;
    exp_33_ram[3332] = 19;
    exp_33_ram[3333] = 103;
    exp_33_ram[3334] = 19;
    exp_33_ram[3335] = 35;
    exp_33_ram[3336] = 35;
    exp_33_ram[3337] = 35;
    exp_33_ram[3338] = 35;
    exp_33_ram[3339] = 35;
    exp_33_ram[3340] = 19;
    exp_33_ram[3341] = 35;
    exp_33_ram[3342] = 147;
    exp_33_ram[3343] = 19;
    exp_33_ram[3344] = 35;
    exp_33_ram[3345] = 35;
    exp_33_ram[3346] = 131;
    exp_33_ram[3347] = 3;
    exp_33_ram[3348] = 131;
    exp_33_ram[3349] = 35;
    exp_33_ram[3350] = 35;
    exp_33_ram[3351] = 3;
    exp_33_ram[3352] = 131;
    exp_33_ram[3353] = 239;
    exp_33_ram[3354] = 147;
    exp_33_ram[3355] = 99;
    exp_33_ram[3356] = 55;
    exp_33_ram[3357] = 19;
    exp_33_ram[3358] = 147;
    exp_33_ram[3359] = 35;
    exp_33_ram[3360] = 35;
    exp_33_ram[3361] = 183;
    exp_33_ram[3362] = 131;
    exp_33_ram[3363] = 19;
    exp_33_ram[3364] = 147;
    exp_33_ram[3365] = 147;
    exp_33_ram[3366] = 3;
    exp_33_ram[3367] = 131;
    exp_33_ram[3368] = 51;
    exp_33_ram[3369] = 147;
    exp_33_ram[3370] = 179;
    exp_33_ram[3371] = 179;
    exp_33_ram[3372] = 179;
    exp_33_ram[3373] = 147;
    exp_33_ram[3374] = 19;
    exp_33_ram[3375] = 147;
    exp_33_ram[3376] = 3;
    exp_33_ram[3377] = 131;
    exp_33_ram[3378] = 51;
    exp_33_ram[3379] = 19;
    exp_33_ram[3380] = 51;
    exp_33_ram[3381] = 179;
    exp_33_ram[3382] = 179;
    exp_33_ram[3383] = 147;
    exp_33_ram[3384] = 35;
    exp_33_ram[3385] = 35;
    exp_33_ram[3386] = 183;
    exp_33_ram[3387] = 147;
    exp_33_ram[3388] = 147;
    exp_33_ram[3389] = 131;
    exp_33_ram[3390] = 3;
    exp_33_ram[3391] = 19;
    exp_33_ram[3392] = 239;
    exp_33_ram[3393] = 3;
    exp_33_ram[3394] = 131;
    exp_33_ram[3395] = 3;
    exp_33_ram[3396] = 3;
    exp_33_ram[3397] = 131;
    exp_33_ram[3398] = 3;
    exp_33_ram[3399] = 131;
    exp_33_ram[3400] = 3;
    exp_33_ram[3401] = 131;
    exp_33_ram[3402] = 35;
    exp_33_ram[3403] = 35;
    exp_33_ram[3404] = 35;
    exp_33_ram[3405] = 35;
    exp_33_ram[3406] = 35;
    exp_33_ram[3407] = 35;
    exp_33_ram[3408] = 35;
    exp_33_ram[3409] = 35;
    exp_33_ram[3410] = 35;
    exp_33_ram[3411] = 3;
    exp_33_ram[3412] = 131;
    exp_33_ram[3413] = 239;
    exp_33_ram[3414] = 19;
    exp_33_ram[3415] = 183;
    exp_33_ram[3416] = 147;
    exp_33_ram[3417] = 35;
    exp_33_ram[3418] = 183;
    exp_33_ram[3419] = 147;
    exp_33_ram[3420] = 19;
    exp_33_ram[3421] = 131;
    exp_33_ram[3422] = 3;
    exp_33_ram[3423] = 131;
    exp_33_ram[3424] = 3;
    exp_33_ram[3425] = 131;
    exp_33_ram[3426] = 19;
    exp_33_ram[3427] = 103;
    exp_33_ram[3428] = 19;
    exp_33_ram[3429] = 35;
    exp_33_ram[3430] = 35;
    exp_33_ram[3431] = 19;
    exp_33_ram[3432] = 35;
    exp_33_ram[3433] = 35;
    exp_33_ram[3434] = 3;
    exp_33_ram[3435] = 239;
    exp_33_ram[3436] = 147;
    exp_33_ram[3437] = 163;
    exp_33_ram[3438] = 131;
    exp_33_ram[3439] = 19;
    exp_33_ram[3440] = 147;
    exp_33_ram[3441] = 99;
    exp_33_ram[3442] = 3;
    exp_33_ram[3443] = 147;
    exp_33_ram[3444] = 147;
    exp_33_ram[3445] = 179;
    exp_33_ram[3446] = 147;
    exp_33_ram[3447] = 35;
    exp_33_ram[3448] = 3;
    exp_33_ram[3449] = 131;
    exp_33_ram[3450] = 179;
    exp_33_ram[3451] = 147;
    exp_33_ram[3452] = 35;
    exp_33_ram[3453] = 111;
    exp_33_ram[3454] = 19;
    exp_33_ram[3455] = 131;
    exp_33_ram[3456] = 19;
    exp_33_ram[3457] = 131;
    exp_33_ram[3458] = 3;
    exp_33_ram[3459] = 19;
    exp_33_ram[3460] = 103;
    exp_33_ram[3461] = 19;
    exp_33_ram[3462] = 35;
    exp_33_ram[3463] = 35;
    exp_33_ram[3464] = 19;
    exp_33_ram[3465] = 183;
    exp_33_ram[3466] = 131;
    exp_33_ram[3467] = 19;
    exp_33_ram[3468] = 239;
    exp_33_ram[3469] = 147;
    exp_33_ram[3470] = 19;
    exp_33_ram[3471] = 131;
    exp_33_ram[3472] = 3;
    exp_33_ram[3473] = 19;
    exp_33_ram[3474] = 103;
    exp_33_ram[3475] = 19;
    exp_33_ram[3476] = 35;
    exp_33_ram[3477] = 35;
    exp_33_ram[3478] = 35;
    exp_33_ram[3479] = 35;
    exp_33_ram[3480] = 19;
    exp_33_ram[3481] = 35;
    exp_33_ram[3482] = 239;
    exp_33_ram[3483] = 35;
    exp_33_ram[3484] = 35;
    exp_33_ram[3485] = 19;
    exp_33_ram[3486] = 239;
    exp_33_ram[3487] = 19;
    exp_33_ram[3488] = 147;
    exp_33_ram[3489] = 3;
    exp_33_ram[3490] = 131;
    exp_33_ram[3491] = 51;
    exp_33_ram[3492] = 19;
    exp_33_ram[3493] = 51;
    exp_33_ram[3494] = 179;
    exp_33_ram[3495] = 179;
    exp_33_ram[3496] = 147;
    exp_33_ram[3497] = 131;
    exp_33_ram[3498] = 19;
    exp_33_ram[3499] = 147;
    exp_33_ram[3500] = 19;
    exp_33_ram[3501] = 147;
    exp_33_ram[3502] = 227;
    exp_33_ram[3503] = 19;
    exp_33_ram[3504] = 147;
    exp_33_ram[3505] = 99;
    exp_33_ram[3506] = 147;
    exp_33_ram[3507] = 147;
    exp_33_ram[3508] = 227;
    exp_33_ram[3509] = 19;
    exp_33_ram[3510] = 19;
    exp_33_ram[3511] = 131;
    exp_33_ram[3512] = 3;
    exp_33_ram[3513] = 3;
    exp_33_ram[3514] = 131;
    exp_33_ram[3515] = 19;
    exp_33_ram[3516] = 103;
    exp_33_ram[3517] = 19;
    exp_33_ram[3518] = 35;
    exp_33_ram[3519] = 35;
    exp_33_ram[3520] = 19;
    exp_33_ram[3521] = 183;
    exp_33_ram[3522] = 19;
    exp_33_ram[3523] = 239;
    exp_33_ram[3524] = 19;
    exp_33_ram[3525] = 131;
    exp_33_ram[3526] = 3;
    exp_33_ram[3527] = 19;
    exp_33_ram[3528] = 103;
    exp_33_ram[3529] = 19;
    exp_33_ram[3530] = 35;
    exp_33_ram[3531] = 35;
    exp_33_ram[3532] = 19;
    exp_33_ram[3533] = 183;
    exp_33_ram[3534] = 19;
    exp_33_ram[3535] = 239;
    exp_33_ram[3536] = 147;
    exp_33_ram[3537] = 35;
    exp_33_ram[3538] = 35;
    exp_33_ram[3539] = 111;
    exp_33_ram[3540] = 131;
    exp_33_ram[3541] = 183;
    exp_33_ram[3542] = 19;
    exp_33_ram[3543] = 239;
    exp_33_ram[3544] = 111;
    exp_33_ram[3545] = 131;
    exp_33_ram[3546] = 147;
    exp_33_ram[3547] = 35;
    exp_33_ram[3548] = 183;
    exp_33_ram[3549] = 131;
    exp_33_ram[3550] = 147;
    exp_33_ram[3551] = 3;
    exp_33_ram[3552] = 239;
    exp_33_ram[3553] = 183;
    exp_33_ram[3554] = 3;
    exp_33_ram[3555] = 147;
    exp_33_ram[3556] = 179;
    exp_33_ram[3557] = 19;
    exp_33_ram[3558] = 239;
    exp_33_ram[3559] = 3;
    exp_33_ram[3560] = 147;
    exp_33_ram[3561] = 227;
    exp_33_ram[3562] = 111;
    exp_33_ram[3563] = 131;
    exp_33_ram[3564] = 147;
    exp_33_ram[3565] = 35;
    exp_33_ram[3566] = 183;
    exp_33_ram[3567] = 131;
    exp_33_ram[3568] = 147;
    exp_33_ram[3569] = 3;
    exp_33_ram[3570] = 239;
    exp_33_ram[3571] = 183;
    exp_33_ram[3572] = 3;
    exp_33_ram[3573] = 147;
    exp_33_ram[3574] = 179;
    exp_33_ram[3575] = 19;
    exp_33_ram[3576] = 239;
    exp_33_ram[3577] = 3;
    exp_33_ram[3578] = 147;
    exp_33_ram[3579] = 227;
    exp_33_ram[3580] = 131;
    exp_33_ram[3581] = 147;
    exp_33_ram[3582] = 35;
    exp_33_ram[3583] = 3;
    exp_33_ram[3584] = 147;
    exp_33_ram[3585] = 227;
    exp_33_ram[3586] = 183;
    exp_33_ram[3587] = 131;
    exp_33_ram[3588] = 147;
    exp_33_ram[3589] = 19;
    exp_33_ram[3590] = 239;
    exp_33_ram[3591] = 19;
    exp_33_ram[3592] = 131;
    exp_33_ram[3593] = 3;
    exp_33_ram[3594] = 19;
    exp_33_ram[3595] = 103;
    exp_33_ram[3596] = 19;
    exp_33_ram[3597] = 35;
    exp_33_ram[3598] = 35;
    exp_33_ram[3599] = 35;
    exp_33_ram[3600] = 35;
    exp_33_ram[3601] = 35;
    exp_33_ram[3602] = 35;
    exp_33_ram[3603] = 35;
    exp_33_ram[3604] = 35;
    exp_33_ram[3605] = 35;
    exp_33_ram[3606] = 35;
    exp_33_ram[3607] = 35;
    exp_33_ram[3608] = 35;
    exp_33_ram[3609] = 19;
    exp_33_ram[3610] = 147;
    exp_33_ram[3611] = 35;
    exp_33_ram[3612] = 19;
    exp_33_ram[3613] = 147;
    exp_33_ram[3614] = 35;
    exp_33_ram[3615] = 35;
    exp_33_ram[3616] = 239;
    exp_33_ram[3617] = 35;
    exp_33_ram[3618] = 35;
    exp_33_ram[3619] = 35;
    exp_33_ram[3620] = 111;
    exp_33_ram[3621] = 3;
    exp_33_ram[3622] = 183;
    exp_33_ram[3623] = 147;
    exp_33_ram[3624] = 179;
    exp_33_ram[3625] = 35;
    exp_33_ram[3626] = 3;
    exp_33_ram[3627] = 183;
    exp_33_ram[3628] = 147;
    exp_33_ram[3629] = 179;
    exp_33_ram[3630] = 35;
    exp_33_ram[3631] = 3;
    exp_33_ram[3632] = 183;
    exp_33_ram[3633] = 147;
    exp_33_ram[3634] = 179;
    exp_33_ram[3635] = 35;
    exp_33_ram[3636] = 3;
    exp_33_ram[3637] = 183;
    exp_33_ram[3638] = 147;
    exp_33_ram[3639] = 179;
    exp_33_ram[3640] = 35;
    exp_33_ram[3641] = 131;
    exp_33_ram[3642] = 147;
    exp_33_ram[3643] = 35;
    exp_33_ram[3644] = 239;
    exp_33_ram[3645] = 19;
    exp_33_ram[3646] = 147;
    exp_33_ram[3647] = 3;
    exp_33_ram[3648] = 131;
    exp_33_ram[3649] = 51;
    exp_33_ram[3650] = 19;
    exp_33_ram[3651] = 51;
    exp_33_ram[3652] = 179;
    exp_33_ram[3653] = 179;
    exp_33_ram[3654] = 147;
    exp_33_ram[3655] = 183;
    exp_33_ram[3656] = 131;
    exp_33_ram[3657] = 35;
    exp_33_ram[3658] = 35;
    exp_33_ram[3659] = 3;
    exp_33_ram[3660] = 131;
    exp_33_ram[3661] = 19;
    exp_33_ram[3662] = 147;
    exp_33_ram[3663] = 227;
    exp_33_ram[3664] = 19;
    exp_33_ram[3665] = 147;
    exp_33_ram[3666] = 99;
    exp_33_ram[3667] = 147;
    exp_33_ram[3668] = 147;
    exp_33_ram[3669] = 227;
    exp_33_ram[3670] = 131;
    exp_33_ram[3671] = 183;
    exp_33_ram[3672] = 19;
    exp_33_ram[3673] = 239;
    exp_33_ram[3674] = 239;
    exp_33_ram[3675] = 35;
    exp_33_ram[3676] = 35;
    exp_33_ram[3677] = 35;
    exp_33_ram[3678] = 111;
    exp_33_ram[3679] = 3;
    exp_33_ram[3680] = 131;
    exp_33_ram[3681] = 183;
    exp_33_ram[3682] = 147;
    exp_33_ram[3683] = 51;
    exp_33_ram[3684] = 147;
    exp_33_ram[3685] = 179;
    exp_33_ram[3686] = 51;
    exp_33_ram[3687] = 183;
    exp_33_ram[3688] = 147;
    exp_33_ram[3689] = 179;
    exp_33_ram[3690] = 179;
    exp_33_ram[3691] = 19;
    exp_33_ram[3692] = 179;
    exp_33_ram[3693] = 147;
    exp_33_ram[3694] = 35;
    exp_33_ram[3695] = 35;
    exp_33_ram[3696] = 3;
    exp_33_ram[3697] = 131;
    exp_33_ram[3698] = 183;
    exp_33_ram[3699] = 147;
    exp_33_ram[3700] = 51;
    exp_33_ram[3701] = 147;
    exp_33_ram[3702] = 179;
    exp_33_ram[3703] = 51;
    exp_33_ram[3704] = 183;
    exp_33_ram[3705] = 147;
    exp_33_ram[3706] = 179;
    exp_33_ram[3707] = 179;
    exp_33_ram[3708] = 19;
    exp_33_ram[3709] = 179;
    exp_33_ram[3710] = 147;
    exp_33_ram[3711] = 35;
    exp_33_ram[3712] = 35;
    exp_33_ram[3713] = 3;
    exp_33_ram[3714] = 131;
    exp_33_ram[3715] = 183;
    exp_33_ram[3716] = 147;
    exp_33_ram[3717] = 51;
    exp_33_ram[3718] = 147;
    exp_33_ram[3719] = 179;
    exp_33_ram[3720] = 51;
    exp_33_ram[3721] = 183;
    exp_33_ram[3722] = 147;
    exp_33_ram[3723] = 179;
    exp_33_ram[3724] = 179;
    exp_33_ram[3725] = 19;
    exp_33_ram[3726] = 179;
    exp_33_ram[3727] = 147;
    exp_33_ram[3728] = 35;
    exp_33_ram[3729] = 35;
    exp_33_ram[3730] = 3;
    exp_33_ram[3731] = 131;
    exp_33_ram[3732] = 183;
    exp_33_ram[3733] = 147;
    exp_33_ram[3734] = 51;
    exp_33_ram[3735] = 147;
    exp_33_ram[3736] = 179;
    exp_33_ram[3737] = 51;
    exp_33_ram[3738] = 183;
    exp_33_ram[3739] = 147;
    exp_33_ram[3740] = 179;
    exp_33_ram[3741] = 179;
    exp_33_ram[3742] = 19;
    exp_33_ram[3743] = 179;
    exp_33_ram[3744] = 147;
    exp_33_ram[3745] = 35;
    exp_33_ram[3746] = 35;
    exp_33_ram[3747] = 131;
    exp_33_ram[3748] = 147;
    exp_33_ram[3749] = 35;
    exp_33_ram[3750] = 239;
    exp_33_ram[3751] = 19;
    exp_33_ram[3752] = 147;
    exp_33_ram[3753] = 3;
    exp_33_ram[3754] = 131;
    exp_33_ram[3755] = 51;
    exp_33_ram[3756] = 19;
    exp_33_ram[3757] = 51;
    exp_33_ram[3758] = 179;
    exp_33_ram[3759] = 179;
    exp_33_ram[3760] = 147;
    exp_33_ram[3761] = 183;
    exp_33_ram[3762] = 131;
    exp_33_ram[3763] = 35;
    exp_33_ram[3764] = 35;
    exp_33_ram[3765] = 3;
    exp_33_ram[3766] = 131;
    exp_33_ram[3767] = 19;
    exp_33_ram[3768] = 147;
    exp_33_ram[3769] = 227;
    exp_33_ram[3770] = 19;
    exp_33_ram[3771] = 147;
    exp_33_ram[3772] = 99;
    exp_33_ram[3773] = 147;
    exp_33_ram[3774] = 147;
    exp_33_ram[3775] = 227;
    exp_33_ram[3776] = 131;
    exp_33_ram[3777] = 183;
    exp_33_ram[3778] = 19;
    exp_33_ram[3779] = 239;
    exp_33_ram[3780] = 239;
    exp_33_ram[3781] = 35;
    exp_33_ram[3782] = 35;
    exp_33_ram[3783] = 35;
    exp_33_ram[3784] = 111;
    exp_33_ram[3785] = 3;
    exp_33_ram[3786] = 183;
    exp_33_ram[3787] = 147;
    exp_33_ram[3788] = 179;
    exp_33_ram[3789] = 35;
    exp_33_ram[3790] = 3;
    exp_33_ram[3791] = 183;
    exp_33_ram[3792] = 147;
    exp_33_ram[3793] = 179;
    exp_33_ram[3794] = 35;
    exp_33_ram[3795] = 3;
    exp_33_ram[3796] = 183;
    exp_33_ram[3797] = 147;
    exp_33_ram[3798] = 179;
    exp_33_ram[3799] = 35;
    exp_33_ram[3800] = 3;
    exp_33_ram[3801] = 183;
    exp_33_ram[3802] = 147;
    exp_33_ram[3803] = 179;
    exp_33_ram[3804] = 35;
    exp_33_ram[3805] = 131;
    exp_33_ram[3806] = 147;
    exp_33_ram[3807] = 35;
    exp_33_ram[3808] = 239;
    exp_33_ram[3809] = 19;
    exp_33_ram[3810] = 147;
    exp_33_ram[3811] = 3;
    exp_33_ram[3812] = 131;
    exp_33_ram[3813] = 51;
    exp_33_ram[3814] = 19;
    exp_33_ram[3815] = 51;
    exp_33_ram[3816] = 179;
    exp_33_ram[3817] = 179;
    exp_33_ram[3818] = 147;
    exp_33_ram[3819] = 183;
    exp_33_ram[3820] = 131;
    exp_33_ram[3821] = 35;
    exp_33_ram[3822] = 35;
    exp_33_ram[3823] = 3;
    exp_33_ram[3824] = 131;
    exp_33_ram[3825] = 19;
    exp_33_ram[3826] = 147;
    exp_33_ram[3827] = 227;
    exp_33_ram[3828] = 19;
    exp_33_ram[3829] = 147;
    exp_33_ram[3830] = 99;
    exp_33_ram[3831] = 147;
    exp_33_ram[3832] = 147;
    exp_33_ram[3833] = 227;
    exp_33_ram[3834] = 131;
    exp_33_ram[3835] = 183;
    exp_33_ram[3836] = 19;
    exp_33_ram[3837] = 239;
    exp_33_ram[3838] = 239;
    exp_33_ram[3839] = 35;
    exp_33_ram[3840] = 35;
    exp_33_ram[3841] = 35;
    exp_33_ram[3842] = 111;
    exp_33_ram[3843] = 3;
    exp_33_ram[3844] = 131;
    exp_33_ram[3845] = 55;
    exp_33_ram[3846] = 19;
    exp_33_ram[3847] = 147;
    exp_33_ram[3848] = 19;
    exp_33_ram[3849] = 147;
    exp_33_ram[3850] = 239;
    exp_33_ram[3851] = 19;
    exp_33_ram[3852] = 147;
    exp_33_ram[3853] = 35;
    exp_33_ram[3854] = 35;
    exp_33_ram[3855] = 3;
    exp_33_ram[3856] = 131;
    exp_33_ram[3857] = 55;
    exp_33_ram[3858] = 19;
    exp_33_ram[3859] = 147;
    exp_33_ram[3860] = 19;
    exp_33_ram[3861] = 147;
    exp_33_ram[3862] = 239;
    exp_33_ram[3863] = 19;
    exp_33_ram[3864] = 147;
    exp_33_ram[3865] = 35;
    exp_33_ram[3866] = 35;
    exp_33_ram[3867] = 3;
    exp_33_ram[3868] = 131;
    exp_33_ram[3869] = 55;
    exp_33_ram[3870] = 19;
    exp_33_ram[3871] = 147;
    exp_33_ram[3872] = 19;
    exp_33_ram[3873] = 147;
    exp_33_ram[3874] = 239;
    exp_33_ram[3875] = 19;
    exp_33_ram[3876] = 147;
    exp_33_ram[3877] = 35;
    exp_33_ram[3878] = 35;
    exp_33_ram[3879] = 3;
    exp_33_ram[3880] = 131;
    exp_33_ram[3881] = 55;
    exp_33_ram[3882] = 19;
    exp_33_ram[3883] = 147;
    exp_33_ram[3884] = 19;
    exp_33_ram[3885] = 147;
    exp_33_ram[3886] = 239;
    exp_33_ram[3887] = 19;
    exp_33_ram[3888] = 147;
    exp_33_ram[3889] = 35;
    exp_33_ram[3890] = 35;
    exp_33_ram[3891] = 131;
    exp_33_ram[3892] = 147;
    exp_33_ram[3893] = 35;
    exp_33_ram[3894] = 239;
    exp_33_ram[3895] = 19;
    exp_33_ram[3896] = 147;
    exp_33_ram[3897] = 3;
    exp_33_ram[3898] = 131;
    exp_33_ram[3899] = 51;
    exp_33_ram[3900] = 19;
    exp_33_ram[3901] = 51;
    exp_33_ram[3902] = 179;
    exp_33_ram[3903] = 179;
    exp_33_ram[3904] = 147;
    exp_33_ram[3905] = 183;
    exp_33_ram[3906] = 131;
    exp_33_ram[3907] = 19;
    exp_33_ram[3908] = 147;
    exp_33_ram[3909] = 19;
    exp_33_ram[3910] = 147;
    exp_33_ram[3911] = 227;
    exp_33_ram[3912] = 19;
    exp_33_ram[3913] = 147;
    exp_33_ram[3914] = 99;
    exp_33_ram[3915] = 147;
    exp_33_ram[3916] = 147;
    exp_33_ram[3917] = 227;
    exp_33_ram[3918] = 131;
    exp_33_ram[3919] = 183;
    exp_33_ram[3920] = 19;
    exp_33_ram[3921] = 239;
    exp_33_ram[3922] = 19;
    exp_33_ram[3923] = 131;
    exp_33_ram[3924] = 3;
    exp_33_ram[3925] = 3;
    exp_33_ram[3926] = 131;
    exp_33_ram[3927] = 3;
    exp_33_ram[3928] = 131;
    exp_33_ram[3929] = 3;
    exp_33_ram[3930] = 131;
    exp_33_ram[3931] = 3;
    exp_33_ram[3932] = 131;
    exp_33_ram[3933] = 3;
    exp_33_ram[3934] = 131;
    exp_33_ram[3935] = 19;
    exp_33_ram[3936] = 103;
    exp_33_ram[3937] = 19;
    exp_33_ram[3938] = 35;
    exp_33_ram[3939] = 35;
    exp_33_ram[3940] = 35;
    exp_33_ram[3941] = 35;
    exp_33_ram[3942] = 35;
    exp_33_ram[3943] = 35;
    exp_33_ram[3944] = 19;
    exp_33_ram[3945] = 183;
    exp_33_ram[3946] = 19;
    exp_33_ram[3947] = 239;
    exp_33_ram[3948] = 239;
    exp_33_ram[3949] = 147;
    exp_33_ram[3950] = 147;
    exp_33_ram[3951] = 35;
    exp_33_ram[3952] = 183;
    exp_33_ram[3953] = 19;
    exp_33_ram[3954] = 239;
    exp_33_ram[3955] = 239;
    exp_33_ram[3956] = 147;
    exp_33_ram[3957] = 147;
    exp_33_ram[3958] = 35;
    exp_33_ram[3959] = 183;
    exp_33_ram[3960] = 19;
    exp_33_ram[3961] = 239;
    exp_33_ram[3962] = 239;
    exp_33_ram[3963] = 147;
    exp_33_ram[3964] = 35;
    exp_33_ram[3965] = 183;
    exp_33_ram[3966] = 19;
    exp_33_ram[3967] = 239;
    exp_33_ram[3968] = 239;
    exp_33_ram[3969] = 147;
    exp_33_ram[3970] = 35;
    exp_33_ram[3971] = 183;
    exp_33_ram[3972] = 19;
    exp_33_ram[3973] = 239;
    exp_33_ram[3974] = 239;
    exp_33_ram[3975] = 147;
    exp_33_ram[3976] = 35;
    exp_33_ram[3977] = 147;
    exp_33_ram[3978] = 35;
    exp_33_ram[3979] = 147;
    exp_33_ram[3980] = 35;
    exp_33_ram[3981] = 147;
    exp_33_ram[3982] = 19;
    exp_33_ram[3983] = 239;
    exp_33_ram[3984] = 19;
    exp_33_ram[3985] = 147;
    exp_33_ram[3986] = 35;
    exp_33_ram[3987] = 35;
    exp_33_ram[3988] = 147;
    exp_33_ram[3989] = 19;
    exp_33_ram[3990] = 239;
    exp_33_ram[3991] = 147;
    exp_33_ram[3992] = 19;
    exp_33_ram[3993] = 239;
    exp_33_ram[3994] = 147;
    exp_33_ram[3995] = 19;
    exp_33_ram[3996] = 239;
    exp_33_ram[3997] = 147;
    exp_33_ram[3998] = 19;
    exp_33_ram[3999] = 239;
    exp_33_ram[4000] = 3;
    exp_33_ram[4001] = 131;
    exp_33_ram[4002] = 19;
    exp_33_ram[4003] = 147;
    exp_33_ram[4004] = 239;
    exp_33_ram[4005] = 19;
    exp_33_ram[4006] = 239;
    exp_33_ram[4007] = 19;
    exp_33_ram[4008] = 147;
    exp_33_ram[4009] = 35;
    exp_33_ram[4010] = 35;
    exp_33_ram[4011] = 147;
    exp_33_ram[4012] = 19;
    exp_33_ram[4013] = 239;
    exp_33_ram[4014] = 147;
    exp_33_ram[4015] = 19;
    exp_33_ram[4016] = 239;
    exp_33_ram[4017] = 239;
    exp_33_ram[4018] = 35;
    exp_33_ram[4019] = 35;
    exp_33_ram[4020] = 35;
    exp_33_ram[4021] = 111;
    exp_33_ram[4022] = 19;
    exp_33_ram[4023] = 239;
    exp_33_ram[4024] = 19;
    exp_33_ram[4025] = 147;
    exp_33_ram[4026] = 3;
    exp_33_ram[4027] = 131;
    exp_33_ram[4028] = 19;
    exp_33_ram[4029] = 147;
    exp_33_ram[4030] = 239;
    exp_33_ram[4031] = 19;
    exp_33_ram[4032] = 147;
    exp_33_ram[4033] = 183;
    exp_33_ram[4034] = 131;
    exp_33_ram[4035] = 19;
    exp_33_ram[4036] = 239;
    exp_33_ram[4037] = 19;
    exp_33_ram[4038] = 147;
    exp_33_ram[4039] = 19;
    exp_33_ram[4040] = 147;
    exp_33_ram[4041] = 19;
    exp_33_ram[4042] = 147;
    exp_33_ram[4043] = 239;
    exp_33_ram[4044] = 147;
    exp_33_ram[4045] = 227;
    exp_33_ram[4046] = 183;
    exp_33_ram[4047] = 131;
    exp_33_ram[4048] = 19;
    exp_33_ram[4049] = 147;
    exp_33_ram[4050] = 3;
    exp_33_ram[4051] = 131;
    exp_33_ram[4052] = 51;
    exp_33_ram[4053] = 147;
    exp_33_ram[4054] = 179;
    exp_33_ram[4055] = 179;
    exp_33_ram[4056] = 179;
    exp_33_ram[4057] = 147;
    exp_33_ram[4058] = 35;
    exp_33_ram[4059] = 35;
    exp_33_ram[4060] = 19;
    exp_33_ram[4061] = 239;
    exp_33_ram[4062] = 19;
    exp_33_ram[4063] = 147;
    exp_33_ram[4064] = 35;
    exp_33_ram[4065] = 35;
    exp_33_ram[4066] = 147;
    exp_33_ram[4067] = 19;
    exp_33_ram[4068] = 239;
    exp_33_ram[4069] = 147;
    exp_33_ram[4070] = 19;
    exp_33_ram[4071] = 239;
    exp_33_ram[4072] = 131;
    exp_33_ram[4073] = 147;
    exp_33_ram[4074] = 35;
    exp_33_ram[4075] = 3;
    exp_33_ram[4076] = 147;
    exp_33_ram[4077] = 227;
    exp_33_ram[4078] = 19;
    exp_33_ram[4079] = 19;
    exp_33_ram[4080] = 131;
    exp_33_ram[4081] = 3;
    exp_33_ram[4082] = 3;
    exp_33_ram[4083] = 131;
    exp_33_ram[4084] = 3;
    exp_33_ram[4085] = 131;
    exp_33_ram[4086] = 19;
    exp_33_ram[4087] = 103;
    exp_33_ram[4088] = 19;
    exp_33_ram[4089] = 35;
    exp_33_ram[4090] = 35;
    exp_33_ram[4091] = 19;
    exp_33_ram[4092] = 183;
    exp_33_ram[4093] = 19;
    exp_33_ram[4094] = 239;
    exp_33_ram[4095] = 183;
    exp_33_ram[4096] = 19;
    exp_33_ram[4097] = 239;
    exp_33_ram[4098] = 183;
    exp_33_ram[4099] = 19;
    exp_33_ram[4100] = 239;
    exp_33_ram[4101] = 183;
    exp_33_ram[4102] = 19;
    exp_33_ram[4103] = 239;
    exp_33_ram[4104] = 183;
    exp_33_ram[4105] = 19;
    exp_33_ram[4106] = 239;
    exp_33_ram[4107] = 239;
    exp_33_ram[4108] = 147;
    exp_33_ram[4109] = 163;
    exp_33_ram[4110] = 131;
    exp_33_ram[4111] = 19;
    exp_33_ram[4112] = 99;
    exp_33_ram[4113] = 19;
    exp_33_ram[4114] = 227;
    exp_33_ram[4115] = 19;
    exp_33_ram[4116] = 99;
    exp_33_ram[4117] = 19;
    exp_33_ram[4118] = 227;
    exp_33_ram[4119] = 19;
    exp_33_ram[4120] = 99;
    exp_33_ram[4121] = 19;
    exp_33_ram[4122] = 99;
    exp_33_ram[4123] = 111;
    exp_33_ram[4124] = 239;
    exp_33_ram[4125] = 111;
    exp_33_ram[4126] = 239;
    exp_33_ram[4127] = 111;
    exp_33_ram[4128] = 239;
    exp_33_ram[4129] = 111;
    exp_33_ram[4130] = 239;
    exp_33_ram[4131] = 19;
    exp_33_ram[4132] = 111;
    exp_33_ram[4133] = 19;
    exp_33_ram[4134] = 147;
    exp_33_ram[4135] = 51;
    exp_33_ram[4136] = 19;
    exp_33_ram[4137] = 179;
    exp_33_ram[4138] = 99;
    exp_33_ram[4139] = 99;
    exp_33_ram[4140] = 19;
    exp_33_ram[4141] = 179;
    exp_33_ram[4142] = 19;
    exp_33_ram[4143] = 103;
    exp_33_ram[4144] = 227;
    exp_33_ram[4145] = 19;
    exp_33_ram[4146] = 179;
    exp_33_ram[4147] = 111;
    exp_33_ram[4148] = 128;
    exp_33_ram[4149] = 8;
    exp_33_ram[4150] = 12;
    exp_33_ram[4151] = 16;
    exp_33_ram[4152] = 40;
    exp_33_ram[4153] = 112;
    exp_33_ram[4154] = 112;
    exp_33_ram[4155] = 76;
    exp_33_ram[4156] = 112;
    exp_33_ram[4157] = 112;
    exp_33_ram[4158] = 112;
    exp_33_ram[4159] = 112;
    exp_33_ram[4160] = 112;
    exp_33_ram[4161] = 112;
    exp_33_ram[4162] = 112;
    exp_33_ram[4163] = 4;
    exp_33_ram[4164] = 112;
    exp_33_ram[4165] = 224;
    exp_33_ram[4166] = 112;
    exp_33_ram[4167] = 112;
    exp_33_ram[4168] = 188;
    exp_33_ram[4169] = 20;
    exp_33_ram[4170] = 172;
    exp_33_ram[4171] = 116;
    exp_33_ram[4172] = 172;
    exp_33_ram[4173] = 208;
    exp_33_ram[4174] = 172;
    exp_33_ram[4175] = 172;
    exp_33_ram[4176] = 172;
    exp_33_ram[4177] = 172;
    exp_33_ram[4178] = 172;
    exp_33_ram[4179] = 172;
    exp_33_ram[4180] = 172;
    exp_33_ram[4181] = 88;
    exp_33_ram[4182] = 172;
    exp_33_ram[4183] = 172;
    exp_33_ram[4184] = 172;
    exp_33_ram[4185] = 172;
    exp_33_ram[4186] = 172;
    exp_33_ram[4187] = 144;
    exp_33_ram[4188] = 212;
    exp_33_ram[4189] = 8;
    exp_33_ram[4190] = 8;
    exp_33_ram[4191] = 8;
    exp_33_ram[4192] = 8;
    exp_33_ram[4193] = 8;
    exp_33_ram[4194] = 8;
    exp_33_ram[4195] = 8;
    exp_33_ram[4196] = 8;
    exp_33_ram[4197] = 8;
    exp_33_ram[4198] = 8;
    exp_33_ram[4199] = 8;
    exp_33_ram[4200] = 8;
    exp_33_ram[4201] = 8;
    exp_33_ram[4202] = 8;
    exp_33_ram[4203] = 8;
    exp_33_ram[4204] = 8;
    exp_33_ram[4205] = 8;
    exp_33_ram[4206] = 8;
    exp_33_ram[4207] = 8;
    exp_33_ram[4208] = 8;
    exp_33_ram[4209] = 8;
    exp_33_ram[4210] = 8;
    exp_33_ram[4211] = 8;
    exp_33_ram[4212] = 8;
    exp_33_ram[4213] = 8;
    exp_33_ram[4214] = 8;
    exp_33_ram[4215] = 8;
    exp_33_ram[4216] = 8;
    exp_33_ram[4217] = 8;
    exp_33_ram[4218] = 8;
    exp_33_ram[4219] = 8;
    exp_33_ram[4220] = 8;
    exp_33_ram[4221] = 8;
    exp_33_ram[4222] = 8;
    exp_33_ram[4223] = 8;
    exp_33_ram[4224] = 8;
    exp_33_ram[4225] = 8;
    exp_33_ram[4226] = 8;
    exp_33_ram[4227] = 8;
    exp_33_ram[4228] = 8;
    exp_33_ram[4229] = 8;
    exp_33_ram[4230] = 8;
    exp_33_ram[4231] = 8;
    exp_33_ram[4232] = 8;
    exp_33_ram[4233] = 8;
    exp_33_ram[4234] = 8;
    exp_33_ram[4235] = 8;
    exp_33_ram[4236] = 8;
    exp_33_ram[4237] = 8;
    exp_33_ram[4238] = 8;
    exp_33_ram[4239] = 236;
    exp_33_ram[4240] = 8;
    exp_33_ram[4241] = 8;
    exp_33_ram[4242] = 8;
    exp_33_ram[4243] = 8;
    exp_33_ram[4244] = 8;
    exp_33_ram[4245] = 8;
    exp_33_ram[4246] = 8;
    exp_33_ram[4247] = 8;
    exp_33_ram[4248] = 8;
    exp_33_ram[4249] = 236;
    exp_33_ram[4250] = 56;
    exp_33_ram[4251] = 236;
    exp_33_ram[4252] = 8;
    exp_33_ram[4253] = 8;
    exp_33_ram[4254] = 8;
    exp_33_ram[4255] = 8;
    exp_33_ram[4256] = 236;
    exp_33_ram[4257] = 8;
    exp_33_ram[4258] = 8;
    exp_33_ram[4259] = 8;
    exp_33_ram[4260] = 8;
    exp_33_ram[4261] = 8;
    exp_33_ram[4262] = 236;
    exp_33_ram[4263] = 104;
    exp_33_ram[4264] = 8;
    exp_33_ram[4265] = 8;
    exp_33_ram[4266] = 20;
    exp_33_ram[4267] = 8;
    exp_33_ram[4268] = 236;
    exp_33_ram[4269] = 8;
    exp_33_ram[4270] = 8;
    exp_33_ram[4271] = 236;
    exp_33_ram[4272] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_179;

  reg [31:0] exp_179_reg;
  always@(*) begin
    case (exp_177)
      0:exp_179_reg <= exp_157;
      1:exp_179_reg <= exp_167;
      default:exp_179_reg <= exp_178;
    endcase
  end
  assign exp_179 = exp_179_reg;
  assign exp_177 = exp_139[2:2];
  assign exp_139 = exp_1;
  assign exp_178 = 0;

      reg [31:0] exp_157_reg = 0;
      always@(posedge clk) begin
        if (exp_156) begin
          exp_157_reg <= exp_164;
        end
      end
      assign exp_157 = exp_157_reg;
    
  reg [31:0] exp_164_reg;
  always@(*) begin
    case (exp_159)
      0:exp_164_reg <= exp_161;
      1:exp_164_reg <= exp_162;
      default:exp_164_reg <= exp_163;
    endcase
  end
  assign exp_164 = exp_164_reg;
  assign exp_159 = exp_157 == exp_158;
  assign exp_158 = 4294967295;
  assign exp_163 = 0;
  assign exp_161 = exp_157 + exp_160;
  assign exp_160 = 1;
  assign exp_162 = 0;
  assign exp_156 = 1;

      reg [31:0] exp_167_reg = 0;
      always@(posedge clk) begin
        if (exp_166) begin
          exp_167_reg <= exp_174;
        end
      end
      assign exp_167 = exp_167_reg;
    
  reg [31:0] exp_174_reg;
  always@(*) begin
    case (exp_169)
      0:exp_174_reg <= exp_171;
      1:exp_174_reg <= exp_172;
      default:exp_174_reg <= exp_173;
    endcase
  end
  assign exp_174 = exp_174_reg;
  assign exp_169 = exp_167 == exp_168;
  assign exp_168 = 4294967295;
  assign exp_173 = 0;
  assign exp_171 = exp_167 + exp_170;
  assign exp_170 = 1;
  assign exp_172 = 0;
  assign exp_166 = exp_159 & exp_165;
  assign exp_165 = 1;
  assign exp_182 = exp_281;
  assign exp_281 = 0;
  assign exp_284 = exp_302;
  assign exp_302 = 0;
  assign exp_307 = exp_391;
  assign exp_391 = exp_388;

      reg [7:0] exp_388_reg = 0;
      always@(posedge clk) begin
        if (exp_387) begin
          exp_388_reg <= exp_390;
        end
      end
      assign exp_388 = exp_388_reg;
      assign exp_390 = {exp_329, exp_389};  assign exp_389 = exp_388[7:1];
  assign exp_387 = exp_352 & exp_386;
  assign exp_386 = exp_353 == exp_385;
  assign exp_385 = 0;
  assign exp_607 = exp_394[15:8];
  assign exp_608 = exp_394[23:16];
  assign exp_609 = exp_394[31:24];
  assign exp_621 = $signed(exp_620);
  assign exp_620 = exp_619 + exp_615;
  assign exp_619 = 0;

  reg [15:0] exp_615_reg;
  always@(*) begin
    case (exp_605)
      0:exp_615_reg <= exp_612;
      1:exp_615_reg <= exp_613;
      default:exp_615_reg <= exp_614;
    endcase
  end
  assign exp_615 = exp_615_reg;
  assign exp_614 = 0;
  assign exp_612 = exp_394[15:0];
  assign exp_613 = exp_394[31:16];
  assign exp_622 = 0;
  assign exp_623 = exp_611;
  assign exp_624 = exp_615;
  assign exp_625 = 0;
  assign exp_626 = 0;

  reg [31:0] exp_985_reg;
  always@(*) begin
    case (exp_775)
      0:exp_985_reg <= exp_981;
      1:exp_985_reg <= exp_983;
      default:exp_985_reg <= exp_984;
    endcase
  end
  assign exp_985 = exp_985_reg;
  assign exp_984 = 0;

  reg [31:0] exp_981_reg;
  always@(*) begin
    case (exp_752)
      0:exp_981_reg <= exp_976;
      1:exp_981_reg <= exp_977;
      default:exp_981_reg <= exp_980;
    endcase
  end
  assign exp_981 = exp_981_reg;
  assign exp_752 = exp_751 & exp_749;
  assign exp_751 = exp_744 == exp_750;
  assign exp_750 = 0;
  assign exp_980 = 0;
  assign exp_976 = exp_975[63:32];

  reg [63:0] exp_975_reg;
  always@(*) begin
    case (exp_972)
      0:exp_975_reg <= exp_971;
      1:exp_975_reg <= exp_973;
      default:exp_975_reg <= exp_974;
    endcase
  end
  assign exp_975 = exp_975_reg;

      reg [0:0] exp_972_reg = 0;
      always@(posedge clk) begin
        if (exp_957) begin
          exp_972_reg <= exp_955;
        end
      end
      assign exp_972 = exp_972_reg;
    
      reg [0:0] exp_955_reg = 0;
      always@(posedge clk) begin
        if (exp_934) begin
          exp_955_reg <= exp_932;
        end
      end
      assign exp_955 = exp_955_reg;
    
      reg [0:0] exp_932_reg = 0;
      always@(posedge clk) begin
        if (exp_914) begin
          exp_932_reg <= exp_929;
        end
      end
      assign exp_932 = exp_932_reg;
      assign exp_929 = exp_927 ^ exp_928;
  assign exp_927 = exp_909 & exp_892;
  assign exp_909 = exp_908 + exp_907;
  assign exp_908 = 0;
  assign exp_907 = exp_905[31:31];

      reg [31:0] exp_905_reg = 0;
      always@(posedge clk) begin
        if (exp_904) begin
          exp_905_reg <= exp_522;
        end
      end
      assign exp_905 = exp_905_reg;
      assign exp_904 = exp_894 == exp_903;
  assign exp_903 = 0;
  assign exp_892 = exp_891 | exp_758;
  assign exp_891 = exp_752 | exp_755;
  assign exp_755 = exp_754 & exp_749;
  assign exp_754 = exp_744 == exp_753;
  assign exp_753 = 1;
  assign exp_758 = exp_757 & exp_749;
  assign exp_757 = exp_744 == exp_756;
  assign exp_756 = 2;
  assign exp_928 = exp_912 & exp_893;
  assign exp_912 = exp_911 + exp_910;
  assign exp_911 = 0;
  assign exp_910 = exp_906[31:31];

      reg [31:0] exp_906_reg = 0;
      always@(posedge clk) begin
        if (exp_904) begin
          exp_906_reg <= exp_523;
        end
      end
      assign exp_906 = exp_906_reg;
      assign exp_893 = exp_752 | exp_755;
  assign exp_914 = exp_894 == exp_913;
  assign exp_913 = 1;
  assign exp_934 = exp_894 == exp_933;
  assign exp_933 = 2;
  assign exp_957 = exp_894 == exp_956;
  assign exp_956 = 3;
  assign exp_974 = 0;

      reg [63:0] exp_971_reg = 0;
      always@(posedge clk) begin
        if (exp_957) begin
          exp_971_reg <= exp_970;
        end
      end
      assign exp_971 = exp_971_reg;
      assign exp_970 = exp_966 + exp_969;
  assign exp_966 = exp_962 + exp_965;
  assign exp_962 = exp_958 + exp_961;
  assign exp_958 = exp_951;

      reg [31:0] exp_951_reg = 0;
      always@(posedge clk) begin
        if (exp_934) begin
          exp_951_reg <= exp_938;
        end
      end
      assign exp_951 = exp_951_reg;
      assign exp_938 = exp_936 * exp_937;
  assign exp_936 = exp_935;
  assign exp_935 = exp_930[15:0];

      reg [31:0] exp_930_reg = 0;
      always@(posedge clk) begin
        if (exp_914) begin
          exp_930_reg <= exp_920;
        end
      end
      assign exp_930 = exp_930_reg;
      assign exp_920 = exp_919 + exp_918;
  assign exp_919 = 0;

  reg [31:0] exp_918_reg;
  always@(*) begin
    case (exp_915)
      0:exp_918_reg <= exp_905;
      1:exp_918_reg <= exp_916;
      default:exp_918_reg <= exp_917;
    endcase
  end
  assign exp_918 = exp_918_reg;
  assign exp_915 = exp_909 & exp_892;
  assign exp_917 = 0;
  assign exp_916 = -exp_905;
  assign exp_937 = exp_931[15:0];

      reg [31:0] exp_931_reg = 0;
      always@(posedge clk) begin
        if (exp_914) begin
          exp_931_reg <= exp_926;
        end
      end
      assign exp_931 = exp_931_reg;
      assign exp_926 = exp_925 + exp_924;
  assign exp_925 = 0;

  reg [31:0] exp_924_reg;
  always@(*) begin
    case (exp_921)
      0:exp_924_reg <= exp_906;
      1:exp_924_reg <= exp_922;
      default:exp_924_reg <= exp_923;
    endcase
  end
  assign exp_924 = exp_924_reg;
  assign exp_921 = exp_912 & exp_893;
  assign exp_923 = 0;
  assign exp_922 = -exp_906;
  assign exp_961 = exp_959 << exp_960;
  assign exp_959 = exp_952;

      reg [31:0] exp_952_reg = 0;
      always@(posedge clk) begin
        if (exp_934) begin
          exp_952_reg <= exp_942;
        end
      end
      assign exp_952 = exp_952_reg;
      assign exp_942 = exp_940 * exp_941;
  assign exp_940 = exp_939;
  assign exp_939 = exp_930[15:0];
  assign exp_941 = exp_931[31:16];
  assign exp_960 = 16;
  assign exp_965 = exp_963 << exp_964;
  assign exp_963 = exp_953;

      reg [31:0] exp_953_reg = 0;
      always@(posedge clk) begin
        if (exp_934) begin
          exp_953_reg <= exp_946;
        end
      end
      assign exp_953 = exp_953_reg;
      assign exp_946 = exp_944 * exp_945;
  assign exp_944 = exp_943;
  assign exp_943 = exp_930[31:16];
  assign exp_945 = exp_931[15:0];
  assign exp_964 = 16;
  assign exp_969 = exp_967 << exp_968;
  assign exp_967 = exp_954;

      reg [31:0] exp_954_reg = 0;
      always@(posedge clk) begin
        if (exp_934) begin
          exp_954_reg <= exp_950;
        end
      end
      assign exp_954 = exp_954_reg;
      assign exp_950 = exp_948 * exp_949;
  assign exp_948 = exp_947;
  assign exp_947 = exp_930[31:16];
  assign exp_949 = exp_931[31:16];
  assign exp_968 = 32;
  assign exp_973 = -exp_971;
  assign exp_977 = exp_975[31:0];

  reg [31:0] exp_983_reg;
  always@(*) begin
    case (exp_776)
      0:exp_983_reg <= exp_886;
      1:exp_983_reg <= exp_887;
      default:exp_983_reg <= exp_982;
    endcase
  end
  assign exp_983 = exp_983_reg;
  assign exp_776 = exp_744[1:1];
  assign exp_982 = 0;

      reg [31:0] exp_886_reg = 0;
      always@(posedge clk) begin
        if (exp_795) begin
          exp_886_reg <= exp_880;
        end
      end
      assign exp_886 = exp_886_reg;
    
  reg [31:0] exp_880_reg;
  always@(*) begin
    case (exp_876)
      0:exp_880_reg <= exp_867;
      1:exp_880_reg <= exp_878;
      default:exp_880_reg <= exp_879;
    endcase
  end
  assign exp_880 = exp_880_reg;
  assign exp_876 = exp_875 & exp_778;
  assign exp_875 = exp_824 == exp_874;

      reg [31:0] exp_824_reg = 0;
      always@(posedge clk) begin
        if (exp_809) begin
          exp_824_reg <= exp_821;
        end
      end
      assign exp_824 = exp_824_reg;
      assign exp_821 = exp_820 + exp_819;
  assign exp_820 = 0;

  reg [31:0] exp_819_reg;
  always@(*) begin
    case (exp_816)
      0:exp_819_reg <= exp_801;
      1:exp_819_reg <= exp_817;
      default:exp_819_reg <= exp_818;
    endcase
  end
  assign exp_819 = exp_819_reg;
  assign exp_816 = exp_807 & exp_778;
  assign exp_807 = exp_806 + exp_805;
  assign exp_806 = 0;
  assign exp_805 = exp_801[31:31];

      reg [31:0] exp_801_reg = 0;
      always@(posedge clk) begin
        if (exp_799) begin
          exp_801_reg <= exp_523;
        end
      end
      assign exp_801 = exp_801_reg;
      assign exp_799 = exp_781 == exp_798;
  assign exp_798 = 0;
  assign exp_778 = ~exp_777;
  assign exp_777 = exp_744[0:0];
  assign exp_818 = 0;
  assign exp_817 = -exp_801;
  assign exp_809 = exp_781 == exp_808;
  assign exp_808 = 1;
  assign exp_874 = 0;
  assign exp_879 = 0;
  assign exp_867 = exp_866 + exp_865;
  assign exp_866 = 0;

  reg [31:0] exp_865_reg;
  always@(*) begin
    case (exp_862)
      0:exp_865_reg <= exp_860;
      1:exp_865_reg <= exp_863;
      default:exp_865_reg <= exp_864;
    endcase
  end
  assign exp_865 = exp_865_reg;
  assign exp_862 = exp_826 & exp_778;

      reg [0:0] exp_826_reg = 0;
      always@(posedge clk) begin
        if (exp_809) begin
          exp_826_reg <= exp_822;
        end
      end
      assign exp_826 = exp_826_reg;
      assign exp_822 = exp_804 ^ exp_807;
  assign exp_804 = exp_803 + exp_802;
  assign exp_803 = 0;
  assign exp_802 = exp_800[31:31];

      reg [31:0] exp_800_reg = 0;
      always@(posedge clk) begin
        if (exp_799) begin
          exp_800_reg <= exp_522;
        end
      end
      assign exp_800 = exp_800_reg;
      assign exp_864 = 0;

      reg [31:0] exp_860_reg = 0;
      always@(posedge clk) begin
        if (exp_793) begin
          exp_860_reg <= exp_830;
        end
      end
      assign exp_860 = exp_860_reg;
    
      reg [31:0] exp_830_reg = 0;
      always@(posedge clk) begin
        if (exp_829) begin
          exp_830_reg <= exp_857;
        end
      end
      assign exp_830 = exp_830_reg;
    
  reg [31:0] exp_857_reg;
  always@(*) begin
    case (exp_791)
      0:exp_857_reg <= exp_849;
      1:exp_857_reg <= exp_855;
      default:exp_857_reg <= exp_856;
    endcase
  end
  assign exp_857 = exp_857_reg;
  assign exp_791 = exp_781 == exp_790;
  assign exp_790 = 2;
  assign exp_856 = 0;

  reg [31:0] exp_849_reg;
  always@(*) begin
    case (exp_839)
      0:exp_849_reg <= exp_843;
      1:exp_849_reg <= exp_847;
      default:exp_849_reg <= exp_848;
    endcase
  end
  assign exp_849 = exp_849_reg;
  assign exp_839 = ~exp_838;
  assign exp_838 = exp_837[32:32];
  assign exp_837 = exp_836 - exp_824;
  assign exp_836 = exp_835;
  assign exp_835 = {exp_833, exp_834};  assign exp_833 = exp_828[31:0];

      reg [31:0] exp_828_reg = 0;
      always@(posedge clk) begin
        if (exp_827) begin
          exp_828_reg <= exp_854;
        end
      end
      assign exp_828 = exp_828_reg;
    
  reg [32:0] exp_854_reg;
  always@(*) begin
    case (exp_791)
      0:exp_854_reg <= exp_841;
      1:exp_854_reg <= exp_852;
      default:exp_854_reg <= exp_853;
    endcase
  end
  assign exp_854 = exp_854_reg;
  assign exp_853 = 0;

  reg [32:0] exp_841_reg;
  always@(*) begin
    case (exp_839)
      0:exp_841_reg <= exp_835;
      1:exp_841_reg <= exp_837;
      default:exp_841_reg <= exp_840;
    endcase
  end
  assign exp_841 = exp_841_reg;
  assign exp_840 = 0;
  assign exp_852 = 0;
  assign exp_827 = 1;
  assign exp_834 = exp_832[31:31];

      reg [31:0] exp_832_reg = 0;
      always@(posedge clk) begin
        if (exp_831) begin
          exp_832_reg <= exp_859;
        end
      end
      assign exp_832 = exp_832_reg;
    
  reg [31:0] exp_859_reg;
  always@(*) begin
    case (exp_791)
      0:exp_859_reg <= exp_851;
      1:exp_859_reg <= exp_823;
      default:exp_859_reg <= exp_858;
    endcase
  end
  assign exp_859 = exp_859_reg;
  assign exp_858 = 0;
  assign exp_851 = exp_832 << exp_850;
  assign exp_850 = 1;

      reg [31:0] exp_823_reg = 0;
      always@(posedge clk) begin
        if (exp_809) begin
          exp_823_reg <= exp_815;
        end
      end
      assign exp_823 = exp_823_reg;
      assign exp_815 = exp_814 + exp_813;
  assign exp_814 = 0;

  reg [31:0] exp_813_reg;
  always@(*) begin
    case (exp_810)
      0:exp_813_reg <= exp_800;
      1:exp_813_reg <= exp_811;
      default:exp_813_reg <= exp_812;
    endcase
  end
  assign exp_813 = exp_813_reg;
  assign exp_810 = exp_804 & exp_778;
  assign exp_812 = 0;
  assign exp_811 = -exp_800;
  assign exp_831 = 1;
  assign exp_848 = 0;
  assign exp_843 = exp_830 << exp_842;
  assign exp_842 = 1;
  assign exp_847 = exp_845 | exp_846;
  assign exp_845 = exp_830 << exp_844;
  assign exp_844 = 1;
  assign exp_846 = 1;
  assign exp_855 = 0;
  assign exp_829 = 1;
  assign exp_793 = exp_781 == exp_792;
  assign exp_792 = 35;
  assign exp_863 = -exp_860;
  assign exp_878 = $signed(exp_877);
  assign exp_877 = -1;
  assign exp_795 = exp_781 == exp_794;
  assign exp_794 = 36;

      reg [31:0] exp_887_reg = 0;
      always@(posedge clk) begin
        if (exp_795) begin
          exp_887_reg <= exp_885;
        end
      end
      assign exp_887 = exp_887_reg;
    
  reg [31:0] exp_885_reg;
  always@(*) begin
    case (exp_883)
      0:exp_885_reg <= exp_873;
      1:exp_885_reg <= exp_800;
      default:exp_885_reg <= exp_884;
    endcase
  end
  assign exp_885 = exp_885_reg;
  assign exp_883 = exp_882 & exp_778;
  assign exp_882 = exp_824 == exp_881;
  assign exp_881 = 0;
  assign exp_884 = 0;
  assign exp_873 = exp_872 + exp_871;
  assign exp_872 = 0;

  reg [31:0] exp_871_reg;
  always@(*) begin
    case (exp_868)
      0:exp_871_reg <= exp_861;
      1:exp_871_reg <= exp_869;
      default:exp_871_reg <= exp_870;
    endcase
  end
  assign exp_871 = exp_871_reg;
  assign exp_868 = exp_825 & exp_778;

      reg [0:0] exp_825_reg = 0;
      always@(posedge clk) begin
        if (exp_809) begin
          exp_825_reg <= exp_804;
        end
      end
      assign exp_825 = exp_825_reg;
      assign exp_870 = 0;

      reg [31:0] exp_861_reg = 0;
      always@(posedge clk) begin
        if (exp_793) begin
          exp_861_reg <= exp_828;
        end
      end
      assign exp_861 = exp_861_reg;
      assign exp_869 = -exp_861;
  assign exp_456 = $signed(exp_455);
  assign exp_455 = 0;
  assign exp_685 = exp_520 != exp_521;
  assign exp_698 = 0;
  assign exp_699 = 0;
  assign exp_686 = $signed(exp_520) < $signed(exp_521);
  assign exp_687 = $signed(exp_520) >= $signed(exp_521);
  assign exp_692 = exp_689 < exp_691;
  assign exp_689 = exp_688 + exp_520;
  assign exp_688 = 0;
  assign exp_691 = exp_690 + exp_521;
  assign exp_690 = 0;
  assign exp_697 = exp_694 >= exp_696;
  assign exp_694 = exp_693 + exp_520;
  assign exp_693 = 0;
  assign exp_696 = exp_695 + exp_521;
  assign exp_695 = 0;
  assign exp_1012 = 0;
  assign exp_1011 = exp_410 + exp_1010;
  assign exp_1010 = 4;

  reg [32:0] exp_742_reg;
  always@(*) begin
    case (exp_543)
      0:exp_742_reg <= exp_732;
      1:exp_742_reg <= exp_740;
      default:exp_742_reg <= exp_741;
    endcase
  end
  assign exp_742 = exp_742_reg;
  assign exp_741 = 0;
  assign exp_732 = exp_731 + exp_529;

  reg [31:0] exp_731_reg;
  always@(*) begin
    case (exp_541)
      0:exp_731_reg <= exp_717;
      1:exp_731_reg <= exp_729;
      default:exp_731_reg <= exp_730;
    endcase
  end
  assign exp_731 = exp_731_reg;
  assign exp_730 = 0;
  assign exp_717 = $signed(exp_716);
  assign exp_716 = exp_715 + exp_714;
  assign exp_715 = 0;
  assign exp_714 = {exp_713, exp_710};  assign exp_713 = {exp_712, exp_709};  assign exp_712 = {exp_711, exp_708};  assign exp_711 = {exp_706, exp_707};  assign exp_706 = exp_528[31:31];
  assign exp_707 = exp_528[7:7];
  assign exp_708 = exp_528[30:25];
  assign exp_709 = exp_528[11:8];
  assign exp_710 = 0;
  assign exp_729 = $signed(exp_728);
  assign exp_728 = exp_727 + exp_726;
  assign exp_727 = 0;
  assign exp_726 = {exp_725, exp_722};  assign exp_725 = {exp_724, exp_721};  assign exp_724 = {exp_723, exp_720};  assign exp_723 = {exp_718, exp_719};  assign exp_718 = exp_528[31:31];
  assign exp_719 = exp_528[19:12];
  assign exp_720 = exp_528[20:20];
  assign exp_721 = exp_528[30:21];
  assign exp_722 = 0;

      reg [31:0] exp_529_reg = 0;
      always@(posedge clk) begin
        if (exp_519) begin
          exp_529_reg <= exp_412;
        end
      end
      assign exp_529 = exp_529_reg;
      assign exp_740 = exp_739 & exp_738;
  assign exp_739 = $signed(exp_737);
  assign exp_737 = exp_520 + exp_736;
  assign exp_736 = $signed(exp_735);
  assign exp_735 = exp_734 + exp_733;
  assign exp_734 = 0;
  assign exp_733 = exp_528[31:20];
  assign exp_738 = 4294967294;
  assign exp_409 = exp_402 & exp_400;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_411;
  assign exp_544 = 3;
  assign exp_185 = exp_6;
  assign exp_218 = exp_206 & exp_217;
  assign exp_217 = ~exp_215;
  assign exp_215 = exp_209 & exp_206;
  assign exp_209 = exp_207 == exp_208;

      reg [8:0] exp_207_reg = 0;
      always@(posedge clk) begin
        if (exp_206) begin
          exp_207_reg <= exp_214;
        end
      end
      assign exp_207 = exp_207_reg;
    
  reg [8:0] exp_214_reg;
  always@(*) begin
    case (exp_209)
      0:exp_214_reg <= exp_211;
      1:exp_214_reg <= exp_212;
      default:exp_214_reg <= exp_213;
    endcase
  end
  assign exp_214 = exp_214_reg;
  assign exp_213 = 0;
  assign exp_211 = exp_207 + exp_210;
  assign exp_210 = 1;
  assign exp_212 = 0;
  assign exp_208 = 433;
  assign exp_205 = 1;
  assign exp_244 = exp_221 & exp_243;
  assign exp_243 = ~exp_242;
  assign exp_242 = exp_230 & exp_240;
  assign exp_230 = exp_224 & exp_221;
  assign exp_224 = exp_222 == exp_223;

      reg [8:0] exp_222_reg = 0;
      always@(posedge clk) begin
        if (exp_221) begin
          exp_222_reg <= exp_229;
        end
      end
      assign exp_222 = exp_222_reg;
    
  reg [8:0] exp_229_reg;
  always@(*) begin
    case (exp_224)
      0:exp_229_reg <= exp_226;
      1:exp_229_reg <= exp_227;
      default:exp_229_reg <= exp_228;
    endcase
  end
  assign exp_229 = exp_229_reg;
  assign exp_228 = 0;
  assign exp_226 = exp_222 + exp_225;
  assign exp_225 = 1;
  assign exp_227 = 0;
  assign exp_223 = 433;
  assign exp_240 = exp_234 & exp_231;
  assign exp_234 = exp_232 == exp_233;

      reg [2:0] exp_232_reg = 0;
      always@(posedge clk) begin
        if (exp_231) begin
          exp_232_reg <= exp_239;
        end
      end
      assign exp_232 = exp_232_reg;
    
  reg [2:0] exp_239_reg;
  always@(*) begin
    case (exp_234)
      0:exp_239_reg <= exp_236;
      1:exp_239_reg <= exp_237;
      default:exp_239_reg <= exp_238;
    endcase
  end
  assign exp_239 = exp_239_reg;
  assign exp_238 = 0;
  assign exp_236 = exp_232 + exp_235;
  assign exp_235 = 1;
  assign exp_237 = 0;
  assign exp_231 = exp_221 & exp_230;
  assign exp_233 = 7;
  assign exp_220 = 1;
  assign exp_260 = exp_247 & exp_259;
  assign exp_259 = ~exp_256;
  assign exp_256 = exp_250 & exp_247;
  assign exp_250 = exp_248 == exp_249;

      reg [8:0] exp_248_reg = 0;
      always@(posedge clk) begin
        if (exp_247) begin
          exp_248_reg <= exp_255;
        end
      end
      assign exp_248 = exp_248_reg;
    
  reg [8:0] exp_255_reg;
  always@(*) begin
    case (exp_250)
      0:exp_255_reg <= exp_252;
      1:exp_255_reg <= exp_253;
      default:exp_255_reg <= exp_254;
    endcase
  end
  assign exp_255 = exp_255_reg;
  assign exp_254 = 0;
  assign exp_252 = exp_248 + exp_251;
  assign exp_251 = 1;
  assign exp_253 = 0;
  assign exp_249 = 433;
  assign exp_246 = 1;
  assign exp_203 = exp_201 & exp_202;
  assign exp_202 = ~exp_198;
  assign exp_200 = 1;
  assign exp_279 = 0;

  reg [0:0] exp_276_reg;
  always@(*) begin
    case (exp_206)
      0:exp_276_reg <= exp_273;
      1:exp_276_reg <= exp_274;
      default:exp_276_reg <= exp_275;
    endcase
  end
  assign exp_276 = exp_276_reg;
  assign exp_275 = 0;
  assign exp_273 = exp_264[0:0];

      reg [7:0] exp_264_reg = 0;
      always@(posedge clk) begin
        if (exp_263) begin
          exp_264_reg <= exp_272;
        end
      end
      assign exp_264 = exp_264_reg;
    
  reg [7:0] exp_272_reg;
  always@(*) begin
    case (exp_270)
      0:exp_272_reg <= exp_269;
      1:exp_272_reg <= exp_197;
      default:exp_272_reg <= exp_271;
    endcase
  end
  assign exp_272 = exp_272_reg;
  assign exp_270 = exp_201 & exp_198;
  assign exp_271 = 0;

  reg [7:0] exp_269_reg;
  always@(*) begin
    case (exp_265)
      0:exp_269_reg <= exp_264;
      1:exp_269_reg <= exp_267;
      default:exp_269_reg <= exp_268;
    endcase
  end
  assign exp_269 = exp_269_reg;
  assign exp_265 = exp_221 & exp_230;
  assign exp_268 = 0;
  assign exp_267 = exp_264 >> exp_266;
  assign exp_266 = 1;
  assign exp_197 = exp_181[7:0];
  assign exp_181 = exp_2;
  assign exp_263 = 1;
  assign exp_274 = 0;
  assign exp_278 = 1;

      reg [31:0] exp_301_reg = 0;
      always@(posedge clk) begin
        if (exp_300) begin
          exp_301_reg <= exp_283;
        end
      end
      assign exp_301 = exp_301_reg;
      assign exp_283 = exp_2;
  assign exp_300 = exp_286 & exp_287;
  assign exp_286 = exp_294;
  assign exp_294 = exp_5 & exp_293;
  assign exp_287 = exp_6;
  assign stdout_tx = exp_280;
  assign leds_out = exp_301;

endmodule