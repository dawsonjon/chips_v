
module blink(clk, stdin_valid_in, stdin_in, buttons_rx, stdout_ready_in, stdin_ready_out, stdout_valid_out, stdout_out, leds_tx);
  input [0:0] stdin_valid_in;
  input [31:0] stdin_in;
  input [0:0] buttons_rx;
  input [0:0] stdout_ready_in;
  input [0:0] clk;
  output [0:0] stdin_ready_out;
  output [0:0] stdout_valid_out;
  output [31:0] stdout_out;
  output [0:0] leds_tx;
  wire [0:0] exp_324;
  wire [0:0] exp_307;
  wire [0:0] exp_315;
  wire [0:0] exp_5;
  wire [0:0] exp_410;
  wire [0:0] exp_757;
  wire [0:0] exp_694;
  wire [0:0] exp_559;
  wire [6:0] exp_544;
  wire [31:0] exp_542;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [10:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_424;
  wire [32:0] exp_1027;
  wire [0:0] exp_1023;
  wire [0:0] exp_719;
  wire [0:0] exp_697;
  wire [0:0] exp_555;
  wire [6:0] exp_554;
  wire [0:0] exp_557;
  wire [6:0] exp_556;
  wire [0:0] exp_718;
  wire [0:0] exp_563;
  wire [6:0] exp_562;
  wire [0:0] exp_717;
  wire [0:0] exp_716;
  wire [0:0] exp_715;
  wire [2:0] exp_545;
  wire [0:0] exp_714;
  wire [0:0] exp_698;
  wire [31:0] exp_534;
  wire [31:0] exp_472;
  wire [0:0] exp_468;
  wire [4:0] exp_448;
  wire [0:0] exp_467;
  wire [0:0] exp_471;
  wire [31:0] exp_464;
  wire [0:0] exp_445;
  wire [0:0] exp_1018;
  wire [0:0] exp_1017;
  wire [0:0] exp_1016;
  wire [0:0] exp_1015;
  wire [4:0] exp_427;
  wire [4:0] exp_1010;
  wire [0:0] exp_1009;
  wire [0:0] exp_601;
  wire [0:0] exp_600;
  wire [0:0] exp_599;
  wire [0:0] exp_598;
  wire [0:0] exp_597;
  wire [0:0] exp_596;
  wire [0:0] exp_547;
  wire [4:0] exp_546;
  wire [0:0] exp_549;
  wire [5:0] exp_548;
  wire [0:0] exp_551;
  wire [5:0] exp_550;
  wire [0:0] exp_553;
  wire [4:0] exp_552;
  wire [0:0] exp_1004;
  wire [0:0] exp_1003;
  wire [0:0] exp_789;
  wire [0:0] exp_763;
  wire [0:0] exp_761;
  wire [6:0] exp_759;
  wire [5:0] exp_760;
  wire [0:0] exp_762;
  wire [0:0] exp_788;
  wire [2:0] exp_758;
  wire [0:0] exp_1002;
  wire [0:0] exp_1000;
  wire [0:0] exp_993;
  wire [2:0] exp_908;
  wire [2:0] exp_915;
  wire [0:0] exp_910;
  wire [2:0] exp_909;
  wire [0:0] exp_914;
  wire [2:0] exp_912;
  wire [0:0] exp_911;
  wire [0:0] exp_913;
  wire [0:0] exp_904;
  wire [0:0] exp_903;
  wire [0:0] exp_902;
  wire [2:0] exp_992;
  wire [0:0] exp_1001;
  wire [0:0] exp_811;
  wire [5:0] exp_795;
  wire [5:0] exp_802;
  wire [0:0] exp_797;
  wire [5:0] exp_796;
  wire [0:0] exp_801;
  wire [5:0] exp_799;
  wire [0:0] exp_798;
  wire [0:0] exp_800;
  wire [5:0] exp_810;
  wire [0:0] exp_422;
  wire [0:0] exp_421;
  wire [0:0] exp_419;
  wire [0:0] exp_418;
  wire [0:0] exp_416;
  wire [0:0] exp_417;
  wire [0:0] exp_415;
  wire [0:0] exp_1028;
  wire [0:0] exp_414;
  wire [0:0] exp_413;
  wire [0:0] exp_1032;
  wire [0:0] exp_1031;
  wire [0:0] exp_1030;
  wire [0:0] exp_1029;
  wire [0:0] exp_409;
  wire [0:0] exp_342;
  wire [0:0] exp_337;
  wire [0:0] exp_334;
  wire [31:0] exp_1;
  wire [31:0] exp_406;
  wire [31:0] exp_613;
  wire [31:0] exp_612;
  wire [31:0] exp_611;
  wire [31:0] exp_610;
  wire [11:0] exp_609;
  wire [11:0] exp_608;
  wire [11:0] exp_607;
  wire [0:0] exp_561;
  wire [5:0] exp_560;
  wire [0:0] exp_606;
  wire [11:0] exp_602;
  wire [11:0] exp_605;
  wire [6:0] exp_603;
  wire [4:0] exp_604;
  wire [31:0] exp_333;
  wire [0:0] exp_336;
  wire [31:0] exp_335;
  wire [0:0] exp_341;
  wire [0:0] exp_319;
  wire [0:0] exp_314;
  wire [0:0] exp_311;
  wire [31:0] exp_310;
  wire [0:0] exp_313;
  wire [31:0] exp_312;
  wire [0:0] exp_318;
  wire [0:0] exp_218;
  wire [0:0] exp_213;
  wire [0:0] exp_210;
  wire [31:0] exp_209;
  wire [0:0] exp_212;
  wire [31:0] exp_211;
  wire [0:0] exp_217;
  wire [0:0] exp_196;
  wire [0:0] exp_191;
  wire [0:0] exp_188;
  wire [31:0] exp_187;
  wire [0:0] exp_190;
  wire [31:0] exp_189;
  wire [0:0] exp_195;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [31:0] exp_146;
  wire [0:0] exp_149;
  wire [31:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [12:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_411;
  wire [0:0] exp_696;
  wire [0:0] exp_695;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_176;
  wire [0:0] exp_183;
  wire [0:0] exp_198;
  wire [0:0] exp_205;
  wire [0:0] exp_222;
  wire [0:0] exp_225;
  wire [0:0] exp_220;
  wire [0:0] exp_283;
  wire [0:0] exp_268;
  wire [0:0] exp_282;
  wire [0:0] exp_279;
  wire [0:0] exp_278;
  wire [0:0] exp_242;
  wire [0:0] exp_266;
  wire [0:0] exp_262;
  wire [0:0] exp_227;
  wire [0:0] exp_240;
  wire [0:0] exp_237;
  wire [0:0] exp_219;
  wire [0:0] exp_206;
  wire [0:0] exp_214;
  wire [0:0] exp_207;
  wire [0:0] exp_239;
  wire [0:0] exp_238;
  wire [0:0] exp_236;
  wire [0:0] exp_230;
  wire [8:0] exp_228;
  wire [8:0] exp_235;
  wire [0:0] exp_234;
  wire [8:0] exp_232;
  wire [0:0] exp_231;
  wire [0:0] exp_233;
  wire [8:0] exp_229;
  wire [0:0] exp_226;
  wire [0:0] exp_265;
  wire [0:0] exp_264;
  wire [0:0] exp_263;
  wire [0:0] exp_251;
  wire [0:0] exp_245;
  wire [8:0] exp_243;
  wire [8:0] exp_250;
  wire [0:0] exp_249;
  wire [8:0] exp_247;
  wire [0:0] exp_246;
  wire [0:0] exp_248;
  wire [8:0] exp_244;
  wire [0:0] exp_261;
  wire [0:0] exp_255;
  wire [2:0] exp_253;
  wire [2:0] exp_260;
  wire [0:0] exp_259;
  wire [2:0] exp_257;
  wire [0:0] exp_256;
  wire [0:0] exp_258;
  wire [0:0] exp_252;
  wire [2:0] exp_254;
  wire [0:0] exp_241;
  wire [0:0] exp_281;
  wire [0:0] exp_280;
  wire [0:0] exp_277;
  wire [0:0] exp_271;
  wire [8:0] exp_269;
  wire [8:0] exp_276;
  wire [0:0] exp_275;
  wire [8:0] exp_273;
  wire [0:0] exp_272;
  wire [0:0] exp_274;
  wire [8:0] exp_270;
  wire [0:0] exp_267;
  wire [0:0] exp_224;
  wire [0:0] exp_223;
  wire [0:0] exp_221;
  wire [0:0] exp_306;
  wire [0:0] exp_322;
  wire [0:0] exp_329;
  wire [7:0] exp_403;
  wire [7:0] exp_405;
  wire [0:0] exp_325;
  wire [6:0] exp_404;
  wire [0:0] exp_402;
  wire [0:0] exp_367;
  wire [0:0] exp_391;
  wire [0:0] exp_387;
  wire [0:0] exp_351;
  wire [0:0] exp_365;
  wire [0:0] exp_362;
  wire [0:0] exp_347;
  wire [0:0] exp_349;
  wire [0:0] exp_345;
  wire [0:0] exp_399;
  wire [0:0] exp_393;
  wire [0:0] exp_398;
  wire [0:0] exp_395;
  wire [0:0] exp_394;
  wire [0:0] exp_376;
  wire [0:0] exp_370;
  wire [8:0] exp_368;
  wire [8:0] exp_375;
  wire [0:0] exp_374;
  wire [8:0] exp_372;
  wire [0:0] exp_371;
  wire [0:0] exp_373;
  wire [8:0] exp_369;
  wire [0:0] exp_386;
  wire [0:0] exp_380;
  wire [2:0] exp_378;
  wire [2:0] exp_385;
  wire [0:0] exp_384;
  wire [2:0] exp_382;
  wire [0:0] exp_381;
  wire [0:0] exp_383;
  wire [0:0] exp_377;
  wire [2:0] exp_379;
  wire [0:0] exp_397;
  wire [0:0] exp_396;
  wire [0:0] exp_344;
  wire [0:0] exp_330;
  wire [0:0] exp_338;
  wire [0:0] exp_343;
  wire [0:0] exp_331;
  wire [0:0] exp_392;
  wire [0:0] exp_348;
  wire [0:0] exp_346;
  wire [0:0] exp_361;
  wire [0:0] exp_364;
  wire [0:0] exp_363;
  wire [0:0] exp_360;
  wire [0:0] exp_354;
  wire [9:0] exp_352;
  wire [9:0] exp_359;
  wire [0:0] exp_358;
  wire [9:0] exp_356;
  wire [0:0] exp_355;
  wire [0:0] exp_357;
  wire [9:0] exp_353;
  wire [0:0] exp_350;
  wire [0:0] exp_390;
  wire [0:0] exp_389;
  wire [0:0] exp_388;
  wire [0:0] exp_366;
  wire [0:0] exp_401;
  wire [0:0] exp_400;
  wire [0:0] exp_1006;
  wire [0:0] exp_1005;
  wire [0:0] exp_420;
  wire [0:0] exp_463;
  wire [31:0] exp_435;
  wire [0:0] exp_434;
  wire [1:0] exp_443;
  wire [4:0] exp_430;
  wire [0:0] exp_433;
  wire [0:0] exp_1012;
  wire [0:0] exp_1011;
  wire [4:0] exp_429;
  wire [31:0] exp_431;
  wire [31:0] exp_1008;
  wire [0:0] exp_1007;
  wire [31:0] exp_644;
  wire [0:0] exp_643;
  wire [31:0] exp_595;
  wire [2:0] exp_538;
  wire [2:0] exp_529;
  wire [0:0] exp_526;
  wire [0:0] exp_460;
  wire [6:0] exp_450;
  wire [6:0] exp_459;
  wire [0:0] exp_462;
  wire [6:0] exp_461;
  wire [0:0] exp_528;
  wire [2:0] exp_516;
  wire [0:0] exp_458;
  wire [4:0] exp_457;
  wire [0:0] exp_515;
  wire [2:0] exp_503;
  wire [0:0] exp_456;
  wire [5:0] exp_455;
  wire [0:0] exp_502;
  wire [2:0] exp_452;
  wire [0:0] exp_501;
  wire [0:0] exp_514;
  wire [0:0] exp_527;
  wire [0:0] exp_533;
  wire [0:0] exp_594;
  wire [31:0] exp_574;
  wire [0:0] exp_540;
  wire [0:0] exp_532;
  wire [0:0] exp_518;
  wire [0:0] exp_505;
  wire [0:0] exp_491;
  wire [0:0] exp_489;
  wire [0:0] exp_490;
  wire [0:0] exp_454;
  wire [4:0] exp_453;
  wire [0:0] exp_504;
  wire [0:0] exp_517;
  wire [0:0] exp_531;
  wire [0:0] exp_530;
  wire [0:0] exp_573;
  wire [31:0] exp_571;
  wire [31:0] exp_536;
  wire [31:0] exp_522;
  wire [0:0] exp_519;
  wire [0:0] exp_521;
  wire [31:0] exp_511;
  wire [0:0] exp_510;
  wire [31:0] exp_497;
  wire [0:0] exp_496;
  wire [31:0] exp_495;
  wire [31:0] exp_493;
  wire [19:0] exp_492;
  wire [3:0] exp_494;
  wire [31:0] exp_509;
  wire [31:0] exp_507;
  wire [19:0] exp_506;
  wire [3:0] exp_508;
  wire [31:0] exp_520;
  wire [31:0] exp_537;
  wire [31:0] exp_525;
  wire [0:0] exp_523;
  wire [0:0] exp_524;
  wire [31:0] exp_513;
  wire [0:0] exp_512;
  wire [31:0] exp_500;
  wire [0:0] exp_499;
  wire [31:0] exp_484;
  wire [0:0] exp_483;
  wire [31:0] exp_478;
  wire [0:0] exp_474;
  wire [4:0] exp_449;
  wire [0:0] exp_473;
  wire [0:0] exp_477;
  wire [31:0] exp_466;
  wire [0:0] exp_446;
  wire [0:0] exp_1022;
  wire [0:0] exp_1021;
  wire [0:0] exp_1020;
  wire [0:0] exp_1019;
  wire [4:0] exp_428;
  wire [0:0] exp_465;
  wire [31:0] exp_442;
  wire [0:0] exp_441;
  wire [1:0] exp_444;
  wire [4:0] exp_437;
  wire [0:0] exp_440;
  wire [0:0] exp_1014;
  wire [0:0] exp_1013;
  wire [4:0] exp_436;
  wire [31:0] exp_438;
  wire [31:0] exp_447;
  wire [31:0] exp_476;
  wire [0:0] exp_475;
  wire [31:0] exp_482;
  wire [31:0] exp_479;
  wire [31:0] exp_481;
  wire [11:0] exp_480;
  wire [31:0] exp_498;
  wire [31:0] exp_426;
  wire [0:0] exp_425;
  wire [31:0] exp_572;
  wire [31:0] exp_576;
  wire [31:0] exp_575;
  wire [5:0] exp_570;
  wire [5:0] exp_569;
  wire [5:0] exp_568;
  wire [4:0] exp_539;
  wire [4:0] exp_488;
  wire [0:0] exp_487;
  wire [4:0] exp_486;
  wire [4:0] exp_451;
  wire [31:0] exp_592;
  wire [1:0] exp_578;
  wire [0:0] exp_577;
  wire [31:0] exp_593;
  wire [1:0] exp_584;
  wire [0:0] exp_583;
  wire [31:0] exp_580;
  wire [31:0] exp_579;
  wire [31:0] exp_582;
  wire [31:0] exp_581;
  wire [31:0] exp_585;
  wire [31:0] exp_589;
  wire [32:0] exp_588;
  wire [32:0] exp_586;
  wire [0:0] exp_567;
  wire [0:0] exp_541;
  wire [0:0] exp_485;
  wire [0:0] exp_566;
  wire [0:0] exp_565;
  wire [0:0] exp_564;
  wire [32:0] exp_587;
  wire [31:0] exp_590;
  wire [31:0] exp_591;
  wire [31:0] exp_642;
  wire [0:0] exp_641;
  wire [31:0] exp_632;
  wire [7:0] exp_631;
  wire [7:0] exp_630;
  wire [7:0] exp_625;
  wire [1:0] exp_616;
  wire [1:0] exp_615;
  wire [1:0] exp_614;
  wire [0:0] exp_624;
  wire [7:0] exp_620;
  wire [31:0] exp_408;
  wire [31:0] exp_340;
  wire [0:0] exp_339;
  wire [31:0] exp_317;
  wire [0:0] exp_316;
  wire [31:0] exp_216;
  wire [0:0] exp_215;
  wire [31:0] exp_194;
  wire [0:0] exp_193;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [10:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_412;
  wire [3:0] exp_693;
  wire [0:0] exp_692;
  wire [3:0] exp_680;
  wire [3:0] exp_676;
  wire [1:0] exp_679;
  wire [1:0] exp_678;
  wire [1:0] exp_677;
  wire [3:0] exp_685;
  wire [3:0] exp_681;
  wire [0:0] exp_684;
  wire [0:0] exp_683;
  wire [0:0] exp_682;
  wire [3:0] exp_686;
  wire [3:0] exp_687;
  wire [3:0] exp_688;
  wire [3:0] exp_689;
  wire [3:0] exp_690;
  wire [3:0] exp_691;
  wire [10:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_407;
  wire [31:0] exp_675;
  wire [0:0] exp_674;
  wire [31:0] exp_662;
  wire [0:0] exp_661;
  wire [31:0] exp_648;
  wire [7:0] exp_647;
  wire [7:0] exp_646;
  wire [7:0] exp_645;
  wire [31:0] exp_535;
  wire [31:0] exp_656;
  wire [3:0] exp_655;
  wire [31:0] exp_658;
  wire [4:0] exp_657;
  wire [31:0] exp_660;
  wire [4:0] exp_659;
  wire [31:0] exp_666;
  wire [0:0] exp_619;
  wire [0:0] exp_618;
  wire [0:0] exp_617;
  wire [0:0] exp_665;
  wire [31:0] exp_652;
  wire [15:0] exp_651;
  wire [15:0] exp_650;
  wire [15:0] exp_649;
  wire [31:0] exp_664;
  wire [4:0] exp_663;
  wire [31:0] exp_668;
  wire [31:0] exp_667;
  wire [31:0] exp_654;
  wire [31:0] exp_653;
  wire [31:0] exp_669;
  wire [31:0] exp_670;
  wire [31:0] exp_671;
  wire [31:0] exp_672;
  wire [31:0] exp_673;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [10:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [10:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [10:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [10:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [10:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [10:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [10:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [10:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [10:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [10:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [10:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [10:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_179;
  wire [0:0] exp_177;
  wire [31:0] exp_139;
  wire [0:0] exp_178;
  wire [31:0] exp_157;
  wire [31:0] exp_164;
  wire [0:0] exp_159;
  wire [31:0] exp_158;
  wire [0:0] exp_163;
  wire [31:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [31:0] exp_167;
  wire [31:0] exp_174;
  wire [0:0] exp_169;
  wire [31:0] exp_168;
  wire [0:0] exp_173;
  wire [31:0] exp_171;
  wire [0:0] exp_170;
  wire [0:0] exp_172;
  wire [0:0] exp_166;
  wire [0:0] exp_165;
  wire [31:0] exp_182;
  wire [31:0] exp_201;
  wire [31:0] exp_204;
  wire [31:0] exp_302;
  wire [31:0] exp_305;
  wire [31:0] exp_320;
  wire [31:0] exp_328;
  wire [7:0] exp_621;
  wire [7:0] exp_622;
  wire [7:0] exp_623;
  wire [31:0] exp_635;
  wire [15:0] exp_634;
  wire [15:0] exp_633;
  wire [15:0] exp_629;
  wire [0:0] exp_628;
  wire [15:0] exp_626;
  wire [15:0] exp_627;
  wire [31:0] exp_636;
  wire [31:0] exp_637;
  wire [31:0] exp_638;
  wire [31:0] exp_639;
  wire [31:0] exp_640;
  wire [31:0] exp_999;
  wire [0:0] exp_998;
  wire [31:0] exp_995;
  wire [0:0] exp_766;
  wire [0:0] exp_765;
  wire [0:0] exp_764;
  wire [0:0] exp_994;
  wire [31:0] exp_990;
  wire [63:0] exp_989;
  wire [0:0] exp_986;
  wire [0:0] exp_969;
  wire [0:0] exp_946;
  wire [0:0] exp_943;
  wire [0:0] exp_941;
  wire [0:0] exp_923;
  wire [0:0] exp_922;
  wire [0:0] exp_921;
  wire [31:0] exp_919;
  wire [0:0] exp_918;
  wire [0:0] exp_917;
  wire [0:0] exp_906;
  wire [0:0] exp_905;
  wire [0:0] exp_769;
  wire [0:0] exp_768;
  wire [0:0] exp_767;
  wire [0:0] exp_772;
  wire [0:0] exp_771;
  wire [1:0] exp_770;
  wire [0:0] exp_942;
  wire [0:0] exp_926;
  wire [0:0] exp_925;
  wire [0:0] exp_924;
  wire [31:0] exp_920;
  wire [0:0] exp_907;
  wire [0:0] exp_928;
  wire [0:0] exp_927;
  wire [0:0] exp_948;
  wire [1:0] exp_947;
  wire [0:0] exp_971;
  wire [1:0] exp_970;
  wire [0:0] exp_988;
  wire [63:0] exp_985;
  wire [63:0] exp_984;
  wire [63:0] exp_980;
  wire [63:0] exp_976;
  wire [63:0] exp_972;
  wire [31:0] exp_965;
  wire [31:0] exp_952;
  wire [31:0] exp_950;
  wire [15:0] exp_949;
  wire [31:0] exp_944;
  wire [31:0] exp_934;
  wire [31:0] exp_933;
  wire [31:0] exp_932;
  wire [0:0] exp_929;
  wire [0:0] exp_931;
  wire [31:0] exp_930;
  wire [15:0] exp_951;
  wire [31:0] exp_945;
  wire [31:0] exp_940;
  wire [31:0] exp_939;
  wire [31:0] exp_938;
  wire [0:0] exp_935;
  wire [0:0] exp_937;
  wire [31:0] exp_936;
  wire [63:0] exp_975;
  wire [63:0] exp_973;
  wire [31:0] exp_966;
  wire [31:0] exp_956;
  wire [31:0] exp_954;
  wire [15:0] exp_953;
  wire [15:0] exp_955;
  wire [4:0] exp_974;
  wire [63:0] exp_979;
  wire [63:0] exp_977;
  wire [31:0] exp_967;
  wire [31:0] exp_960;
  wire [31:0] exp_958;
  wire [15:0] exp_957;
  wire [15:0] exp_959;
  wire [4:0] exp_978;
  wire [63:0] exp_983;
  wire [63:0] exp_981;
  wire [31:0] exp_968;
  wire [31:0] exp_964;
  wire [31:0] exp_962;
  wire [15:0] exp_961;
  wire [15:0] exp_963;
  wire [5:0] exp_982;
  wire [63:0] exp_987;
  wire [31:0] exp_991;
  wire [31:0] exp_997;
  wire [0:0] exp_790;
  wire [0:0] exp_996;
  wire [31:0] exp_900;
  wire [31:0] exp_894;
  wire [0:0] exp_890;
  wire [0:0] exp_889;
  wire [31:0] exp_838;
  wire [31:0] exp_835;
  wire [31:0] exp_834;
  wire [31:0] exp_833;
  wire [0:0] exp_830;
  wire [0:0] exp_821;
  wire [0:0] exp_820;
  wire [0:0] exp_819;
  wire [31:0] exp_815;
  wire [0:0] exp_813;
  wire [0:0] exp_812;
  wire [0:0] exp_792;
  wire [0:0] exp_791;
  wire [0:0] exp_832;
  wire [31:0] exp_831;
  wire [0:0] exp_823;
  wire [0:0] exp_822;
  wire [0:0] exp_888;
  wire [0:0] exp_893;
  wire [31:0] exp_881;
  wire [31:0] exp_880;
  wire [31:0] exp_879;
  wire [0:0] exp_876;
  wire [0:0] exp_840;
  wire [0:0] exp_836;
  wire [0:0] exp_818;
  wire [0:0] exp_817;
  wire [0:0] exp_816;
  wire [31:0] exp_814;
  wire [0:0] exp_878;
  wire [31:0] exp_874;
  wire [31:0] exp_844;
  wire [31:0] exp_871;
  wire [0:0] exp_805;
  wire [1:0] exp_804;
  wire [0:0] exp_870;
  wire [31:0] exp_863;
  wire [0:0] exp_853;
  wire [0:0] exp_852;
  wire [32:0] exp_851;
  wire [32:0] exp_850;
  wire [32:0] exp_849;
  wire [31:0] exp_847;
  wire [31:0] exp_842;
  wire [32:0] exp_868;
  wire [0:0] exp_867;
  wire [32:0] exp_855;
  wire [0:0] exp_854;
  wire [0:0] exp_866;
  wire [0:0] exp_841;
  wire [0:0] exp_848;
  wire [31:0] exp_846;
  wire [31:0] exp_873;
  wire [0:0] exp_872;
  wire [31:0] exp_865;
  wire [0:0] exp_864;
  wire [31:0] exp_837;
  wire [31:0] exp_829;
  wire [31:0] exp_828;
  wire [31:0] exp_827;
  wire [0:0] exp_824;
  wire [0:0] exp_826;
  wire [31:0] exp_825;
  wire [0:0] exp_845;
  wire [0:0] exp_862;
  wire [31:0] exp_857;
  wire [0:0] exp_856;
  wire [31:0] exp_861;
  wire [31:0] exp_859;
  wire [0:0] exp_858;
  wire [0:0] exp_860;
  wire [0:0] exp_869;
  wire [0:0] exp_843;
  wire [0:0] exp_807;
  wire [5:0] exp_806;
  wire [31:0] exp_877;
  wire [31:0] exp_892;
  wire [0:0] exp_891;
  wire [0:0] exp_809;
  wire [5:0] exp_808;
  wire [31:0] exp_901;
  wire [31:0] exp_899;
  wire [0:0] exp_897;
  wire [0:0] exp_896;
  wire [0:0] exp_895;
  wire [0:0] exp_898;
  wire [31:0] exp_887;
  wire [31:0] exp_886;
  wire [31:0] exp_885;
  wire [0:0] exp_882;
  wire [0:0] exp_839;
  wire [0:0] exp_884;
  wire [31:0] exp_875;
  wire [31:0] exp_883;
  wire [31:0] exp_470;
  wire [0:0] exp_469;
  wire [0:0] exp_699;
  wire [0:0] exp_712;
  wire [0:0] exp_713;
  wire [0:0] exp_700;
  wire [0:0] exp_701;
  wire [0:0] exp_706;
  wire [31:0] exp_703;
  wire [31:0] exp_702;
  wire [31:0] exp_705;
  wire [31:0] exp_704;
  wire [0:0] exp_711;
  wire [31:0] exp_708;
  wire [31:0] exp_707;
  wire [31:0] exp_710;
  wire [31:0] exp_709;
  wire [0:0] exp_1026;
  wire [31:0] exp_1025;
  wire [2:0] exp_1024;
  wire [32:0] exp_756;
  wire [0:0] exp_755;
  wire [31:0] exp_746;
  wire [31:0] exp_745;
  wire [0:0] exp_744;
  wire [31:0] exp_731;
  wire [12:0] exp_730;
  wire [12:0] exp_729;
  wire [12:0] exp_728;
  wire [11:0] exp_727;
  wire [7:0] exp_726;
  wire [1:0] exp_725;
  wire [0:0] exp_720;
  wire [0:0] exp_721;
  wire [5:0] exp_722;
  wire [3:0] exp_723;
  wire [0:0] exp_724;
  wire [31:0] exp_743;
  wire [20:0] exp_742;
  wire [20:0] exp_741;
  wire [20:0] exp_740;
  wire [19:0] exp_739;
  wire [9:0] exp_738;
  wire [8:0] exp_737;
  wire [0:0] exp_732;
  wire [7:0] exp_733;
  wire [0:0] exp_734;
  wire [9:0] exp_735;
  wire [0:0] exp_736;
  wire [31:0] exp_543;
  wire [32:0] exp_754;
  wire [32:0] exp_753;
  wire [31:0] exp_751;
  wire [31:0] exp_750;
  wire [11:0] exp_749;
  wire [11:0] exp_748;
  wire [11:0] exp_747;
  wire [32:0] exp_752;
  wire [0:0] exp_423;
  wire [0:0] exp_80;
  wire [10:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_558;
  wire [0:0] exp_323;
  wire [0:0] exp_308;
  wire [0:0] exp_200;
  wire [0:0] exp_184;
  wire [0:0] exp_192;
  wire [0:0] exp_185;
  wire [31:0] exp_181;
  wire [0:0] exp_301;
  wire [0:0] exp_298;
  wire [0:0] exp_300;
  wire [0:0] exp_297;
  wire [0:0] exp_296;
  wire [0:0] exp_294;
  wire [7:0] exp_285;
  wire [31:0] exp_293;
  wire [0:0] exp_291;
  wire [0:0] exp_292;
  wire [7:0] exp_290;
  wire [0:0] exp_286;
  wire [0:0] exp_289;
  wire [7:0] exp_288;
  wire [0:0] exp_287;
  wire [0:0] exp_284;
  wire [0:0] exp_295;
  wire [0:0] exp_299;

  assign exp_324 = exp_307 & exp_323;
  assign exp_307 = exp_315;
  assign exp_315 = exp_5 & exp_314;
  assign exp_5 = exp_410;
  assign exp_410 = exp_757;
  assign exp_757 = exp_694 & exp_422;
  assign exp_694 = exp_559 | exp_561;
  assign exp_559 = exp_544 == exp_558;
  assign exp_544 = exp_542[6:0];

      reg [31:0] exp_542_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_542_reg <= exp_96;
        end
      end
      assign exp_542 = exp_542_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_424;

      reg [31:0] exp_424_reg = 0;
      always@(posedge clk) begin
        if (exp_423) begin
          exp_424_reg <= exp_1027;
        end
      end
      assign exp_424 = exp_424_reg;
    
  reg [32:0] exp_1027_reg;
  always@(*) begin
    case (exp_1023)
      0:exp_1027_reg <= exp_1025;
      1:exp_1027_reg <= exp_756;
      default:exp_1027_reg <= exp_1026;
    endcase
  end
  assign exp_1027 = exp_1027_reg;
  assign exp_1023 = exp_719 & exp_422;
  assign exp_719 = exp_697 | exp_718;
  assign exp_697 = exp_555 | exp_557;
  assign exp_555 = exp_544 == exp_554;
  assign exp_554 = 111;
  assign exp_557 = exp_544 == exp_556;
  assign exp_556 = 103;

  reg [0:0] exp_718_reg;
  always@(*) begin
    case (exp_563)
      0:exp_718_reg <= exp_716;
      1:exp_718_reg <= exp_715;
      default:exp_718_reg <= exp_717;
    endcase
  end
  assign exp_718 = exp_718_reg;
  assign exp_563 = exp_544 == exp_562;
  assign exp_562 = 99;
  assign exp_717 = 0;
  assign exp_716 = 0;

  reg [0:0] exp_715_reg;
  always@(*) begin
    case (exp_545)
      0:exp_715_reg <= exp_698;
      1:exp_715_reg <= exp_699;
      2:exp_715_reg <= exp_712;
      3:exp_715_reg <= exp_713;
      4:exp_715_reg <= exp_700;
      5:exp_715_reg <= exp_701;
      6:exp_715_reg <= exp_706;
      7:exp_715_reg <= exp_711;
      default:exp_715_reg <= exp_714;
    endcase
  end
  assign exp_715 = exp_715_reg;
  assign exp_545 = exp_542[14:12];
  assign exp_714 = 0;
  assign exp_698 = exp_534 == exp_535;

      reg [31:0] exp_534_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_534_reg <= exp_472;
        end
      end
      assign exp_534 = exp_534_reg;
    
  reg [31:0] exp_472_reg;
  always@(*) begin
    case (exp_468)
      0:exp_472_reg <= exp_464;
      1:exp_472_reg <= exp_470;
      default:exp_472_reg <= exp_471;
    endcase
  end
  assign exp_472 = exp_472_reg;
  assign exp_468 = exp_448 == exp_467;
  assign exp_448 = exp_96[19:15];
  assign exp_467 = 0;
  assign exp_471 = 0;

  reg [31:0] exp_464_reg;
  always@(*) begin
    case (exp_445)
      0:exp_464_reg <= exp_435;
      1:exp_464_reg <= exp_447;
      default:exp_464_reg <= exp_463;
    endcase
  end
  assign exp_464 = exp_464_reg;
  assign exp_445 = exp_1018;
  assign exp_1018 = exp_1017 & exp_414;
  assign exp_1017 = exp_1016 & exp_422;
  assign exp_1016 = exp_1015 & exp_1009;
  assign exp_1015 = exp_427 == exp_1010;
  assign exp_427 = exp_96[19:15];
  assign exp_1010 = exp_542[11:7];
  assign exp_1009 = exp_601 | exp_1004;
  assign exp_601 = exp_600 | exp_559;
  assign exp_600 = exp_599 | exp_553;
  assign exp_599 = exp_598 | exp_551;
  assign exp_598 = exp_597 | exp_557;
  assign exp_597 = exp_596 | exp_555;
  assign exp_596 = exp_547 | exp_549;
  assign exp_547 = exp_544 == exp_546;
  assign exp_546 = 19;
  assign exp_549 = exp_544 == exp_548;
  assign exp_548 = 51;
  assign exp_551 = exp_544 == exp_550;
  assign exp_550 = 55;
  assign exp_553 = exp_544 == exp_552;
  assign exp_552 = 23;
  assign exp_1004 = exp_1003 & exp_763;

  reg [0:0] exp_1003_reg;
  always@(*) begin
    case (exp_789)
      0:exp_1003_reg <= exp_1000;
      1:exp_1003_reg <= exp_1001;
      default:exp_1003_reg <= exp_1002;
    endcase
  end
  assign exp_1003 = exp_1003_reg;
  assign exp_789 = exp_763 & exp_788;
  assign exp_763 = exp_761 & exp_762;
  assign exp_761 = exp_759 == exp_760;
  assign exp_759 = exp_542[6:0];
  assign exp_760 = 51;
  assign exp_762 = exp_542[25:25];
  assign exp_788 = exp_758[2:2];
  assign exp_758 = exp_542[14:12];
  assign exp_1002 = 0;
  assign exp_1000 = exp_993 & exp_763;
  assign exp_993 = exp_908 == exp_992;

      reg [2:0] exp_908_reg = 0;
      always@(posedge clk) begin
        if (exp_904) begin
          exp_908_reg <= exp_915;
        end
      end
      assign exp_908 = exp_908_reg;
    
  reg [2:0] exp_915_reg;
  always@(*) begin
    case (exp_910)
      0:exp_915_reg <= exp_912;
      1:exp_915_reg <= exp_913;
      default:exp_915_reg <= exp_914;
    endcase
  end
  assign exp_915 = exp_915_reg;
  assign exp_910 = exp_908 == exp_909;
  assign exp_909 = 4;
  assign exp_914 = 0;
  assign exp_912 = exp_908 + exp_911;
  assign exp_911 = 1;
  assign exp_913 = 0;
  assign exp_904 = exp_763 & exp_903;
  assign exp_903 = ~exp_902;
  assign exp_902 = exp_758[2:2];
  assign exp_992 = 4;
  assign exp_1001 = exp_811 & exp_763;
  assign exp_811 = exp_795 == exp_810;

      reg [5:0] exp_795_reg = 0;
      always@(posedge clk) begin
        if (exp_789) begin
          exp_795_reg <= exp_802;
        end
      end
      assign exp_795 = exp_795_reg;
    
  reg [5:0] exp_802_reg;
  always@(*) begin
    case (exp_797)
      0:exp_802_reg <= exp_799;
      1:exp_802_reg <= exp_800;
      default:exp_802_reg <= exp_801;
    endcase
  end
  assign exp_802 = exp_802_reg;
  assign exp_797 = exp_795 == exp_796;
  assign exp_796 = 37;
  assign exp_801 = 0;
  assign exp_799 = exp_795 + exp_798;
  assign exp_798 = 1;
  assign exp_800 = 0;
  assign exp_810 = 37;

      reg [0:0] exp_422_reg = 0;
      always@(posedge clk) begin
        if (exp_414) begin
          exp_422_reg <= exp_421;
        end
      end
      assign exp_422 = exp_422_reg;
      assign exp_421 = exp_419 & exp_420;

      reg [0:0] exp_419_reg = 0;
      always@(posedge clk) begin
        if (exp_414) begin
          exp_419_reg <= exp_418;
        end
      end
      assign exp_419 = exp_419_reg;
      assign exp_418 = exp_416 & exp_417;
  assign exp_416 = 1;
  assign exp_417 = ~exp_415;
  assign exp_415 = exp_1028;
  assign exp_1028 = exp_422 & exp_719;
  assign exp_414 = ~exp_413;
  assign exp_413 = exp_1032;
  assign exp_1032 = exp_422 & exp_1031;
  assign exp_1031 = exp_1030 | exp_1006;
  assign exp_1030 = exp_410 & exp_1029;
  assign exp_1029 = ~exp_409;
  assign exp_409 = exp_342;

  reg [0:0] exp_342_reg;
  always@(*) begin
    case (exp_337)
      0:exp_342_reg <= exp_319;
      1:exp_342_reg <= exp_329;
      default:exp_342_reg <= exp_341;
    endcase
  end
  assign exp_342 = exp_342_reg;
  assign exp_337 = exp_334 & exp_336;
  assign exp_334 = exp_1 >= exp_333;
  assign exp_1 = exp_406;
  assign exp_406 = exp_613;
  assign exp_613 = exp_612 + exp_611;
  assign exp_612 = 0;
  assign exp_611 = exp_534 + exp_610;
  assign exp_610 = $signed(exp_609);
  assign exp_609 = exp_608 + exp_607;
  assign exp_608 = 0;

  reg [11:0] exp_607_reg;
  always@(*) begin
    case (exp_561)
      0:exp_607_reg <= exp_602;
      1:exp_607_reg <= exp_605;
      default:exp_607_reg <= exp_606;
    endcase
  end
  assign exp_607 = exp_607_reg;
  assign exp_561 = exp_544 == exp_560;
  assign exp_560 = 35;
  assign exp_606 = 0;
  assign exp_602 = exp_542[31:20];
  assign exp_605 = {exp_603, exp_604};  assign exp_603 = exp_542[31:25];
  assign exp_604 = exp_542[11:7];
  assign exp_333 = 2147483668;
  assign exp_336 = exp_1 <= exp_335;
  assign exp_335 = 2147483668;
  assign exp_341 = 0;

  reg [0:0] exp_319_reg;
  always@(*) begin
    case (exp_314)
      0:exp_319_reg <= exp_218;
      1:exp_319_reg <= exp_306;
      default:exp_319_reg <= exp_318;
    endcase
  end
  assign exp_319 = exp_319_reg;
  assign exp_314 = exp_311 & exp_313;
  assign exp_311 = exp_1 >= exp_310;
  assign exp_310 = 2147483664;
  assign exp_313 = exp_1 <= exp_312;
  assign exp_312 = 2147483664;
  assign exp_318 = 0;

  reg [0:0] exp_218_reg;
  always@(*) begin
    case (exp_213)
      0:exp_218_reg <= exp_196;
      1:exp_218_reg <= exp_205;
      default:exp_218_reg <= exp_217;
    endcase
  end
  assign exp_218 = exp_218_reg;
  assign exp_213 = exp_210 & exp_212;
  assign exp_210 = exp_1 >= exp_209;
  assign exp_209 = 2147483660;
  assign exp_212 = exp_1 <= exp_211;
  assign exp_211 = 2147483660;
  assign exp_217 = 0;

  reg [0:0] exp_196_reg;
  always@(*) begin
    case (exp_191)
      0:exp_196_reg <= exp_155;
      1:exp_196_reg <= exp_183;
      default:exp_196_reg <= exp_195;
    endcase
  end
  assign exp_196 = exp_196_reg;
  assign exp_191 = exp_188 & exp_190;
  assign exp_188 = exp_1 >= exp_187;
  assign exp_187 = 2147483656;
  assign exp_190 = exp_1 <= exp_189;
  assign exp_189 = 2147483656;
  assign exp_195 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 2147483648;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 2147483652;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 8188;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_411;
  assign exp_411 = exp_696;
  assign exp_696 = exp_695 + exp_561;
  assign exp_695 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_176;
  assign exp_176 = 1;
  assign exp_183 = exp_198;
  assign exp_198 = stdout_ready_in;
  assign exp_205 = exp_222;

      reg [0:0] exp_222_reg = 1;
      always@(posedge clk) begin
        if (exp_221) begin
          exp_222_reg <= exp_225;
        end
      end
      assign exp_222 = exp_222_reg;
      assign exp_225 = exp_220 | exp_224;
  assign exp_220 = exp_283;
  assign exp_283 = exp_268 & exp_277;

      reg [0:0] exp_268_reg = 0;
      always@(posedge clk) begin
        if (exp_267) begin
          exp_268_reg <= exp_282;
        end
      end
      assign exp_268 = exp_268_reg;
      assign exp_282 = exp_279 | exp_281;
  assign exp_279 = exp_278 & exp_261;
  assign exp_278 = exp_242 & exp_251;

      reg [0:0] exp_242_reg = 0;
      always@(posedge clk) begin
        if (exp_241) begin
          exp_242_reg <= exp_266;
        end
      end
      assign exp_242 = exp_242_reg;
      assign exp_266 = exp_262 | exp_265;
  assign exp_262 = exp_227 & exp_236;

      reg [0:0] exp_227_reg = 0;
      always@(posedge clk) begin
        if (exp_226) begin
          exp_227_reg <= exp_240;
        end
      end
      assign exp_227 = exp_227_reg;
      assign exp_240 = exp_237 | exp_239;
  assign exp_237 = exp_222 & exp_219;
  assign exp_219 = exp_206 & exp_207;
  assign exp_206 = exp_214;
  assign exp_214 = exp_5 & exp_213;
  assign exp_207 = exp_6;
  assign exp_239 = exp_227 & exp_238;
  assign exp_238 = ~exp_236;
  assign exp_236 = exp_230 & exp_227;
  assign exp_230 = exp_228 == exp_229;

      reg [8:0] exp_228_reg = 0;
      always@(posedge clk) begin
        if (exp_227) begin
          exp_228_reg <= exp_235;
        end
      end
      assign exp_228 = exp_228_reg;
    
  reg [8:0] exp_235_reg;
  always@(*) begin
    case (exp_230)
      0:exp_235_reg <= exp_232;
      1:exp_235_reg <= exp_233;
      default:exp_235_reg <= exp_234;
    endcase
  end
  assign exp_235 = exp_235_reg;
  assign exp_234 = 0;
  assign exp_232 = exp_228 + exp_231;
  assign exp_231 = 1;
  assign exp_233 = 0;
  assign exp_229 = 433;
  assign exp_226 = 1;
  assign exp_265 = exp_242 & exp_264;
  assign exp_264 = ~exp_263;
  assign exp_263 = exp_251 & exp_261;
  assign exp_251 = exp_245 & exp_242;
  assign exp_245 = exp_243 == exp_244;

      reg [8:0] exp_243_reg = 0;
      always@(posedge clk) begin
        if (exp_242) begin
          exp_243_reg <= exp_250;
        end
      end
      assign exp_243 = exp_243_reg;
    
  reg [8:0] exp_250_reg;
  always@(*) begin
    case (exp_245)
      0:exp_250_reg <= exp_247;
      1:exp_250_reg <= exp_248;
      default:exp_250_reg <= exp_249;
    endcase
  end
  assign exp_250 = exp_250_reg;
  assign exp_249 = 0;
  assign exp_247 = exp_243 + exp_246;
  assign exp_246 = 1;
  assign exp_248 = 0;
  assign exp_244 = 433;
  assign exp_261 = exp_255 & exp_252;
  assign exp_255 = exp_253 == exp_254;

      reg [2:0] exp_253_reg = 0;
      always@(posedge clk) begin
        if (exp_252) begin
          exp_253_reg <= exp_260;
        end
      end
      assign exp_253 = exp_253_reg;
    
  reg [2:0] exp_260_reg;
  always@(*) begin
    case (exp_255)
      0:exp_260_reg <= exp_257;
      1:exp_260_reg <= exp_258;
      default:exp_260_reg <= exp_259;
    endcase
  end
  assign exp_260 = exp_260_reg;
  assign exp_259 = 0;
  assign exp_257 = exp_253 + exp_256;
  assign exp_256 = 1;
  assign exp_258 = 0;
  assign exp_252 = exp_242 & exp_251;
  assign exp_254 = 7;
  assign exp_241 = 1;
  assign exp_281 = exp_268 & exp_280;
  assign exp_280 = ~exp_277;
  assign exp_277 = exp_271 & exp_268;
  assign exp_271 = exp_269 == exp_270;

      reg [8:0] exp_269_reg = 0;
      always@(posedge clk) begin
        if (exp_268) begin
          exp_269_reg <= exp_276;
        end
      end
      assign exp_269 = exp_269_reg;
    
  reg [8:0] exp_276_reg;
  always@(*) begin
    case (exp_271)
      0:exp_276_reg <= exp_273;
      1:exp_276_reg <= exp_274;
      default:exp_276_reg <= exp_275;
    endcase
  end
  assign exp_276 = exp_276_reg;
  assign exp_275 = 0;
  assign exp_273 = exp_269 + exp_272;
  assign exp_272 = 1;
  assign exp_274 = 0;
  assign exp_270 = 433;
  assign exp_267 = 1;
  assign exp_224 = exp_222 & exp_223;
  assign exp_223 = ~exp_219;
  assign exp_221 = 1;
  assign exp_306 = exp_322;
  assign exp_322 = stdin_valid_in;
  assign exp_329 = exp_403;

      reg [7:0] exp_403_reg = 0;
      always@(posedge clk) begin
        if (exp_402) begin
          exp_403_reg <= exp_405;
        end
      end
      assign exp_403 = exp_403_reg;
      assign exp_405 = {exp_325, exp_404};  assign exp_325 = buttons_rx;
  assign exp_404 = exp_403[7:1];
  assign exp_402 = exp_367 & exp_401;

      reg [0:0] exp_367_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_367_reg <= exp_391;
        end
      end
      assign exp_367 = exp_367_reg;
      assign exp_391 = exp_387 | exp_390;
  assign exp_387 = exp_351 & exp_360;

      reg [0:0] exp_351_reg = 0;
      always@(posedge clk) begin
        if (exp_350) begin
          exp_351_reg <= exp_365;
        end
      end
      assign exp_351 = exp_351_reg;
      assign exp_365 = exp_362 | exp_364;
  assign exp_362 = exp_347 & exp_361;

      reg [0:0] exp_347_reg = 1;
      always@(posedge clk) begin
        if (exp_346) begin
          exp_347_reg <= exp_349;
        end
      end
      assign exp_347 = exp_347_reg;
      assign exp_349 = exp_345 | exp_348;
  assign exp_345 = exp_399;
  assign exp_399 = exp_393 & exp_344;

      reg [0:0] exp_393_reg = 0;
      always@(posedge clk) begin
        if (exp_392) begin
          exp_393_reg <= exp_398;
        end
      end
      assign exp_393 = exp_393_reg;
      assign exp_398 = exp_395 | exp_397;
  assign exp_395 = exp_394 & exp_386;
  assign exp_394 = exp_367 & exp_376;
  assign exp_376 = exp_370 & exp_367;
  assign exp_370 = exp_368 == exp_369;

      reg [8:0] exp_368_reg = 0;
      always@(posedge clk) begin
        if (exp_367) begin
          exp_368_reg <= exp_375;
        end
      end
      assign exp_368 = exp_368_reg;
    
  reg [8:0] exp_375_reg;
  always@(*) begin
    case (exp_370)
      0:exp_375_reg <= exp_372;
      1:exp_375_reg <= exp_373;
      default:exp_375_reg <= exp_374;
    endcase
  end
  assign exp_375 = exp_375_reg;
  assign exp_374 = 0;
  assign exp_372 = exp_368 + exp_371;
  assign exp_371 = 1;
  assign exp_373 = 0;
  assign exp_369 = 433;
  assign exp_386 = exp_380 & exp_377;
  assign exp_380 = exp_378 == exp_379;

      reg [2:0] exp_378_reg = 0;
      always@(posedge clk) begin
        if (exp_377) begin
          exp_378_reg <= exp_385;
        end
      end
      assign exp_378 = exp_378_reg;
    
  reg [2:0] exp_385_reg;
  always@(*) begin
    case (exp_380)
      0:exp_385_reg <= exp_382;
      1:exp_385_reg <= exp_383;
      default:exp_385_reg <= exp_384;
    endcase
  end
  assign exp_385 = exp_385_reg;
  assign exp_384 = 0;
  assign exp_382 = exp_378 + exp_381;
  assign exp_381 = 1;
  assign exp_383 = 0;
  assign exp_377 = exp_367 & exp_376;
  assign exp_379 = 7;
  assign exp_397 = exp_393 & exp_396;
  assign exp_396 = ~exp_344;
  assign exp_344 = exp_330 & exp_343;
  assign exp_330 = exp_338;
  assign exp_338 = exp_5 & exp_337;
  assign exp_343 = ~exp_331;
  assign exp_331 = exp_6;
  assign exp_392 = 1;
  assign exp_348 = exp_347 & exp_325;
  assign exp_346 = 1;
  assign exp_361 = ~exp_325;
  assign exp_364 = exp_351 & exp_363;
  assign exp_363 = ~exp_360;
  assign exp_360 = exp_354 & exp_351;
  assign exp_354 = exp_352 == exp_353;

      reg [9:0] exp_352_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_352_reg <= exp_359;
        end
      end
      assign exp_352 = exp_352_reg;
    
  reg [9:0] exp_359_reg;
  always@(*) begin
    case (exp_354)
      0:exp_359_reg <= exp_356;
      1:exp_359_reg <= exp_357;
      default:exp_359_reg <= exp_358;
    endcase
  end
  assign exp_359 = exp_359_reg;
  assign exp_358 = 0;
  assign exp_356 = exp_352 + exp_355;
  assign exp_355 = 1;
  assign exp_357 = 0;
  assign exp_353 = 650;
  assign exp_350 = 1;
  assign exp_390 = exp_367 & exp_389;
  assign exp_389 = ~exp_388;
  assign exp_388 = exp_376 & exp_386;
  assign exp_366 = 1;
  assign exp_401 = exp_368 == exp_400;
  assign exp_400 = 0;
  assign exp_1006 = exp_763 & exp_1005;
  assign exp_1005 = ~exp_1003;
  assign exp_420 = ~exp_415;
  assign exp_463 = 0;

  //Create RAM
  reg [31:0] exp_435_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_433) begin
      exp_435_ram[exp_429] <= exp_431;
    end
  end
  assign exp_435 = exp_435_ram[exp_430];
  assign exp_434 = exp_443;
  assign exp_443 = 1;
  assign exp_430 = exp_427;
  assign exp_433 = exp_1012;
  assign exp_1012 = exp_1011 & exp_414;
  assign exp_1011 = exp_1009 & exp_422;
  assign exp_429 = exp_1010;
  assign exp_431 = exp_1008;

  reg [31:0] exp_1008_reg;
  always@(*) begin
    case (exp_1004)
      0:exp_1008_reg <= exp_644;
      1:exp_1008_reg <= exp_999;
      default:exp_1008_reg <= exp_1007;
    endcase
  end
  assign exp_1008 = exp_1008_reg;
  assign exp_1007 = 0;

  reg [31:0] exp_644_reg;
  always@(*) begin
    case (exp_559)
      0:exp_644_reg <= exp_595;
      1:exp_644_reg <= exp_642;
      default:exp_644_reg <= exp_643;
    endcase
  end
  assign exp_644 = exp_644_reg;
  assign exp_643 = 0;

  reg [31:0] exp_595_reg;
  always@(*) begin
    case (exp_538)
      0:exp_595_reg <= exp_574;
      1:exp_595_reg <= exp_576;
      2:exp_595_reg <= exp_592;
      3:exp_595_reg <= exp_593;
      4:exp_595_reg <= exp_585;
      5:exp_595_reg <= exp_589;
      6:exp_595_reg <= exp_590;
      7:exp_595_reg <= exp_591;
      default:exp_595_reg <= exp_594;
    endcase
  end
  assign exp_595 = exp_595_reg;

      reg [2:0] exp_538_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_538_reg <= exp_529;
        end
      end
      assign exp_538 = exp_538_reg;
    
  reg [2:0] exp_529_reg;
  always@(*) begin
    case (exp_526)
      0:exp_529_reg <= exp_516;
      1:exp_529_reg <= exp_527;
      default:exp_529_reg <= exp_528;
    endcase
  end
  assign exp_529 = exp_529_reg;
  assign exp_526 = exp_460 | exp_462;
  assign exp_460 = exp_450 == exp_459;
  assign exp_450 = exp_96[6:0];
  assign exp_459 = 111;
  assign exp_462 = exp_450 == exp_461;
  assign exp_461 = 103;
  assign exp_528 = 0;

  reg [2:0] exp_516_reg;
  always@(*) begin
    case (exp_458)
      0:exp_516_reg <= exp_503;
      1:exp_516_reg <= exp_514;
      default:exp_516_reg <= exp_515;
    endcase
  end
  assign exp_516 = exp_516_reg;
  assign exp_458 = exp_450 == exp_457;
  assign exp_457 = 23;
  assign exp_515 = 0;

  reg [2:0] exp_503_reg;
  always@(*) begin
    case (exp_456)
      0:exp_503_reg <= exp_452;
      1:exp_503_reg <= exp_501;
      default:exp_503_reg <= exp_502;
    endcase
  end
  assign exp_503 = exp_503_reg;
  assign exp_456 = exp_450 == exp_455;
  assign exp_455 = 55;
  assign exp_502 = 0;
  assign exp_452 = exp_96[14:12];
  assign exp_501 = 0;
  assign exp_514 = 0;
  assign exp_527 = 0;
  assign exp_533 = exp_414 & exp_419;
  assign exp_594 = 0;

  reg [31:0] exp_574_reg;
  always@(*) begin
    case (exp_540)
      0:exp_574_reg <= exp_571;
      1:exp_574_reg <= exp_572;
      default:exp_574_reg <= exp_573;
    endcase
  end
  assign exp_574 = exp_574_reg;

      reg [0:0] exp_540_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_540_reg <= exp_532;
        end
      end
      assign exp_540 = exp_540_reg;
      assign exp_532 = exp_518 & exp_531;
  assign exp_518 = exp_505 & exp_517;
  assign exp_505 = exp_491 & exp_504;
  assign exp_491 = exp_489 & exp_490;
  assign exp_489 = exp_96[30:30];
  assign exp_490 = ~exp_454;
  assign exp_454 = exp_450 == exp_453;
  assign exp_453 = 19;
  assign exp_504 = ~exp_456;
  assign exp_517 = ~exp_458;
  assign exp_531 = ~exp_530;
  assign exp_530 = exp_460 | exp_462;
  assign exp_573 = 0;
  assign exp_571 = exp_536 + exp_537;

      reg [31:0] exp_536_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_536_reg <= exp_522;
        end
      end
      assign exp_536 = exp_536_reg;
    
  reg [31:0] exp_522_reg;
  always@(*) begin
    case (exp_519)
      0:exp_522_reg <= exp_511;
      1:exp_522_reg <= exp_520;
      default:exp_522_reg <= exp_521;
    endcase
  end
  assign exp_522 = exp_522_reg;
  assign exp_519 = exp_460 | exp_462;
  assign exp_521 = 0;

  reg [31:0] exp_511_reg;
  always@(*) begin
    case (exp_458)
      0:exp_511_reg <= exp_497;
      1:exp_511_reg <= exp_509;
      default:exp_511_reg <= exp_510;
    endcase
  end
  assign exp_511 = exp_511_reg;
  assign exp_510 = 0;

  reg [31:0] exp_497_reg;
  always@(*) begin
    case (exp_456)
      0:exp_497_reg <= exp_472;
      1:exp_497_reg <= exp_495;
      default:exp_497_reg <= exp_496;
    endcase
  end
  assign exp_497 = exp_497_reg;
  assign exp_496 = 0;
  assign exp_495 = exp_493 << exp_494;
  assign exp_493 = exp_492;
  assign exp_492 = exp_96[31:12];
  assign exp_494 = 12;
  assign exp_509 = exp_507 << exp_508;
  assign exp_507 = exp_506;
  assign exp_506 = exp_96[31:12];
  assign exp_508 = 12;
  assign exp_520 = 4;

      reg [31:0] exp_537_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_537_reg <= exp_525;
        end
      end
      assign exp_537 = exp_537_reg;
    
  reg [31:0] exp_525_reg;
  always@(*) begin
    case (exp_523)
      0:exp_525_reg <= exp_513;
      1:exp_525_reg <= exp_426;
      default:exp_525_reg <= exp_524;
    endcase
  end
  assign exp_525 = exp_525_reg;
  assign exp_523 = exp_460 | exp_462;
  assign exp_524 = 0;

  reg [31:0] exp_513_reg;
  always@(*) begin
    case (exp_458)
      0:exp_513_reg <= exp_500;
      1:exp_513_reg <= exp_426;
      default:exp_513_reg <= exp_512;
    endcase
  end
  assign exp_513 = exp_513_reg;
  assign exp_512 = 0;

  reg [31:0] exp_500_reg;
  always@(*) begin
    case (exp_456)
      0:exp_500_reg <= exp_484;
      1:exp_500_reg <= exp_498;
      default:exp_500_reg <= exp_499;
    endcase
  end
  assign exp_500 = exp_500_reg;
  assign exp_499 = 0;

  reg [31:0] exp_484_reg;
  always@(*) begin
    case (exp_454)
      0:exp_484_reg <= exp_478;
      1:exp_484_reg <= exp_482;
      default:exp_484_reg <= exp_483;
    endcase
  end
  assign exp_484 = exp_484_reg;
  assign exp_483 = 0;

  reg [31:0] exp_478_reg;
  always@(*) begin
    case (exp_474)
      0:exp_478_reg <= exp_466;
      1:exp_478_reg <= exp_476;
      default:exp_478_reg <= exp_477;
    endcase
  end
  assign exp_478 = exp_478_reg;
  assign exp_474 = exp_449 == exp_473;
  assign exp_449 = exp_96[24:20];
  assign exp_473 = 0;
  assign exp_477 = 0;

  reg [31:0] exp_466_reg;
  always@(*) begin
    case (exp_446)
      0:exp_466_reg <= exp_442;
      1:exp_466_reg <= exp_447;
      default:exp_466_reg <= exp_465;
    endcase
  end
  assign exp_466 = exp_466_reg;
  assign exp_446 = exp_1022;
  assign exp_1022 = exp_1021 & exp_414;
  assign exp_1021 = exp_1020 & exp_422;
  assign exp_1020 = exp_1019 & exp_1009;
  assign exp_1019 = exp_428 == exp_1010;
  assign exp_428 = exp_96[24:20];
  assign exp_465 = 0;

  //Create RAM
  reg [31:0] exp_442_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_440) begin
      exp_442_ram[exp_436] <= exp_438;
    end
  end
  assign exp_442 = exp_442_ram[exp_437];
  assign exp_441 = exp_444;
  assign exp_444 = 1;
  assign exp_437 = exp_428;
  assign exp_440 = exp_1014;
  assign exp_1014 = exp_1013 & exp_414;
  assign exp_1013 = exp_1009 & exp_422;
  assign exp_436 = exp_1010;
  assign exp_438 = exp_1008;
  assign exp_447 = exp_1008;
  assign exp_476 = $signed(exp_475);
  assign exp_475 = 0;
  assign exp_482 = exp_479 + exp_481;
  assign exp_479 = 0;
  assign exp_481 = $signed(exp_480);
  assign exp_480 = exp_96[31:20];
  assign exp_498 = 0;

      reg [31:0] exp_426_reg = 0;
      always@(posedge clk) begin
        if (exp_425) begin
          exp_426_reg <= exp_424;
        end
      end
      assign exp_426 = exp_426_reg;
      assign exp_425 = exp_416 & exp_414;
  assign exp_572 = exp_536 - exp_537;
  assign exp_576 = exp_536 << exp_575;
  assign exp_575 = $signed(exp_570);
  assign exp_570 = exp_569 + exp_568;
  assign exp_569 = 0;
  assign exp_568 = exp_539;

      reg [4:0] exp_539_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_539_reg <= exp_488;
        end
      end
      assign exp_539 = exp_539_reg;
    
  reg [4:0] exp_488_reg;
  always@(*) begin
    case (exp_454)
      0:exp_488_reg <= exp_486;
      1:exp_488_reg <= exp_451;
      default:exp_488_reg <= exp_487;
    endcase
  end
  assign exp_488 = exp_488_reg;
  assign exp_487 = 0;
  assign exp_486 = exp_484[4:0];
  assign exp_451 = exp_96[24:20];
  assign exp_592 = $signed(exp_578);
  assign exp_578 = exp_577;
  assign exp_577 = $signed(exp_536) < $signed(exp_537);
  assign exp_593 = $signed(exp_584);
  assign exp_584 = exp_583;
  assign exp_583 = exp_580 < exp_582;
  assign exp_580 = exp_579 + exp_536;
  assign exp_579 = 0;
  assign exp_582 = exp_581 + exp_537;
  assign exp_581 = 0;
  assign exp_585 = exp_536 ^ exp_537;
  assign exp_589 = exp_588[31:0];
  assign exp_588 = $signed(exp_586) >>> $signed(exp_587);
  assign exp_586 = {exp_567, exp_536};
  reg [0:0] exp_567_reg;
  always@(*) begin
    case (exp_541)
      0:exp_567_reg <= exp_565;
      1:exp_567_reg <= exp_564;
      default:exp_567_reg <= exp_566;
    endcase
  end
  assign exp_567 = exp_567_reg;

      reg [0:0] exp_541_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_541_reg <= exp_485;
        end
      end
      assign exp_541 = exp_541_reg;
      assign exp_485 = exp_96[30:30];
  assign exp_566 = 0;
  assign exp_565 = 0;
  assign exp_564 = exp_536[31:31];
  assign exp_587 = $signed(exp_570);
  assign exp_590 = exp_536 | exp_537;
  assign exp_591 = exp_536 & exp_537;

  reg [31:0] exp_642_reg;
  always@(*) begin
    case (exp_545)
      0:exp_642_reg <= exp_632;
      1:exp_642_reg <= exp_635;
      2:exp_642_reg <= exp_408;
      3:exp_642_reg <= exp_636;
      4:exp_642_reg <= exp_637;
      5:exp_642_reg <= exp_638;
      6:exp_642_reg <= exp_639;
      7:exp_642_reg <= exp_640;
      default:exp_642_reg <= exp_641;
    endcase
  end
  assign exp_642 = exp_642_reg;
  assign exp_641 = 0;
  assign exp_632 = $signed(exp_631);
  assign exp_631 = exp_630 + exp_625;
  assign exp_630 = 0;

  reg [7:0] exp_625_reg;
  always@(*) begin
    case (exp_616)
      0:exp_625_reg <= exp_620;
      1:exp_625_reg <= exp_621;
      2:exp_625_reg <= exp_622;
      3:exp_625_reg <= exp_623;
      default:exp_625_reg <= exp_624;
    endcase
  end
  assign exp_625 = exp_625_reg;
  assign exp_616 = exp_615 + exp_614;
  assign exp_615 = 0;
  assign exp_614 = exp_613[1:0];
  assign exp_624 = 0;
  assign exp_620 = exp_408[7:0];
  assign exp_408 = exp_340;

  reg [31:0] exp_340_reg;
  always@(*) begin
    case (exp_337)
      0:exp_340_reg <= exp_317;
      1:exp_340_reg <= exp_328;
      default:exp_340_reg <= exp_339;
    endcase
  end
  assign exp_340 = exp_340_reg;
  assign exp_339 = 0;

  reg [31:0] exp_317_reg;
  always@(*) begin
    case (exp_314)
      0:exp_317_reg <= exp_216;
      1:exp_317_reg <= exp_305;
      default:exp_317_reg <= exp_316;
    endcase
  end
  assign exp_317 = exp_317_reg;
  assign exp_316 = 0;

  reg [31:0] exp_216_reg;
  always@(*) begin
    case (exp_213)
      0:exp_216_reg <= exp_194;
      1:exp_216_reg <= exp_204;
      default:exp_216_reg <= exp_215;
    endcase
  end
  assign exp_216 = exp_216_reg;
  assign exp_215 = 0;

  reg [31:0] exp_194_reg;
  always@(*) begin
    case (exp_191)
      0:exp_194_reg <= exp_153;
      1:exp_194_reg <= exp_182;
      default:exp_194_reg <= exp_193;
    endcase
  end
  assign exp_194 = exp_194_reg;
  assign exp_193 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 0;
    exp_54_ram[32] = 252;
    exp_54_ram[33] = 10;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 253;
    exp_54_ram[36] = 2;
    exp_54_ram[37] = 3;
    exp_54_ram[38] = 252;
    exp_54_ram[39] = 252;
    exp_54_ram[40] = 253;
    exp_54_ram[41] = 254;
    exp_54_ram[42] = 253;
    exp_54_ram[43] = 254;
    exp_54_ram[44] = 0;
    exp_54_ram[45] = 253;
    exp_54_ram[46] = 0;
    exp_54_ram[47] = 2;
    exp_54_ram[48] = 3;
    exp_54_ram[49] = 0;
    exp_54_ram[50] = 254;
    exp_54_ram[51] = 0;
    exp_54_ram[52] = 2;
    exp_54_ram[53] = 128;
    exp_54_ram[54] = 254;
    exp_54_ram[55] = 128;
    exp_54_ram[56] = 0;
    exp_54_ram[57] = 254;
    exp_54_ram[58] = 254;
    exp_54_ram[59] = 0;
    exp_54_ram[60] = 0;
    exp_54_ram[61] = 254;
    exp_54_ram[62] = 0;
    exp_54_ram[63] = 0;
    exp_54_ram[64] = 0;
    exp_54_ram[65] = 0;
    exp_54_ram[66] = 0;
    exp_54_ram[67] = 0;
    exp_54_ram[68] = 0;
    exp_54_ram[69] = 0;
    exp_54_ram[70] = 0;
    exp_54_ram[71] = 0;
    exp_54_ram[72] = 1;
    exp_54_ram[73] = 2;
    exp_54_ram[74] = 0;
    exp_54_ram[75] = 252;
    exp_54_ram[76] = 2;
    exp_54_ram[77] = 2;
    exp_54_ram[78] = 3;
    exp_54_ram[79] = 3;
    exp_54_ram[80] = 3;
    exp_54_ram[81] = 3;
    exp_54_ram[82] = 3;
    exp_54_ram[83] = 3;
    exp_54_ram[84] = 1;
    exp_54_ram[85] = 1;
    exp_54_ram[86] = 4;
    exp_54_ram[87] = 246;
    exp_54_ram[88] = 252;
    exp_54_ram[89] = 252;
    exp_54_ram[90] = 0;
    exp_54_ram[91] = 245;
    exp_54_ram[92] = 0;
    exp_54_ram[93] = 0;
    exp_54_ram[94] = 252;
    exp_54_ram[95] = 252;
    exp_54_ram[96] = 64;
    exp_54_ram[97] = 0;
    exp_54_ram[98] = 1;
    exp_54_ram[99] = 64;
    exp_54_ram[100] = 65;
    exp_54_ram[101] = 0;
    exp_54_ram[102] = 42;
    exp_54_ram[103] = 0;
    exp_54_ram[104] = 0;
    exp_54_ram[105] = 0;
    exp_54_ram[106] = 0;
    exp_54_ram[107] = 252;
    exp_54_ram[108] = 0;
    exp_54_ram[109] = 0;
    exp_54_ram[110] = 0;
    exp_54_ram[111] = 0;
    exp_54_ram[112] = 250;
    exp_54_ram[113] = 42;
    exp_54_ram[114] = 0;
    exp_54_ram[115] = 0;
    exp_54_ram[116] = 252;
    exp_54_ram[117] = 252;
    exp_54_ram[118] = 1;
    exp_54_ram[119] = 0;
    exp_54_ram[120] = 0;
    exp_54_ram[121] = 1;
    exp_54_ram[122] = 0;
    exp_54_ram[123] = 0;
    exp_54_ram[124] = 252;
    exp_54_ram[125] = 252;
    exp_54_ram[126] = 43;
    exp_54_ram[127] = 0;
    exp_54_ram[128] = 0;
    exp_54_ram[129] = 232;
    exp_54_ram[130] = 0;
    exp_54_ram[131] = 235;
    exp_54_ram[132] = 0;
    exp_54_ram[133] = 0;
    exp_54_ram[134] = 252;
    exp_54_ram[135] = 252;
    exp_54_ram[136] = 64;
    exp_54_ram[137] = 0;
    exp_54_ram[138] = 1;
    exp_54_ram[139] = 64;
    exp_54_ram[140] = 65;
    exp_54_ram[141] = 0;
    exp_54_ram[142] = 42;
    exp_54_ram[143] = 0;
    exp_54_ram[144] = 0;
    exp_54_ram[145] = 0;
    exp_54_ram[146] = 0;
    exp_54_ram[147] = 252;
    exp_54_ram[148] = 0;
    exp_54_ram[149] = 0;
    exp_54_ram[150] = 0;
    exp_54_ram[151] = 0;
    exp_54_ram[152] = 250;
    exp_54_ram[153] = 42;
    exp_54_ram[154] = 0;
    exp_54_ram[155] = 0;
    exp_54_ram[156] = 252;
    exp_54_ram[157] = 252;
    exp_54_ram[158] = 1;
    exp_54_ram[159] = 0;
    exp_54_ram[160] = 0;
    exp_54_ram[161] = 1;
    exp_54_ram[162] = 0;
    exp_54_ram[163] = 0;
    exp_54_ram[164] = 252;
    exp_54_ram[165] = 252;
    exp_54_ram[166] = 43;
    exp_54_ram[167] = 0;
    exp_54_ram[168] = 0;
    exp_54_ram[169] = 222;
    exp_54_ram[170] = 236;
    exp_54_ram[171] = 2;
    exp_54_ram[172] = 128;
    exp_54_ram[173] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_412;
  assign exp_412 = exp_693;

  reg [3:0] exp_693_reg;
  always@(*) begin
    case (exp_545)
      0:exp_693_reg <= exp_680;
      1:exp_693_reg <= exp_685;
      2:exp_693_reg <= exp_686;
      3:exp_693_reg <= exp_687;
      4:exp_693_reg <= exp_688;
      5:exp_693_reg <= exp_689;
      6:exp_693_reg <= exp_690;
      7:exp_693_reg <= exp_691;
      default:exp_693_reg <= exp_692;
    endcase
  end
  assign exp_693 = exp_693_reg;
  assign exp_692 = 0;
  assign exp_680 = exp_676 << exp_679;
  assign exp_676 = 1;
  assign exp_679 = exp_678 + exp_677;
  assign exp_678 = 0;
  assign exp_677 = exp_613[1:0];
  assign exp_685 = exp_681 << exp_684;
  assign exp_681 = 3;
  assign exp_684 = exp_683 + exp_682;
  assign exp_683 = 0;
  assign exp_682 = exp_613[1:1];
  assign exp_686 = 15;
  assign exp_687 = 0;
  assign exp_688 = 0;
  assign exp_689 = 0;
  assign exp_690 = 0;
  assign exp_691 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_407;
  assign exp_407 = exp_675;

  reg [31:0] exp_675_reg;
  always@(*) begin
    case (exp_545)
      0:exp_675_reg <= exp_662;
      1:exp_675_reg <= exp_666;
      2:exp_675_reg <= exp_668;
      3:exp_675_reg <= exp_669;
      4:exp_675_reg <= exp_670;
      5:exp_675_reg <= exp_671;
      6:exp_675_reg <= exp_672;
      7:exp_675_reg <= exp_673;
      default:exp_675_reg <= exp_674;
    endcase
  end
  assign exp_675 = exp_675_reg;
  assign exp_674 = 0;

  reg [31:0] exp_662_reg;
  always@(*) begin
    case (exp_616)
      0:exp_662_reg <= exp_648;
      1:exp_662_reg <= exp_656;
      2:exp_662_reg <= exp_658;
      3:exp_662_reg <= exp_660;
      default:exp_662_reg <= exp_661;
    endcase
  end
  assign exp_662 = exp_662_reg;
  assign exp_661 = 0;
  assign exp_648 = exp_647;
  assign exp_647 = exp_646 + exp_645;
  assign exp_646 = 0;
  assign exp_645 = exp_535[7:0];

      reg [31:0] exp_535_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_535_reg <= exp_478;
        end
      end
      assign exp_535 = exp_535_reg;
      assign exp_656 = exp_648 << exp_655;
  assign exp_655 = 8;
  assign exp_658 = exp_648 << exp_657;
  assign exp_657 = 16;
  assign exp_660 = exp_648 << exp_659;
  assign exp_659 = 24;

  reg [31:0] exp_666_reg;
  always@(*) begin
    case (exp_619)
      0:exp_666_reg <= exp_652;
      1:exp_666_reg <= exp_664;
      default:exp_666_reg <= exp_665;
    endcase
  end
  assign exp_666 = exp_666_reg;
  assign exp_619 = exp_618 + exp_617;
  assign exp_618 = 0;
  assign exp_617 = exp_613[1:1];
  assign exp_665 = 0;
  assign exp_652 = exp_651;
  assign exp_651 = exp_650 + exp_649;
  assign exp_650 = 0;
  assign exp_649 = exp_535[15:0];
  assign exp_664 = exp_652 << exp_663;
  assign exp_663 = 16;
  assign exp_668 = exp_667 + exp_654;
  assign exp_667 = 0;
  assign exp_654 = exp_653 + exp_535;
  assign exp_653 = 0;
  assign exp_669 = 0;
  assign exp_670 = 0;
  assign exp_671 = 0;
  assign exp_672 = 0;
  assign exp_673 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 0;
    exp_47_ram[32] = 1;
    exp_47_ram[33] = 128;
    exp_47_ram[34] = 0;
    exp_47_ram[35] = 1;
    exp_47_ram[36] = 129;
    exp_47_ram[37] = 1;
    exp_47_ram[38] = 164;
    exp_47_ram[39] = 180;
    exp_47_ram[40] = 132;
    exp_47_ram[41] = 244;
    exp_47_ram[42] = 196;
    exp_47_ram[43] = 196;
    exp_47_ram[44] = 231;
    exp_47_ram[45] = 196;
    exp_47_ram[46] = 7;
    exp_47_ram[47] = 193;
    exp_47_ram[48] = 1;
    exp_47_ram[49] = 0;
    exp_47_ram[50] = 1;
    exp_47_ram[51] = 129;
    exp_47_ram[52] = 1;
    exp_47_ram[53] = 0;
    exp_47_ram[54] = 212;
    exp_47_ram[55] = 0;
    exp_47_ram[56] = 70;
    exp_47_ram[57] = 212;
    exp_47_ram[58] = 196;
    exp_47_ram[59] = 6;
    exp_47_ram[60] = 70;
    exp_47_ram[61] = 132;
    exp_47_ram[62] = 72;
    exp_47_ram[63] = 8;
    exp_47_ram[64] = 8;
    exp_47_ram[65] = 0;
    exp_47_ram[66] = 230;
    exp_47_ram[67] = 246;
    exp_47_ram[68] = 5;
    exp_47_ram[69] = 5;
    exp_47_ram[70] = 7;
    exp_47_ram[71] = 7;
    exp_47_ram[72] = 193;
    exp_47_ram[73] = 1;
    exp_47_ram[74] = 0;
    exp_47_ram[75] = 1;
    exp_47_ram[76] = 17;
    exp_47_ram[77] = 129;
    exp_47_ram[78] = 33;
    exp_47_ram[79] = 49;
    exp_47_ram[80] = 65;
    exp_47_ram[81] = 81;
    exp_47_ram[82] = 97;
    exp_47_ram[83] = 113;
    exp_47_ram[84] = 129;
    exp_47_ram[85] = 145;
    exp_47_ram[86] = 1;
    exp_47_ram[87] = 223;
    exp_47_ram[88] = 164;
    exp_47_ram[89] = 180;
    exp_47_ram[90] = 0;
    exp_47_ram[91] = 223;
    exp_47_ram[92] = 5;
    exp_47_ram[93] = 5;
    exp_47_ram[94] = 132;
    exp_47_ram[95] = 196;
    exp_47_ram[96] = 166;
    exp_47_ram[97] = 7;
    exp_47_ram[98] = 6;
    exp_47_ram[99] = 182;
    exp_47_ram[100] = 7;
    exp_47_ram[101] = 6;
    exp_47_ram[102] = 192;
    exp_47_ram[103] = 6;
    exp_47_ram[104] = 0;
    exp_47_ram[105] = 7;
    exp_47_ram[106] = 11;
    exp_47_ram[107] = 198;
    exp_47_ram[108] = 7;
    exp_47_ram[109] = 11;
    exp_47_ram[110] = 214;
    exp_47_ram[111] = 11;
    exp_47_ram[112] = 231;
    exp_47_ram[113] = 192;
    exp_47_ram[114] = 7;
    exp_47_ram[115] = 0;
    exp_47_ram[116] = 132;
    exp_47_ram[117] = 196;
    exp_47_ram[118] = 70;
    exp_47_ram[119] = 7;
    exp_47_ram[120] = 197;
    exp_47_ram[121] = 86;
    exp_47_ram[122] = 245;
    exp_47_ram[123] = 6;
    exp_47_ram[124] = 228;
    exp_47_ram[125] = 244;
    exp_47_ram[126] = 0;
    exp_47_ram[127] = 7;
    exp_47_ram[128] = 16;
    exp_47_ram[129] = 159;
    exp_47_ram[130] = 0;
    exp_47_ram[131] = 223;
    exp_47_ram[132] = 5;
    exp_47_ram[133] = 5;
    exp_47_ram[134] = 132;
    exp_47_ram[135] = 196;
    exp_47_ram[136] = 166;
    exp_47_ram[137] = 7;
    exp_47_ram[138] = 6;
    exp_47_ram[139] = 182;
    exp_47_ram[140] = 7;
    exp_47_ram[141] = 6;
    exp_47_ram[142] = 192;
    exp_47_ram[143] = 6;
    exp_47_ram[144] = 0;
    exp_47_ram[145] = 7;
    exp_47_ram[146] = 12;
    exp_47_ram[147] = 198;
    exp_47_ram[148] = 7;
    exp_47_ram[149] = 12;
    exp_47_ram[150] = 214;
    exp_47_ram[151] = 12;
    exp_47_ram[152] = 231;
    exp_47_ram[153] = 192;
    exp_47_ram[154] = 7;
    exp_47_ram[155] = 0;
    exp_47_ram[156] = 132;
    exp_47_ram[157] = 196;
    exp_47_ram[158] = 38;
    exp_47_ram[159] = 7;
    exp_47_ram[160] = 197;
    exp_47_ram[161] = 54;
    exp_47_ram[162] = 245;
    exp_47_ram[163] = 6;
    exp_47_ram[164] = 228;
    exp_47_ram[165] = 244;
    exp_47_ram[166] = 0;
    exp_47_ram[167] = 7;
    exp_47_ram[168] = 0;
    exp_47_ram[169] = 159;
    exp_47_ram[170] = 31;
    exp_47_ram[171] = 250;
    exp_47_ram[172] = 0;
    exp_47_ram[173] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 33;
    exp_40_ram[32] = 1;
    exp_40_ram[33] = 0;
    exp_40_ram[34] = 0;
    exp_40_ram[35] = 1;
    exp_40_ram[36] = 38;
    exp_40_ram[37] = 4;
    exp_40_ram[38] = 46;
    exp_40_ram[39] = 44;
    exp_40_ram[40] = 39;
    exp_40_ram[41] = 38;
    exp_40_ram[42] = 39;
    exp_40_ram[43] = 39;
    exp_40_ram[44] = 160;
    exp_40_ram[45] = 39;
    exp_40_ram[46] = 133;
    exp_40_ram[47] = 36;
    exp_40_ram[48] = 1;
    exp_40_ram[49] = 128;
    exp_40_ram[50] = 1;
    exp_40_ram[51] = 46;
    exp_40_ram[52] = 4;
    exp_40_ram[53] = 6;
    exp_40_ram[54] = 38;
    exp_40_ram[55] = 6;
    exp_40_ram[56] = 134;
    exp_40_ram[57] = 36;
    exp_40_ram[58] = 38;
    exp_40_ram[59] = 166;
    exp_40_ram[60] = 166;
    exp_40_ram[61] = 40;
    exp_40_ram[62] = 40;
    exp_40_ram[63] = 40;
    exp_40_ram[64] = 23;
    exp_40_ram[65] = 7;
    exp_40_ram[66] = 101;
    exp_40_ram[67] = 229;
    exp_40_ram[68] = 7;
    exp_40_ram[69] = 135;
    exp_40_ram[70] = 5;
    exp_40_ram[71] = 133;
    exp_40_ram[72] = 36;
    exp_40_ram[73] = 1;
    exp_40_ram[74] = 128;
    exp_40_ram[75] = 1;
    exp_40_ram[76] = 46;
    exp_40_ram[77] = 44;
    exp_40_ram[78] = 42;
    exp_40_ram[79] = 40;
    exp_40_ram[80] = 38;
    exp_40_ram[81] = 36;
    exp_40_ram[82] = 34;
    exp_40_ram[83] = 32;
    exp_40_ram[84] = 46;
    exp_40_ram[85] = 44;
    exp_40_ram[86] = 4;
    exp_40_ram[87] = 240;
    exp_40_ram[88] = 36;
    exp_40_ram[89] = 38;
    exp_40_ram[90] = 0;
    exp_40_ram[91] = 240;
    exp_40_ram[92] = 6;
    exp_40_ram[93] = 134;
    exp_40_ram[94] = 37;
    exp_40_ram[95] = 37;
    exp_40_ram[96] = 7;
    exp_40_ram[97] = 8;
    exp_40_ram[98] = 56;
    exp_40_ram[99] = 135;
    exp_40_ram[100] = 134;
    exp_40_ram[101] = 135;
    exp_40_ram[102] = 38;
    exp_40_ram[103] = 139;
    exp_40_ram[104] = 11;
    exp_40_ram[105] = 134;
    exp_40_ram[106] = 134;
    exp_40_ram[107] = 224;
    exp_40_ram[108] = 134;
    exp_40_ram[109] = 134;
    exp_40_ram[110] = 22;
    exp_40_ram[111] = 7;
    exp_40_ram[112] = 230;
    exp_40_ram[113] = 39;
    exp_40_ram[114] = 138;
    exp_40_ram[115] = 10;
    exp_40_ram[116] = 38;
    exp_40_ram[117] = 38;
    exp_40_ram[118] = 7;
    exp_40_ram[119] = 5;
    exp_40_ram[120] = 181;
    exp_40_ram[121] = 135;
    exp_40_ram[122] = 134;
    exp_40_ram[123] = 135;
    exp_40_ram[124] = 36;
    exp_40_ram[125] = 38;
    exp_40_ram[126] = 39;
    exp_40_ram[127] = 133;
    exp_40_ram[128] = 5;
    exp_40_ram[129] = 240;
    exp_40_ram[130] = 0;
    exp_40_ram[131] = 240;
    exp_40_ram[132] = 6;
    exp_40_ram[133] = 134;
    exp_40_ram[134] = 37;
    exp_40_ram[135] = 37;
    exp_40_ram[136] = 7;
    exp_40_ram[137] = 8;
    exp_40_ram[138] = 56;
    exp_40_ram[139] = 135;
    exp_40_ram[140] = 134;
    exp_40_ram[141] = 135;
    exp_40_ram[142] = 38;
    exp_40_ram[143] = 140;
    exp_40_ram[144] = 12;
    exp_40_ram[145] = 134;
    exp_40_ram[146] = 134;
    exp_40_ram[147] = 224;
    exp_40_ram[148] = 134;
    exp_40_ram[149] = 134;
    exp_40_ram[150] = 22;
    exp_40_ram[151] = 7;
    exp_40_ram[152] = 230;
    exp_40_ram[153] = 39;
    exp_40_ram[154] = 137;
    exp_40_ram[155] = 9;
    exp_40_ram[156] = 38;
    exp_40_ram[157] = 38;
    exp_40_ram[158] = 7;
    exp_40_ram[159] = 5;
    exp_40_ram[160] = 181;
    exp_40_ram[161] = 135;
    exp_40_ram[162] = 134;
    exp_40_ram[163] = 135;
    exp_40_ram[164] = 36;
    exp_40_ram[165] = 38;
    exp_40_ram[166] = 39;
    exp_40_ram[167] = 133;
    exp_40_ram[168] = 5;
    exp_40_ram[169] = 240;
    exp_40_ram[170] = 240;
    exp_40_ram[171] = 240;
    exp_40_ram[172] = 0;
    exp_40_ram[173] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 55;
    exp_33_ram[32] = 19;
    exp_33_ram[33] = 239;
    exp_33_ram[34] = 111;
    exp_33_ram[35] = 19;
    exp_33_ram[36] = 35;
    exp_33_ram[37] = 19;
    exp_33_ram[38] = 35;
    exp_33_ram[39] = 35;
    exp_33_ram[40] = 131;
    exp_33_ram[41] = 35;
    exp_33_ram[42] = 3;
    exp_33_ram[43] = 131;
    exp_33_ram[44] = 35;
    exp_33_ram[45] = 131;
    exp_33_ram[46] = 19;
    exp_33_ram[47] = 3;
    exp_33_ram[48] = 19;
    exp_33_ram[49] = 103;
    exp_33_ram[50] = 19;
    exp_33_ram[51] = 35;
    exp_33_ram[52] = 19;
    exp_33_ram[53] = 183;
    exp_33_ram[54] = 35;
    exp_33_ram[55] = 183;
    exp_33_ram[56] = 147;
    exp_33_ram[57] = 35;
    exp_33_ram[58] = 131;
    exp_33_ram[59] = 3;
    exp_33_ram[60] = 131;
    exp_33_ram[61] = 3;
    exp_33_ram[62] = 131;
    exp_33_ram[63] = 3;
    exp_33_ram[64] = 147;
    exp_33_ram[65] = 19;
    exp_33_ram[66] = 51;
    exp_33_ram[67] = 179;
    exp_33_ram[68] = 19;
    exp_33_ram[69] = 147;
    exp_33_ram[70] = 19;
    exp_33_ram[71] = 147;
    exp_33_ram[72] = 3;
    exp_33_ram[73] = 19;
    exp_33_ram[74] = 103;
    exp_33_ram[75] = 19;
    exp_33_ram[76] = 35;
    exp_33_ram[77] = 35;
    exp_33_ram[78] = 35;
    exp_33_ram[79] = 35;
    exp_33_ram[80] = 35;
    exp_33_ram[81] = 35;
    exp_33_ram[82] = 35;
    exp_33_ram[83] = 35;
    exp_33_ram[84] = 35;
    exp_33_ram[85] = 35;
    exp_33_ram[86] = 19;
    exp_33_ram[87] = 239;
    exp_33_ram[88] = 35;
    exp_33_ram[89] = 35;
    exp_33_ram[90] = 19;
    exp_33_ram[91] = 239;
    exp_33_ram[92] = 19;
    exp_33_ram[93] = 147;
    exp_33_ram[94] = 3;
    exp_33_ram[95] = 131;
    exp_33_ram[96] = 51;
    exp_33_ram[97] = 19;
    exp_33_ram[98] = 51;
    exp_33_ram[99] = 179;
    exp_33_ram[100] = 179;
    exp_33_ram[101] = 147;
    exp_33_ram[102] = 131;
    exp_33_ram[103] = 19;
    exp_33_ram[104] = 147;
    exp_33_ram[105] = 19;
    exp_33_ram[106] = 147;
    exp_33_ram[107] = 227;
    exp_33_ram[108] = 19;
    exp_33_ram[109] = 147;
    exp_33_ram[110] = 99;
    exp_33_ram[111] = 147;
    exp_33_ram[112] = 227;
    exp_33_ram[113] = 131;
    exp_33_ram[114] = 19;
    exp_33_ram[115] = 147;
    exp_33_ram[116] = 3;
    exp_33_ram[117] = 131;
    exp_33_ram[118] = 51;
    exp_33_ram[119] = 147;
    exp_33_ram[120] = 179;
    exp_33_ram[121] = 179;
    exp_33_ram[122] = 179;
    exp_33_ram[123] = 147;
    exp_33_ram[124] = 35;
    exp_33_ram[125] = 35;
    exp_33_ram[126] = 131;
    exp_33_ram[127] = 147;
    exp_33_ram[128] = 19;
    exp_33_ram[129] = 239;
    exp_33_ram[130] = 19;
    exp_33_ram[131] = 239;
    exp_33_ram[132] = 19;
    exp_33_ram[133] = 147;
    exp_33_ram[134] = 3;
    exp_33_ram[135] = 131;
    exp_33_ram[136] = 51;
    exp_33_ram[137] = 19;
    exp_33_ram[138] = 51;
    exp_33_ram[139] = 179;
    exp_33_ram[140] = 179;
    exp_33_ram[141] = 147;
    exp_33_ram[142] = 131;
    exp_33_ram[143] = 19;
    exp_33_ram[144] = 147;
    exp_33_ram[145] = 19;
    exp_33_ram[146] = 147;
    exp_33_ram[147] = 227;
    exp_33_ram[148] = 19;
    exp_33_ram[149] = 147;
    exp_33_ram[150] = 99;
    exp_33_ram[151] = 147;
    exp_33_ram[152] = 227;
    exp_33_ram[153] = 131;
    exp_33_ram[154] = 19;
    exp_33_ram[155] = 147;
    exp_33_ram[156] = 3;
    exp_33_ram[157] = 131;
    exp_33_ram[158] = 51;
    exp_33_ram[159] = 147;
    exp_33_ram[160] = 179;
    exp_33_ram[161] = 179;
    exp_33_ram[162] = 179;
    exp_33_ram[163] = 147;
    exp_33_ram[164] = 35;
    exp_33_ram[165] = 35;
    exp_33_ram[166] = 131;
    exp_33_ram[167] = 147;
    exp_33_ram[168] = 19;
    exp_33_ram[169] = 239;
    exp_33_ram[170] = 111;
    exp_33_ram[171] = 128;
    exp_33_ram[172] = 12;
    exp_33_ram[173] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_179;

  reg [31:0] exp_179_reg;
  always@(*) begin
    case (exp_177)
      0:exp_179_reg <= exp_157;
      1:exp_179_reg <= exp_167;
      default:exp_179_reg <= exp_178;
    endcase
  end
  assign exp_179 = exp_179_reg;
  assign exp_177 = exp_139[2:2];
  assign exp_139 = exp_1;
  assign exp_178 = 0;

      reg [31:0] exp_157_reg = 0;
      always@(posedge clk) begin
        if (exp_156) begin
          exp_157_reg <= exp_164;
        end
      end
      assign exp_157 = exp_157_reg;
    
  reg [31:0] exp_164_reg;
  always@(*) begin
    case (exp_159)
      0:exp_164_reg <= exp_161;
      1:exp_164_reg <= exp_162;
      default:exp_164_reg <= exp_163;
    endcase
  end
  assign exp_164 = exp_164_reg;
  assign exp_159 = exp_157 == exp_158;
  assign exp_158 = 4294967295;
  assign exp_163 = 0;
  assign exp_161 = exp_157 + exp_160;
  assign exp_160 = 1;
  assign exp_162 = 0;
  assign exp_156 = 1;

      reg [31:0] exp_167_reg = 0;
      always@(posedge clk) begin
        if (exp_166) begin
          exp_167_reg <= exp_174;
        end
      end
      assign exp_167 = exp_167_reg;
    
  reg [31:0] exp_174_reg;
  always@(*) begin
    case (exp_169)
      0:exp_174_reg <= exp_171;
      1:exp_174_reg <= exp_172;
      default:exp_174_reg <= exp_173;
    endcase
  end
  assign exp_174 = exp_174_reg;
  assign exp_169 = exp_167 == exp_168;
  assign exp_168 = 4294967295;
  assign exp_173 = 0;
  assign exp_171 = exp_167 + exp_170;
  assign exp_170 = 1;
  assign exp_172 = 0;
  assign exp_166 = exp_159 & exp_165;
  assign exp_165 = 1;
  assign exp_182 = exp_201;
  assign exp_201 = 0;
  assign exp_204 = exp_302;
  assign exp_302 = 0;
  assign exp_305 = exp_320;
  assign exp_320 = stdin_in;
  assign exp_328 = exp_393;
  assign exp_621 = exp_408[15:8];
  assign exp_622 = exp_408[23:16];
  assign exp_623 = exp_408[31:24];
  assign exp_635 = $signed(exp_634);
  assign exp_634 = exp_633 + exp_629;
  assign exp_633 = 0;

  reg [15:0] exp_629_reg;
  always@(*) begin
    case (exp_619)
      0:exp_629_reg <= exp_626;
      1:exp_629_reg <= exp_627;
      default:exp_629_reg <= exp_628;
    endcase
  end
  assign exp_629 = exp_629_reg;
  assign exp_628 = 0;
  assign exp_626 = exp_408[15:0];
  assign exp_627 = exp_408[31:16];
  assign exp_636 = 0;
  assign exp_637 = exp_625;
  assign exp_638 = exp_629;
  assign exp_639 = 0;
  assign exp_640 = 0;

  reg [31:0] exp_999_reg;
  always@(*) begin
    case (exp_789)
      0:exp_999_reg <= exp_995;
      1:exp_999_reg <= exp_997;
      default:exp_999_reg <= exp_998;
    endcase
  end
  assign exp_999 = exp_999_reg;
  assign exp_998 = 0;

  reg [31:0] exp_995_reg;
  always@(*) begin
    case (exp_766)
      0:exp_995_reg <= exp_990;
      1:exp_995_reg <= exp_991;
      default:exp_995_reg <= exp_994;
    endcase
  end
  assign exp_995 = exp_995_reg;
  assign exp_766 = exp_765 & exp_763;
  assign exp_765 = exp_758 == exp_764;
  assign exp_764 = 0;
  assign exp_994 = 0;
  assign exp_990 = exp_989[63:32];

  reg [63:0] exp_989_reg;
  always@(*) begin
    case (exp_986)
      0:exp_989_reg <= exp_985;
      1:exp_989_reg <= exp_987;
      default:exp_989_reg <= exp_988;
    endcase
  end
  assign exp_989 = exp_989_reg;

      reg [0:0] exp_986_reg = 0;
      always@(posedge clk) begin
        if (exp_971) begin
          exp_986_reg <= exp_969;
        end
      end
      assign exp_986 = exp_986_reg;
    
      reg [0:0] exp_969_reg = 0;
      always@(posedge clk) begin
        if (exp_948) begin
          exp_969_reg <= exp_946;
        end
      end
      assign exp_969 = exp_969_reg;
    
      reg [0:0] exp_946_reg = 0;
      always@(posedge clk) begin
        if (exp_928) begin
          exp_946_reg <= exp_943;
        end
      end
      assign exp_946 = exp_946_reg;
      assign exp_943 = exp_941 ^ exp_942;
  assign exp_941 = exp_923 & exp_906;
  assign exp_923 = exp_922 + exp_921;
  assign exp_922 = 0;
  assign exp_921 = exp_919[31:31];

      reg [31:0] exp_919_reg = 0;
      always@(posedge clk) begin
        if (exp_918) begin
          exp_919_reg <= exp_536;
        end
      end
      assign exp_919 = exp_919_reg;
      assign exp_918 = exp_908 == exp_917;
  assign exp_917 = 0;
  assign exp_906 = exp_905 | exp_772;
  assign exp_905 = exp_766 | exp_769;
  assign exp_769 = exp_768 & exp_763;
  assign exp_768 = exp_758 == exp_767;
  assign exp_767 = 1;
  assign exp_772 = exp_771 & exp_763;
  assign exp_771 = exp_758 == exp_770;
  assign exp_770 = 2;
  assign exp_942 = exp_926 & exp_907;
  assign exp_926 = exp_925 + exp_924;
  assign exp_925 = 0;
  assign exp_924 = exp_920[31:31];

      reg [31:0] exp_920_reg = 0;
      always@(posedge clk) begin
        if (exp_918) begin
          exp_920_reg <= exp_537;
        end
      end
      assign exp_920 = exp_920_reg;
      assign exp_907 = exp_766 | exp_769;
  assign exp_928 = exp_908 == exp_927;
  assign exp_927 = 1;
  assign exp_948 = exp_908 == exp_947;
  assign exp_947 = 2;
  assign exp_971 = exp_908 == exp_970;
  assign exp_970 = 3;
  assign exp_988 = 0;

      reg [63:0] exp_985_reg = 0;
      always@(posedge clk) begin
        if (exp_971) begin
          exp_985_reg <= exp_984;
        end
      end
      assign exp_985 = exp_985_reg;
      assign exp_984 = exp_980 + exp_983;
  assign exp_980 = exp_976 + exp_979;
  assign exp_976 = exp_972 + exp_975;
  assign exp_972 = exp_965;

      reg [31:0] exp_965_reg = 0;
      always@(posedge clk) begin
        if (exp_948) begin
          exp_965_reg <= exp_952;
        end
      end
      assign exp_965 = exp_965_reg;
      assign exp_952 = exp_950 * exp_951;
  assign exp_950 = exp_949;
  assign exp_949 = exp_944[15:0];

      reg [31:0] exp_944_reg = 0;
      always@(posedge clk) begin
        if (exp_928) begin
          exp_944_reg <= exp_934;
        end
      end
      assign exp_944 = exp_944_reg;
      assign exp_934 = exp_933 + exp_932;
  assign exp_933 = 0;

  reg [31:0] exp_932_reg;
  always@(*) begin
    case (exp_929)
      0:exp_932_reg <= exp_919;
      1:exp_932_reg <= exp_930;
      default:exp_932_reg <= exp_931;
    endcase
  end
  assign exp_932 = exp_932_reg;
  assign exp_929 = exp_923 & exp_906;
  assign exp_931 = 0;
  assign exp_930 = -exp_919;
  assign exp_951 = exp_945[15:0];

      reg [31:0] exp_945_reg = 0;
      always@(posedge clk) begin
        if (exp_928) begin
          exp_945_reg <= exp_940;
        end
      end
      assign exp_945 = exp_945_reg;
      assign exp_940 = exp_939 + exp_938;
  assign exp_939 = 0;

  reg [31:0] exp_938_reg;
  always@(*) begin
    case (exp_935)
      0:exp_938_reg <= exp_920;
      1:exp_938_reg <= exp_936;
      default:exp_938_reg <= exp_937;
    endcase
  end
  assign exp_938 = exp_938_reg;
  assign exp_935 = exp_926 & exp_907;
  assign exp_937 = 0;
  assign exp_936 = -exp_920;
  assign exp_975 = exp_973 << exp_974;
  assign exp_973 = exp_966;

      reg [31:0] exp_966_reg = 0;
      always@(posedge clk) begin
        if (exp_948) begin
          exp_966_reg <= exp_956;
        end
      end
      assign exp_966 = exp_966_reg;
      assign exp_956 = exp_954 * exp_955;
  assign exp_954 = exp_953;
  assign exp_953 = exp_944[15:0];
  assign exp_955 = exp_945[31:16];
  assign exp_974 = 16;
  assign exp_979 = exp_977 << exp_978;
  assign exp_977 = exp_967;

      reg [31:0] exp_967_reg = 0;
      always@(posedge clk) begin
        if (exp_948) begin
          exp_967_reg <= exp_960;
        end
      end
      assign exp_967 = exp_967_reg;
      assign exp_960 = exp_958 * exp_959;
  assign exp_958 = exp_957;
  assign exp_957 = exp_944[31:16];
  assign exp_959 = exp_945[15:0];
  assign exp_978 = 16;
  assign exp_983 = exp_981 << exp_982;
  assign exp_981 = exp_968;

      reg [31:0] exp_968_reg = 0;
      always@(posedge clk) begin
        if (exp_948) begin
          exp_968_reg <= exp_964;
        end
      end
      assign exp_968 = exp_968_reg;
      assign exp_964 = exp_962 * exp_963;
  assign exp_962 = exp_961;
  assign exp_961 = exp_944[31:16];
  assign exp_963 = exp_945[31:16];
  assign exp_982 = 32;
  assign exp_987 = -exp_985;
  assign exp_991 = exp_989[31:0];

  reg [31:0] exp_997_reg;
  always@(*) begin
    case (exp_790)
      0:exp_997_reg <= exp_900;
      1:exp_997_reg <= exp_901;
      default:exp_997_reg <= exp_996;
    endcase
  end
  assign exp_997 = exp_997_reg;
  assign exp_790 = exp_758[1:1];
  assign exp_996 = 0;

      reg [31:0] exp_900_reg = 0;
      always@(posedge clk) begin
        if (exp_809) begin
          exp_900_reg <= exp_894;
        end
      end
      assign exp_900 = exp_900_reg;
    
  reg [31:0] exp_894_reg;
  always@(*) begin
    case (exp_890)
      0:exp_894_reg <= exp_881;
      1:exp_894_reg <= exp_892;
      default:exp_894_reg <= exp_893;
    endcase
  end
  assign exp_894 = exp_894_reg;
  assign exp_890 = exp_889 & exp_792;
  assign exp_889 = exp_838 == exp_888;

      reg [31:0] exp_838_reg = 0;
      always@(posedge clk) begin
        if (exp_823) begin
          exp_838_reg <= exp_835;
        end
      end
      assign exp_838 = exp_838_reg;
      assign exp_835 = exp_834 + exp_833;
  assign exp_834 = 0;

  reg [31:0] exp_833_reg;
  always@(*) begin
    case (exp_830)
      0:exp_833_reg <= exp_815;
      1:exp_833_reg <= exp_831;
      default:exp_833_reg <= exp_832;
    endcase
  end
  assign exp_833 = exp_833_reg;
  assign exp_830 = exp_821 & exp_792;
  assign exp_821 = exp_820 + exp_819;
  assign exp_820 = 0;
  assign exp_819 = exp_815[31:31];

      reg [31:0] exp_815_reg = 0;
      always@(posedge clk) begin
        if (exp_813) begin
          exp_815_reg <= exp_537;
        end
      end
      assign exp_815 = exp_815_reg;
      assign exp_813 = exp_795 == exp_812;
  assign exp_812 = 0;
  assign exp_792 = ~exp_791;
  assign exp_791 = exp_758[0:0];
  assign exp_832 = 0;
  assign exp_831 = -exp_815;
  assign exp_823 = exp_795 == exp_822;
  assign exp_822 = 1;
  assign exp_888 = 0;
  assign exp_893 = 0;
  assign exp_881 = exp_880 + exp_879;
  assign exp_880 = 0;

  reg [31:0] exp_879_reg;
  always@(*) begin
    case (exp_876)
      0:exp_879_reg <= exp_874;
      1:exp_879_reg <= exp_877;
      default:exp_879_reg <= exp_878;
    endcase
  end
  assign exp_879 = exp_879_reg;
  assign exp_876 = exp_840 & exp_792;

      reg [0:0] exp_840_reg = 0;
      always@(posedge clk) begin
        if (exp_823) begin
          exp_840_reg <= exp_836;
        end
      end
      assign exp_840 = exp_840_reg;
      assign exp_836 = exp_818 ^ exp_821;
  assign exp_818 = exp_817 + exp_816;
  assign exp_817 = 0;
  assign exp_816 = exp_814[31:31];

      reg [31:0] exp_814_reg = 0;
      always@(posedge clk) begin
        if (exp_813) begin
          exp_814_reg <= exp_536;
        end
      end
      assign exp_814 = exp_814_reg;
      assign exp_878 = 0;

      reg [31:0] exp_874_reg = 0;
      always@(posedge clk) begin
        if (exp_807) begin
          exp_874_reg <= exp_844;
        end
      end
      assign exp_874 = exp_874_reg;
    
      reg [31:0] exp_844_reg = 0;
      always@(posedge clk) begin
        if (exp_843) begin
          exp_844_reg <= exp_871;
        end
      end
      assign exp_844 = exp_844_reg;
    
  reg [31:0] exp_871_reg;
  always@(*) begin
    case (exp_805)
      0:exp_871_reg <= exp_863;
      1:exp_871_reg <= exp_869;
      default:exp_871_reg <= exp_870;
    endcase
  end
  assign exp_871 = exp_871_reg;
  assign exp_805 = exp_795 == exp_804;
  assign exp_804 = 2;
  assign exp_870 = 0;

  reg [31:0] exp_863_reg;
  always@(*) begin
    case (exp_853)
      0:exp_863_reg <= exp_857;
      1:exp_863_reg <= exp_861;
      default:exp_863_reg <= exp_862;
    endcase
  end
  assign exp_863 = exp_863_reg;
  assign exp_853 = ~exp_852;
  assign exp_852 = exp_851[32:32];
  assign exp_851 = exp_850 - exp_838;
  assign exp_850 = exp_849;
  assign exp_849 = {exp_847, exp_848};  assign exp_847 = exp_842[31:0];

      reg [31:0] exp_842_reg = 0;
      always@(posedge clk) begin
        if (exp_841) begin
          exp_842_reg <= exp_868;
        end
      end
      assign exp_842 = exp_842_reg;
    
  reg [32:0] exp_868_reg;
  always@(*) begin
    case (exp_805)
      0:exp_868_reg <= exp_855;
      1:exp_868_reg <= exp_866;
      default:exp_868_reg <= exp_867;
    endcase
  end
  assign exp_868 = exp_868_reg;
  assign exp_867 = 0;

  reg [32:0] exp_855_reg;
  always@(*) begin
    case (exp_853)
      0:exp_855_reg <= exp_849;
      1:exp_855_reg <= exp_851;
      default:exp_855_reg <= exp_854;
    endcase
  end
  assign exp_855 = exp_855_reg;
  assign exp_854 = 0;
  assign exp_866 = 0;
  assign exp_841 = 1;
  assign exp_848 = exp_846[31:31];

      reg [31:0] exp_846_reg = 0;
      always@(posedge clk) begin
        if (exp_845) begin
          exp_846_reg <= exp_873;
        end
      end
      assign exp_846 = exp_846_reg;
    
  reg [31:0] exp_873_reg;
  always@(*) begin
    case (exp_805)
      0:exp_873_reg <= exp_865;
      1:exp_873_reg <= exp_837;
      default:exp_873_reg <= exp_872;
    endcase
  end
  assign exp_873 = exp_873_reg;
  assign exp_872 = 0;
  assign exp_865 = exp_846 << exp_864;
  assign exp_864 = 1;

      reg [31:0] exp_837_reg = 0;
      always@(posedge clk) begin
        if (exp_823) begin
          exp_837_reg <= exp_829;
        end
      end
      assign exp_837 = exp_837_reg;
      assign exp_829 = exp_828 + exp_827;
  assign exp_828 = 0;

  reg [31:0] exp_827_reg;
  always@(*) begin
    case (exp_824)
      0:exp_827_reg <= exp_814;
      1:exp_827_reg <= exp_825;
      default:exp_827_reg <= exp_826;
    endcase
  end
  assign exp_827 = exp_827_reg;
  assign exp_824 = exp_818 & exp_792;
  assign exp_826 = 0;
  assign exp_825 = -exp_814;
  assign exp_845 = 1;
  assign exp_862 = 0;
  assign exp_857 = exp_844 << exp_856;
  assign exp_856 = 1;
  assign exp_861 = exp_859 | exp_860;
  assign exp_859 = exp_844 << exp_858;
  assign exp_858 = 1;
  assign exp_860 = 1;
  assign exp_869 = 0;
  assign exp_843 = 1;
  assign exp_807 = exp_795 == exp_806;
  assign exp_806 = 35;
  assign exp_877 = -exp_874;
  assign exp_892 = $signed(exp_891);
  assign exp_891 = -1;
  assign exp_809 = exp_795 == exp_808;
  assign exp_808 = 36;

      reg [31:0] exp_901_reg = 0;
      always@(posedge clk) begin
        if (exp_809) begin
          exp_901_reg <= exp_899;
        end
      end
      assign exp_901 = exp_901_reg;
    
  reg [31:0] exp_899_reg;
  always@(*) begin
    case (exp_897)
      0:exp_899_reg <= exp_887;
      1:exp_899_reg <= exp_814;
      default:exp_899_reg <= exp_898;
    endcase
  end
  assign exp_899 = exp_899_reg;
  assign exp_897 = exp_896 & exp_792;
  assign exp_896 = exp_838 == exp_895;
  assign exp_895 = 0;
  assign exp_898 = 0;
  assign exp_887 = exp_886 + exp_885;
  assign exp_886 = 0;

  reg [31:0] exp_885_reg;
  always@(*) begin
    case (exp_882)
      0:exp_885_reg <= exp_875;
      1:exp_885_reg <= exp_883;
      default:exp_885_reg <= exp_884;
    endcase
  end
  assign exp_885 = exp_885_reg;
  assign exp_882 = exp_839 & exp_792;

      reg [0:0] exp_839_reg = 0;
      always@(posedge clk) begin
        if (exp_823) begin
          exp_839_reg <= exp_818;
        end
      end
      assign exp_839 = exp_839_reg;
      assign exp_884 = 0;

      reg [31:0] exp_875_reg = 0;
      always@(posedge clk) begin
        if (exp_807) begin
          exp_875_reg <= exp_842;
        end
      end
      assign exp_875 = exp_875_reg;
      assign exp_883 = -exp_875;
  assign exp_470 = $signed(exp_469);
  assign exp_469 = 0;
  assign exp_699 = exp_534 != exp_535;
  assign exp_712 = 0;
  assign exp_713 = 0;
  assign exp_700 = $signed(exp_534) < $signed(exp_535);
  assign exp_701 = $signed(exp_534) >= $signed(exp_535);
  assign exp_706 = exp_703 < exp_705;
  assign exp_703 = exp_702 + exp_534;
  assign exp_702 = 0;
  assign exp_705 = exp_704 + exp_535;
  assign exp_704 = 0;
  assign exp_711 = exp_708 >= exp_710;
  assign exp_708 = exp_707 + exp_534;
  assign exp_707 = 0;
  assign exp_710 = exp_709 + exp_535;
  assign exp_709 = 0;
  assign exp_1026 = 0;
  assign exp_1025 = exp_424 + exp_1024;
  assign exp_1024 = 4;

  reg [32:0] exp_756_reg;
  always@(*) begin
    case (exp_557)
      0:exp_756_reg <= exp_746;
      1:exp_756_reg <= exp_754;
      default:exp_756_reg <= exp_755;
    endcase
  end
  assign exp_756 = exp_756_reg;
  assign exp_755 = 0;
  assign exp_746 = exp_745 + exp_543;

  reg [31:0] exp_745_reg;
  always@(*) begin
    case (exp_555)
      0:exp_745_reg <= exp_731;
      1:exp_745_reg <= exp_743;
      default:exp_745_reg <= exp_744;
    endcase
  end
  assign exp_745 = exp_745_reg;
  assign exp_744 = 0;
  assign exp_731 = $signed(exp_730);
  assign exp_730 = exp_729 + exp_728;
  assign exp_729 = 0;
  assign exp_728 = {exp_727, exp_724};  assign exp_727 = {exp_726, exp_723};  assign exp_726 = {exp_725, exp_722};  assign exp_725 = {exp_720, exp_721};  assign exp_720 = exp_542[31:31];
  assign exp_721 = exp_542[7:7];
  assign exp_722 = exp_542[30:25];
  assign exp_723 = exp_542[11:8];
  assign exp_724 = 0;
  assign exp_743 = $signed(exp_742);
  assign exp_742 = exp_741 + exp_740;
  assign exp_741 = 0;
  assign exp_740 = {exp_739, exp_736};  assign exp_739 = {exp_738, exp_735};  assign exp_738 = {exp_737, exp_734};  assign exp_737 = {exp_732, exp_733};  assign exp_732 = exp_542[31:31];
  assign exp_733 = exp_542[19:12];
  assign exp_734 = exp_542[20:20];
  assign exp_735 = exp_542[30:21];
  assign exp_736 = 0;

      reg [31:0] exp_543_reg = 0;
      always@(posedge clk) begin
        if (exp_533) begin
          exp_543_reg <= exp_426;
        end
      end
      assign exp_543 = exp_543_reg;
      assign exp_754 = exp_753 & exp_752;
  assign exp_753 = $signed(exp_751);
  assign exp_751 = exp_534 + exp_750;
  assign exp_750 = $signed(exp_749);
  assign exp_749 = exp_748 + exp_747;
  assign exp_748 = 0;
  assign exp_747 = exp_542[31:20];
  assign exp_752 = 4294967294;
  assign exp_423 = exp_416 & exp_414;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_425;
  assign exp_558 = 3;
  assign exp_323 = ~exp_308;
  assign exp_308 = exp_6;
  assign exp_200 = exp_184 & exp_185;
  assign exp_184 = exp_192;
  assign exp_192 = exp_5 & exp_191;
  assign exp_185 = exp_6;
  assign exp_181 = exp_2;

  reg [0:0] exp_301_reg;
  always@(*) begin
    case (exp_298)
      0:exp_301_reg <= exp_297;
      1:exp_301_reg <= exp_299;
      default:exp_301_reg <= exp_300;
    endcase
  end
  assign exp_301 = exp_301_reg;
  assign exp_298 = exp_222 | exp_268;
  assign exp_300 = 0;

  reg [0:0] exp_297_reg;
  always@(*) begin
    case (exp_227)
      0:exp_297_reg <= exp_294;
      1:exp_297_reg <= exp_295;
      default:exp_297_reg <= exp_296;
    endcase
  end
  assign exp_297 = exp_297_reg;
  assign exp_296 = 0;
  assign exp_294 = exp_285[0:0];

      reg [7:0] exp_285_reg = 0;
      always@(posedge clk) begin
        if (exp_284) begin
          exp_285_reg <= exp_293;
        end
      end
      assign exp_285 = exp_285_reg;
    
  reg [31:0] exp_293_reg;
  always@(*) begin
    case (exp_291)
      0:exp_293_reg <= exp_290;
      1:exp_293_reg <= exp_204;
      default:exp_293_reg <= exp_292;
    endcase
  end
  assign exp_293 = exp_293_reg;
  assign exp_291 = exp_222 & exp_219;
  assign exp_292 = 0;

  reg [7:0] exp_290_reg;
  always@(*) begin
    case (exp_286)
      0:exp_290_reg <= exp_285;
      1:exp_290_reg <= exp_288;
      default:exp_290_reg <= exp_289;
    endcase
  end
  assign exp_290 = exp_290_reg;
  assign exp_286 = exp_242 & exp_251;
  assign exp_289 = 0;
  assign exp_288 = exp_285 >> exp_287;
  assign exp_287 = 1;
  assign exp_284 = 1;
  assign exp_295 = 0;
  assign exp_299 = 1;
  assign stdin_ready_out = exp_324;
  assign stdout_valid_out = exp_200;
  assign stdout_out = exp_181;
  assign leds_tx = exp_301;

endmodule