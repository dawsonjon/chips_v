
module cpu(clk, data_in, data_ready, data_out, address, byte_enable, data_valid, write_read);
  input [31:0] data_in;
  input [0:0] data_ready;
  input [0:0] clk;
  output [31:0] data_out;
  output [31:0] address;
  output [3:0] byte_enable;
  output [0:0] data_valid;
  output [0:0] write_read;
  wire [31:0] exp_268;
  wire [2:0] exp_140;
  wire [31:0] exp_134;
  wire [31:0] exp_17;
  wire [31:0] exp_15;
  wire [31:0] exp_14;
  wire [31:0] exp_12;
  wire [31:0] exp_362;
  wire [0:0] exp_358;
  wire [0:0] exp_310;
  wire [0:0] exp_288;
  wire [0:0] exp_150;
  wire [6:0] exp_138;
  wire [6:0] exp_149;
  wire [0:0] exp_152;
  wire [6:0] exp_151;
  wire [0:0] exp_309;
  wire [0:0] exp_158;
  wire [6:0] exp_157;
  wire [0:0] exp_308;
  wire [0:0] exp_307;
  wire [0:0] exp_306;
  wire [0:0] exp_305;
  wire [0:0] exp_289;
  wire [31:0] exp_126;
  wire [31:0] exp_64;
  wire [0:0] exp_60;
  wire [4:0] exp_40;
  wire [0:0] exp_59;
  wire [0:0] exp_63;
  wire [31:0] exp_56;
  wire [0:0] exp_37;
  wire [0:0] exp_353;
  wire [4:0] exp_19;
  wire [4:0] exp_352;
  wire [4:0] exp_351;
  wire [4:0] exp_350;
  wire [4:0] exp_345;
  wire [0:0] exp_196;
  wire [0:0] exp_195;
  wire [0:0] exp_194;
  wire [0:0] exp_193;
  wire [0:0] exp_192;
  wire [0:0] exp_191;
  wire [0:0] exp_142;
  wire [4:0] exp_141;
  wire [0:0] exp_144;
  wire [5:0] exp_143;
  wire [0:0] exp_146;
  wire [5:0] exp_145;
  wire [0:0] exp_148;
  wire [4:0] exp_147;
  wire [0:0] exp_154;
  wire [1:0] exp_153;
  wire [0:0] exp_10;
  wire [0:0] exp_9;
  wire [0:0] exp_7;
  wire [0:0] exp_6;
  wire [0:0] exp_4;
  wire [0:0] exp_5;
  wire [0:0] exp_3;
  wire [0:0] exp_363;
  wire [0:0] exp_2;
  wire [0:0] exp_1;
  wire [0:0] exp_366;
  wire [0:0] exp_364;
  wire [0:0] exp_287;
  wire [0:0] exp_156;
  wire [5:0] exp_155;
  wire [0:0] exp_365;
  wire [0:0] exp_8;
  wire [0:0] exp_55;
  wire [31:0] exp_27;
  wire [0:0] exp_26;
  wire [1:0] exp_35;
  wire [4:0] exp_22;
  wire [0:0] exp_25;
  wire [0:0] exp_347;
  wire [0:0] exp_346;
  wire [4:0] exp_21;
  wire [31:0] exp_23;
  wire [31:0] exp_237;
  wire [0:0] exp_236;
  wire [31:0] exp_190;
  wire [2:0] exp_130;
  wire [2:0] exp_121;
  wire [0:0] exp_118;
  wire [0:0] exp_52;
  wire [6:0] exp_42;
  wire [6:0] exp_51;
  wire [0:0] exp_54;
  wire [6:0] exp_53;
  wire [0:0] exp_120;
  wire [2:0] exp_108;
  wire [0:0] exp_50;
  wire [4:0] exp_49;
  wire [0:0] exp_107;
  wire [2:0] exp_95;
  wire [0:0] exp_48;
  wire [5:0] exp_47;
  wire [0:0] exp_94;
  wire [2:0] exp_44;
  wire [0:0] exp_93;
  wire [0:0] exp_106;
  wire [0:0] exp_119;
  wire [0:0] exp_125;
  wire [0:0] exp_189;
  wire [31:0] exp_169;
  wire [0:0] exp_132;
  wire [0:0] exp_124;
  wire [0:0] exp_110;
  wire [0:0] exp_97;
  wire [0:0] exp_83;
  wire [0:0] exp_81;
  wire [0:0] exp_82;
  wire [0:0] exp_46;
  wire [4:0] exp_45;
  wire [0:0] exp_96;
  wire [0:0] exp_109;
  wire [0:0] exp_123;
  wire [0:0] exp_122;
  wire [0:0] exp_168;
  wire [31:0] exp_166;
  wire [31:0] exp_128;
  wire [31:0] exp_114;
  wire [0:0] exp_111;
  wire [0:0] exp_113;
  wire [31:0] exp_103;
  wire [0:0] exp_102;
  wire [31:0] exp_89;
  wire [0:0] exp_88;
  wire [31:0] exp_87;
  wire [31:0] exp_85;
  wire [19:0] exp_84;
  wire [3:0] exp_86;
  wire [31:0] exp_101;
  wire [31:0] exp_99;
  wire [19:0] exp_98;
  wire [3:0] exp_100;
  wire [31:0] exp_112;
  wire [31:0] exp_129;
  wire [31:0] exp_117;
  wire [0:0] exp_115;
  wire [0:0] exp_116;
  wire [31:0] exp_105;
  wire [0:0] exp_104;
  wire [31:0] exp_92;
  wire [0:0] exp_91;
  wire [31:0] exp_76;
  wire [0:0] exp_75;
  wire [31:0] exp_70;
  wire [0:0] exp_66;
  wire [4:0] exp_41;
  wire [0:0] exp_65;
  wire [0:0] exp_69;
  wire [31:0] exp_58;
  wire [0:0] exp_38;
  wire [0:0] exp_357;
  wire [4:0] exp_20;
  wire [4:0] exp_356;
  wire [4:0] exp_355;
  wire [4:0] exp_354;
  wire [0:0] exp_57;
  wire [31:0] exp_34;
  wire [0:0] exp_33;
  wire [1:0] exp_36;
  wire [4:0] exp_29;
  wire [0:0] exp_32;
  wire [0:0] exp_349;
  wire [0:0] exp_348;
  wire [4:0] exp_28;
  wire [31:0] exp_30;
  wire [31:0] exp_39;
  wire [31:0] exp_68;
  wire [0:0] exp_67;
  wire [31:0] exp_74;
  wire [31:0] exp_71;
  wire [31:0] exp_73;
  wire [11:0] exp_72;
  wire [31:0] exp_90;
  wire [31:0] exp_18;
  wire [0:0] exp_16;
  wire [31:0] exp_167;
  wire [31:0] exp_171;
  wire [31:0] exp_170;
  wire [5:0] exp_165;
  wire [5:0] exp_164;
  wire [5:0] exp_163;
  wire [4:0] exp_131;
  wire [4:0] exp_80;
  wire [0:0] exp_79;
  wire [4:0] exp_78;
  wire [4:0] exp_43;
  wire [31:0] exp_187;
  wire [1:0] exp_173;
  wire [0:0] exp_172;
  wire [31:0] exp_188;
  wire [1:0] exp_179;
  wire [0:0] exp_178;
  wire [31:0] exp_175;
  wire [31:0] exp_174;
  wire [31:0] exp_177;
  wire [31:0] exp_176;
  wire [31:0] exp_180;
  wire [31:0] exp_184;
  wire [32:0] exp_183;
  wire [32:0] exp_181;
  wire [0:0] exp_162;
  wire [0:0] exp_133;
  wire [0:0] exp_77;
  wire [0:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_159;
  wire [32:0] exp_182;
  wire [31:0] exp_185;
  wire [31:0] exp_186;
  wire [31:0] exp_235;
  wire [0:0] exp_234;
  wire [31:0] exp_225;
  wire [7:0] exp_224;
  wire [7:0] exp_223;
  wire [7:0] exp_218;
  wire [1:0] exp_209;
  wire [1:0] exp_208;
  wire [1:0] exp_207;
  wire [31:0] exp_206;
  wire [31:0] exp_205;
  wire [11:0] exp_204;
  wire [11:0] exp_203;
  wire [11:0] exp_202;
  wire [0:0] exp_201;
  wire [11:0] exp_197;
  wire [11:0] exp_200;
  wire [6:0] exp_198;
  wire [4:0] exp_199;
  wire [0:0] exp_217;
  wire [7:0] exp_213;
  wire [7:0] exp_214;
  wire [7:0] exp_215;
  wire [7:0] exp_216;
  wire [31:0] exp_228;
  wire [15:0] exp_227;
  wire [15:0] exp_226;
  wire [15:0] exp_222;
  wire [0:0] exp_212;
  wire [0:0] exp_211;
  wire [0:0] exp_210;
  wire [0:0] exp_221;
  wire [15:0] exp_219;
  wire [15:0] exp_220;
  wire [31:0] exp_229;
  wire [31:0] exp_230;
  wire [31:0] exp_231;
  wire [31:0] exp_232;
  wire [31:0] exp_233;
  wire [31:0] exp_62;
  wire [0:0] exp_61;
  wire [31:0] exp_127;
  wire [0:0] exp_290;
  wire [0:0] exp_303;
  wire [0:0] exp_304;
  wire [0:0] exp_291;
  wire [0:0] exp_292;
  wire [0:0] exp_297;
  wire [31:0] exp_294;
  wire [31:0] exp_293;
  wire [31:0] exp_296;
  wire [31:0] exp_295;
  wire [0:0] exp_302;
  wire [31:0] exp_299;
  wire [31:0] exp_298;
  wire [31:0] exp_301;
  wire [31:0] exp_300;
  wire [0:0] exp_361;
  wire [31:0] exp_360;
  wire [2:0] exp_359;
  wire [31:0] exp_344;
  wire [0:0] exp_343;
  wire [31:0] exp_337;
  wire [31:0] exp_336;
  wire [0:0] exp_335;
  wire [31:0] exp_322;
  wire [12:0] exp_321;
  wire [12:0] exp_320;
  wire [12:0] exp_319;
  wire [11:0] exp_318;
  wire [7:0] exp_317;
  wire [1:0] exp_316;
  wire [0:0] exp_311;
  wire [0:0] exp_312;
  wire [5:0] exp_313;
  wire [3:0] exp_314;
  wire [0:0] exp_315;
  wire [31:0] exp_334;
  wire [20:0] exp_333;
  wire [20:0] exp_332;
  wire [20:0] exp_331;
  wire [19:0] exp_330;
  wire [9:0] exp_329;
  wire [8:0] exp_328;
  wire [0:0] exp_323;
  wire [7:0] exp_324;
  wire [0:0] exp_325;
  wire [9:0] exp_326;
  wire [0:0] exp_327;
  wire [31:0] exp_135;
  wire [31:0] exp_342;
  wire [31:0] exp_341;
  wire [11:0] exp_340;
  wire [11:0] exp_339;
  wire [11:0] exp_338;
  wire [0:0] exp_11;
  wire [1:0] exp_13;
  wire [0:0] exp_267;
  wire [31:0] exp_255;
  wire [0:0] exp_254;
  wire [31:0] exp_241;
  wire [7:0] exp_240;
  wire [7:0] exp_239;
  wire [7:0] exp_238;
  wire [31:0] exp_249;
  wire [3:0] exp_248;
  wire [31:0] exp_251;
  wire [4:0] exp_250;
  wire [31:0] exp_253;
  wire [4:0] exp_252;
  wire [31:0] exp_259;
  wire [0:0] exp_258;
  wire [31:0] exp_245;
  wire [15:0] exp_244;
  wire [15:0] exp_243;
  wire [15:0] exp_242;
  wire [31:0] exp_257;
  wire [4:0] exp_256;
  wire [31:0] exp_261;
  wire [31:0] exp_260;
  wire [31:0] exp_247;
  wire [31:0] exp_246;
  wire [31:0] exp_262;
  wire [31:0] exp_263;
  wire [31:0] exp_264;
  wire [31:0] exp_265;
  wire [31:0] exp_266;
  wire [3:0] exp_286;
  wire [0:0] exp_285;
  wire [3:0] exp_273;
  wire [3:0] exp_269;
  wire [1:0] exp_272;
  wire [1:0] exp_271;
  wire [1:0] exp_270;
  wire [3:0] exp_278;
  wire [3:0] exp_274;
  wire [0:0] exp_277;
  wire [0:0] exp_276;
  wire [0:0] exp_275;
  wire [3:0] exp_279;
  wire [3:0] exp_280;
  wire [3:0] exp_281;
  wire [3:0] exp_282;
  wire [3:0] exp_283;
  wire [3:0] exp_284;


  reg [31:0] exp_268_reg;
  always@(*) begin
    case (exp_140)
      0:exp_268_reg <= exp_255;
      1:exp_268_reg <= exp_259;
      2:exp_268_reg <= exp_261;
      3:exp_268_reg <= exp_262;
      4:exp_268_reg <= exp_263;
      5:exp_268_reg <= exp_264;
      6:exp_268_reg <= exp_265;
      7:exp_268_reg <= exp_266;
      default:exp_268_reg <= exp_267;
    endcase
  end
  assign exp_268 = exp_268_reg;
  assign exp_140 = exp_134[14:12];

      reg [31:0] exp_134_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_134_reg <= exp_17;
        end
      end
      assign exp_134 = exp_134_reg;
    
      reg [31:0] exp_17_reg = 0;
      always@(posedge clk) begin
        if (exp_16) begin
          exp_17_reg <= exp_15;
        end
      end
      assign exp_17 = exp_17_reg;
    
  reg [31:0] exp_15_reg;
  always@(*) begin
    case (exp_14)
      0:exp_15_reg <= 1048723;
      1:exp_15_reg <= 1056803;
      2:exp_15_reg <= 1081491;
      3:exp_15_reg <= 1056803;
      4:exp_15_reg <= 1081491;
      5:exp_15_reg <= 1056803;
      default:exp_15_reg <= 0;
    endcase
  end
  assign exp_15 = exp_15_reg;
  assign exp_14 = exp_12 >> exp_13;

      reg [31:0] exp_12_reg = 0;
      always@(posedge clk) begin
        if (exp_11) begin
          exp_12_reg <= exp_362;
        end
      end
      assign exp_12 = exp_12_reg;
    
  reg [31:0] exp_362_reg;
  always@(*) begin
    case (exp_358)
      0:exp_362_reg <= exp_360;
      1:exp_362_reg <= exp_344;
      default:exp_362_reg <= exp_361;
    endcase
  end
  assign exp_362 = exp_362_reg;
  assign exp_358 = exp_310 & exp_10;
  assign exp_310 = exp_288 | exp_309;
  assign exp_288 = exp_150 | exp_152;
  assign exp_150 = exp_138 == exp_149;
  assign exp_138 = exp_134[6:0];
  assign exp_149 = 111;
  assign exp_152 = exp_138 == exp_151;
  assign exp_151 = 103;

  reg [0:0] exp_309_reg;
  always@(*) begin
    case (exp_158)
      0:exp_309_reg <= exp_307;
      1:exp_309_reg <= exp_306;
      default:exp_309_reg <= exp_308;
    endcase
  end
  assign exp_309 = exp_309_reg;
  assign exp_158 = exp_138 == exp_157;
  assign exp_157 = 99;
  assign exp_308 = 0;
  assign exp_307 = 0;

  reg [0:0] exp_306_reg;
  always@(*) begin
    case (exp_140)
      0:exp_306_reg <= exp_289;
      1:exp_306_reg <= exp_290;
      2:exp_306_reg <= exp_303;
      3:exp_306_reg <= exp_304;
      4:exp_306_reg <= exp_291;
      5:exp_306_reg <= exp_292;
      6:exp_306_reg <= exp_297;
      7:exp_306_reg <= exp_302;
      default:exp_306_reg <= exp_305;
    endcase
  end
  assign exp_306 = exp_306_reg;
  assign exp_305 = 0;
  assign exp_289 = exp_126 == exp_127;

      reg [31:0] exp_126_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_126_reg <= exp_64;
        end
      end
      assign exp_126 = exp_126_reg;
    
  reg [31:0] exp_64_reg;
  always@(*) begin
    case (exp_60)
      0:exp_64_reg <= exp_56;
      1:exp_64_reg <= exp_62;
      default:exp_64_reg <= exp_63;
    endcase
  end
  assign exp_64 = exp_64_reg;
  assign exp_60 = exp_40 == exp_59;
  assign exp_40 = exp_17[19:15];
  assign exp_59 = 0;
  assign exp_63 = 0;

  reg [31:0] exp_56_reg;
  always@(*) begin
    case (exp_37)
      0:exp_56_reg <= exp_27;
      1:exp_56_reg <= exp_39;
      default:exp_56_reg <= exp_55;
    endcase
  end
  assign exp_56 = exp_56_reg;
  assign exp_37 = exp_353;
  assign exp_353 = exp_19 == exp_352;
  assign exp_19 = exp_17[19:15];
  assign exp_352 = exp_351 & exp_2;
  assign exp_351 = exp_350 & exp_10;
  assign exp_350 = exp_345 & exp_196;
  assign exp_345 = exp_134[11:7];
  assign exp_196 = exp_195 | exp_154;
  assign exp_195 = exp_194 | exp_148;
  assign exp_194 = exp_193 | exp_146;
  assign exp_193 = exp_192 | exp_152;
  assign exp_192 = exp_191 | exp_150;
  assign exp_191 = exp_142 | exp_144;
  assign exp_142 = exp_138 == exp_141;
  assign exp_141 = 19;
  assign exp_144 = exp_138 == exp_143;
  assign exp_143 = 51;
  assign exp_146 = exp_138 == exp_145;
  assign exp_145 = 55;
  assign exp_148 = exp_138 == exp_147;
  assign exp_147 = 23;
  assign exp_154 = exp_138 == exp_153;
  assign exp_153 = 3;

      reg [0:0] exp_10_reg = 0;
      always@(posedge clk) begin
        if (exp_2) begin
          exp_10_reg <= exp_9;
        end
      end
      assign exp_10 = exp_10_reg;
      assign exp_9 = exp_7 & exp_8;

      reg [0:0] exp_7_reg = 0;
      always@(posedge clk) begin
        if (exp_2) begin
          exp_7_reg <= exp_6;
        end
      end
      assign exp_7 = exp_7_reg;
      assign exp_6 = exp_4 & exp_5;
  assign exp_4 = 1;
  assign exp_5 = ~exp_3;
  assign exp_3 = exp_363;
  assign exp_363 = exp_10 & exp_310;
  assign exp_2 = ~exp_1;
  assign exp_1 = exp_366;
  assign exp_366 = exp_364 & exp_365;
  assign exp_364 = exp_10 & exp_287;
  assign exp_287 = exp_154 | exp_156;
  assign exp_156 = exp_138 == exp_155;
  assign exp_155 = 35;
  assign exp_365 = ~data_ready;
  assign exp_8 = ~exp_3;
  assign exp_55 = 0;

  reg [31:0] exp_27_ram [31:0];
  always@(posedge clk) begin
    if (exp_25) begin
        exp_27_ram[exp_21] <= exp_23;
    end
  end
  assign exp_27 = exp_27_ram[exp_22];
  assign exp_26 = exp_35;
  assign exp_35 = 1;
  assign exp_22 = exp_19;
  assign exp_25 = exp_347;
  assign exp_347 = exp_346 & exp_2;
  assign exp_346 = exp_196 & exp_10;
  assign exp_21 = exp_345;
  assign exp_23 = exp_237;

  reg [31:0] exp_237_reg;
  always@(*) begin
    case (exp_154)
      0:exp_237_reg <= exp_190;
      1:exp_237_reg <= exp_235;
      default:exp_237_reg <= exp_236;
    endcase
  end
  assign exp_237 = exp_237_reg;
  assign exp_236 = 0;

  reg [31:0] exp_190_reg;
  always@(*) begin
    case (exp_130)
      0:exp_190_reg <= exp_169;
      1:exp_190_reg <= exp_171;
      2:exp_190_reg <= exp_187;
      3:exp_190_reg <= exp_188;
      4:exp_190_reg <= exp_180;
      5:exp_190_reg <= exp_184;
      6:exp_190_reg <= exp_185;
      7:exp_190_reg <= exp_186;
      default:exp_190_reg <= exp_189;
    endcase
  end
  assign exp_190 = exp_190_reg;

      reg [2:0] exp_130_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_130_reg <= exp_121;
        end
      end
      assign exp_130 = exp_130_reg;
    
  reg [2:0] exp_121_reg;
  always@(*) begin
    case (exp_118)
      0:exp_121_reg <= exp_108;
      1:exp_121_reg <= exp_119;
      default:exp_121_reg <= exp_120;
    endcase
  end
  assign exp_121 = exp_121_reg;
  assign exp_118 = exp_52 | exp_54;
  assign exp_52 = exp_42 == exp_51;
  assign exp_42 = exp_17[6:0];
  assign exp_51 = 111;
  assign exp_54 = exp_42 == exp_53;
  assign exp_53 = 103;
  assign exp_120 = 0;

  reg [2:0] exp_108_reg;
  always@(*) begin
    case (exp_50)
      0:exp_108_reg <= exp_95;
      1:exp_108_reg <= exp_106;
      default:exp_108_reg <= exp_107;
    endcase
  end
  assign exp_108 = exp_108_reg;
  assign exp_50 = exp_42 == exp_49;
  assign exp_49 = 23;
  assign exp_107 = 0;

  reg [2:0] exp_95_reg;
  always@(*) begin
    case (exp_48)
      0:exp_95_reg <= exp_44;
      1:exp_95_reg <= exp_93;
      default:exp_95_reg <= exp_94;
    endcase
  end
  assign exp_95 = exp_95_reg;
  assign exp_48 = exp_42 == exp_47;
  assign exp_47 = 55;
  assign exp_94 = 0;
  assign exp_44 = exp_17[14:12];
  assign exp_93 = 0;
  assign exp_106 = 0;
  assign exp_119 = 0;
  assign exp_125 = exp_2 & exp_7;
  assign exp_189 = 0;

  reg [31:0] exp_169_reg;
  always@(*) begin
    case (exp_132)
      0:exp_169_reg <= exp_166;
      1:exp_169_reg <= exp_167;
      default:exp_169_reg <= exp_168;
    endcase
  end
  assign exp_169 = exp_169_reg;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_132_reg <= exp_124;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_124 = exp_110 & exp_123;
  assign exp_110 = exp_97 & exp_109;
  assign exp_97 = exp_83 & exp_96;
  assign exp_83 = exp_81 & exp_82;
  assign exp_81 = exp_17[30:30];
  assign exp_82 = ~exp_46;
  assign exp_46 = exp_42 == exp_45;
  assign exp_45 = 19;
  assign exp_96 = ~exp_48;
  assign exp_109 = ~exp_50;
  assign exp_123 = ~exp_122;
  assign exp_122 = exp_52 | exp_54;
  assign exp_168 = 0;
  assign exp_166 = exp_128 + exp_129;

      reg [31:0] exp_128_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_128_reg <= exp_114;
        end
      end
      assign exp_128 = exp_128_reg;
    
  reg [31:0] exp_114_reg;
  always@(*) begin
    case (exp_111)
      0:exp_114_reg <= exp_103;
      1:exp_114_reg <= exp_112;
      default:exp_114_reg <= exp_113;
    endcase
  end
  assign exp_114 = exp_114_reg;
  assign exp_111 = exp_52 | exp_54;
  assign exp_113 = 0;

  reg [31:0] exp_103_reg;
  always@(*) begin
    case (exp_50)
      0:exp_103_reg <= exp_89;
      1:exp_103_reg <= exp_101;
      default:exp_103_reg <= exp_102;
    endcase
  end
  assign exp_103 = exp_103_reg;
  assign exp_102 = 0;

  reg [31:0] exp_89_reg;
  always@(*) begin
    case (exp_48)
      0:exp_89_reg <= exp_64;
      1:exp_89_reg <= exp_87;
      default:exp_89_reg <= exp_88;
    endcase
  end
  assign exp_89 = exp_89_reg;
  assign exp_88 = 0;
  assign exp_87 = exp_85 << exp_86;
  assign exp_85 = exp_84;
  assign exp_84 = exp_17[31:12];
  assign exp_86 = 12;
  assign exp_101 = exp_99 << exp_100;
  assign exp_99 = exp_98;
  assign exp_98 = exp_17[31:12];
  assign exp_100 = 12;
  assign exp_112 = 4;

      reg [31:0] exp_129_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_129_reg <= exp_117;
        end
      end
      assign exp_129 = exp_129_reg;
    
  reg [31:0] exp_117_reg;
  always@(*) begin
    case (exp_115)
      0:exp_117_reg <= exp_105;
      1:exp_117_reg <= exp_18;
      default:exp_117_reg <= exp_116;
    endcase
  end
  assign exp_117 = exp_117_reg;
  assign exp_115 = exp_52 | exp_54;
  assign exp_116 = 0;

  reg [31:0] exp_105_reg;
  always@(*) begin
    case (exp_50)
      0:exp_105_reg <= exp_92;
      1:exp_105_reg <= exp_18;
      default:exp_105_reg <= exp_104;
    endcase
  end
  assign exp_105 = exp_105_reg;
  assign exp_104 = 0;

  reg [31:0] exp_92_reg;
  always@(*) begin
    case (exp_48)
      0:exp_92_reg <= exp_76;
      1:exp_92_reg <= exp_90;
      default:exp_92_reg <= exp_91;
    endcase
  end
  assign exp_92 = exp_92_reg;
  assign exp_91 = 0;

  reg [31:0] exp_76_reg;
  always@(*) begin
    case (exp_46)
      0:exp_76_reg <= exp_70;
      1:exp_76_reg <= exp_74;
      default:exp_76_reg <= exp_75;
    endcase
  end
  assign exp_76 = exp_76_reg;
  assign exp_75 = 0;

  reg [31:0] exp_70_reg;
  always@(*) begin
    case (exp_66)
      0:exp_70_reg <= exp_58;
      1:exp_70_reg <= exp_68;
      default:exp_70_reg <= exp_69;
    endcase
  end
  assign exp_70 = exp_70_reg;
  assign exp_66 = exp_41 == exp_65;
  assign exp_41 = exp_17[24:20];
  assign exp_65 = 0;
  assign exp_69 = 0;

  reg [31:0] exp_58_reg;
  always@(*) begin
    case (exp_38)
      0:exp_58_reg <= exp_34;
      1:exp_58_reg <= exp_39;
      default:exp_58_reg <= exp_57;
    endcase
  end
  assign exp_58 = exp_58_reg;
  assign exp_38 = exp_357;
  assign exp_357 = exp_20 == exp_356;
  assign exp_20 = exp_17[24:20];
  assign exp_356 = exp_355 & exp_2;
  assign exp_355 = exp_354 & exp_10;
  assign exp_354 = exp_345 & exp_196;
  assign exp_57 = 0;

  reg [31:0] exp_34_ram [31:0];
  always@(posedge clk) begin
    if (exp_32) begin
        exp_34_ram[exp_28] <= exp_30;
    end
  end
  assign exp_34 = exp_34_ram[exp_29];
  assign exp_33 = exp_36;
  assign exp_36 = 1;
  assign exp_29 = exp_20;
  assign exp_32 = exp_349;
  assign exp_349 = exp_348 & exp_2;
  assign exp_348 = exp_196 & exp_10;
  assign exp_28 = exp_345;
  assign exp_30 = exp_237;
  assign exp_39 = exp_237;
  assign exp_68 = $signed(exp_67);
  assign exp_67 = 0;
  assign exp_74 = exp_71 + exp_73;
  assign exp_71 = 0;
  assign exp_73 = $signed(exp_72);
  assign exp_72 = exp_17[31:20];
  assign exp_90 = 0;

      reg [31:0] exp_18_reg = 0;
      always@(posedge clk) begin
        if (exp_16) begin
          exp_18_reg <= exp_12;
        end
      end
      assign exp_18 = exp_18_reg;
      assign exp_16 = exp_4 & exp_2;
  assign exp_167 = exp_128 - exp_129;
  assign exp_171 = exp_128 << exp_170;
  assign exp_170 = $signed(exp_165);
  assign exp_165 = exp_164 + exp_163;
  assign exp_164 = 0;
  assign exp_163 = exp_131;

      reg [4:0] exp_131_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_131_reg <= exp_80;
        end
      end
      assign exp_131 = exp_131_reg;
    
  reg [4:0] exp_80_reg;
  always@(*) begin
    case (exp_46)
      0:exp_80_reg <= exp_78;
      1:exp_80_reg <= exp_43;
      default:exp_80_reg <= exp_79;
    endcase
  end
  assign exp_80 = exp_80_reg;
  assign exp_79 = 0;
  assign exp_78 = exp_76[4:0];
  assign exp_43 = exp_17[24:20];
  assign exp_187 = $signed(exp_173);
  assign exp_173 = exp_172;
  assign exp_172 = $signed(exp_128) < $signed(exp_129);
  assign exp_188 = $signed(exp_179);
  assign exp_179 = exp_178;
  assign exp_178 = exp_175 < exp_177;
  assign exp_175 = exp_174 + exp_128;
  assign exp_174 = 0;
  assign exp_177 = exp_176 + exp_129;
  assign exp_176 = 0;
  assign exp_180 = exp_128 ^ exp_129;
  assign exp_184 = exp_183[31:0];
  assign exp_183 = $signed(exp_181) >>> $signed(exp_182);
  assign exp_181 = {exp_162, exp_128};
  reg [0:0] exp_162_reg;
  always@(*) begin
    case (exp_133)
      0:exp_162_reg <= exp_160;
      1:exp_162_reg <= exp_159;
      default:exp_162_reg <= exp_161;
    endcase
  end
  assign exp_162 = exp_162_reg;

      reg [0:0] exp_133_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_133_reg <= exp_77;
        end
      end
      assign exp_133 = exp_133_reg;
      assign exp_77 = exp_17[30:30];
  assign exp_161 = 0;
  assign exp_160 = 0;
  assign exp_159 = exp_128[31:31];
  assign exp_182 = $signed(exp_165);
  assign exp_185 = exp_128 | exp_129;
  assign exp_186 = exp_128 & exp_129;

  reg [31:0] exp_235_reg;
  always@(*) begin
    case (exp_140)
      0:exp_235_reg <= exp_225;
      1:exp_235_reg <= exp_228;
      2:exp_235_reg <= data_in;
      3:exp_235_reg <= exp_229;
      4:exp_235_reg <= exp_230;
      5:exp_235_reg <= exp_231;
      6:exp_235_reg <= exp_232;
      7:exp_235_reg <= exp_233;
      default:exp_235_reg <= exp_234;
    endcase
  end
  assign exp_235 = exp_235_reg;
  assign exp_234 = 0;
  assign exp_225 = $signed(exp_224);
  assign exp_224 = exp_223 + exp_218;
  assign exp_223 = 0;

  reg [7:0] exp_218_reg;
  always@(*) begin
    case (exp_209)
      0:exp_218_reg <= exp_213;
      1:exp_218_reg <= exp_214;
      2:exp_218_reg <= exp_215;
      3:exp_218_reg <= exp_216;
      default:exp_218_reg <= exp_217;
    endcase
  end
  assign exp_218 = exp_218_reg;
  assign exp_209 = exp_208 + exp_207;
  assign exp_208 = 0;
  assign exp_207 = exp_206[1:0];
  assign exp_206 = exp_126 + exp_205;
  assign exp_205 = $signed(exp_204);
  assign exp_204 = exp_203 + exp_202;
  assign exp_203 = 0;

  reg [11:0] exp_202_reg;
  always@(*) begin
    case (exp_156)
      0:exp_202_reg <= exp_197;
      1:exp_202_reg <= exp_200;
      default:exp_202_reg <= exp_201;
    endcase
  end
  assign exp_202 = exp_202_reg;
  assign exp_201 = 0;
  assign exp_197 = exp_134[31:20];
  assign exp_200 = {exp_198, exp_199};  assign exp_198 = exp_134[31:25];
  assign exp_199 = exp_134[11:7];
  assign exp_217 = 0;
  assign exp_213 = data_in[7:0];
  assign exp_214 = data_in[15:8];
  assign exp_215 = data_in[23:16];
  assign exp_216 = data_in[31:24];
  assign exp_228 = $signed(exp_227);
  assign exp_227 = exp_226 + exp_222;
  assign exp_226 = 0;

  reg [15:0] exp_222_reg;
  always@(*) begin
    case (exp_212)
      0:exp_222_reg <= exp_219;
      1:exp_222_reg <= exp_220;
      default:exp_222_reg <= exp_221;
    endcase
  end
  assign exp_222 = exp_222_reg;
  assign exp_212 = exp_211 + exp_210;
  assign exp_211 = 0;
  assign exp_210 = exp_206[1:1];
  assign exp_221 = 0;
  assign exp_219 = data_in[15:0];
  assign exp_220 = data_in[31:16];
  assign exp_229 = 0;
  assign exp_230 = exp_218;
  assign exp_231 = exp_222;
  assign exp_232 = 0;
  assign exp_233 = 0;
  assign exp_62 = $signed(exp_61);
  assign exp_61 = 0;

      reg [31:0] exp_127_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_127_reg <= exp_70;
        end
      end
      assign exp_127 = exp_127_reg;
      assign exp_290 = exp_126 != exp_127;
  assign exp_303 = 0;
  assign exp_304 = 0;
  assign exp_291 = $signed(exp_126) < $signed(exp_127);
  assign exp_292 = $signed(exp_126) >= $signed(exp_127);
  assign exp_297 = exp_294 < exp_296;
  assign exp_294 = exp_293 + exp_126;
  assign exp_293 = 0;
  assign exp_296 = exp_295 + exp_127;
  assign exp_295 = 0;
  assign exp_302 = exp_299 >= exp_301;
  assign exp_299 = exp_298 + exp_126;
  assign exp_298 = 0;
  assign exp_301 = exp_300 + exp_127;
  assign exp_300 = 0;
  assign exp_361 = 0;
  assign exp_360 = exp_12 + exp_359;
  assign exp_359 = 4;

  reg [31:0] exp_344_reg;
  always@(*) begin
    case (exp_152)
      0:exp_344_reg <= exp_337;
      1:exp_344_reg <= exp_342;
      default:exp_344_reg <= exp_343;
    endcase
  end
  assign exp_344 = exp_344_reg;
  assign exp_343 = 0;
  assign exp_337 = exp_336 + exp_135;

  reg [31:0] exp_336_reg;
  always@(*) begin
    case (exp_150)
      0:exp_336_reg <= exp_322;
      1:exp_336_reg <= exp_334;
      default:exp_336_reg <= exp_335;
    endcase
  end
  assign exp_336 = exp_336_reg;
  assign exp_335 = 0;
  assign exp_322 = $signed(exp_321);
  assign exp_321 = exp_320 + exp_319;
  assign exp_320 = 0;
  assign exp_319 = {exp_318, exp_315};  assign exp_318 = {exp_317, exp_314};  assign exp_317 = {exp_316, exp_313};  assign exp_316 = {exp_311, exp_312};  assign exp_311 = exp_134[31:31];
  assign exp_312 = exp_134[7:7];
  assign exp_313 = exp_134[30:25];
  assign exp_314 = exp_134[11:8];
  assign exp_315 = 0;
  assign exp_334 = $signed(exp_333);
  assign exp_333 = exp_332 + exp_331;
  assign exp_332 = 0;
  assign exp_331 = {exp_330, exp_327};  assign exp_330 = {exp_329, exp_326};  assign exp_329 = {exp_328, exp_325};  assign exp_328 = {exp_323, exp_324};  assign exp_323 = exp_134[31:31];
  assign exp_324 = exp_134[19:12];
  assign exp_325 = exp_134[20:20];
  assign exp_326 = exp_134[30:21];
  assign exp_327 = 0;

      reg [31:0] exp_135_reg = 0;
      always@(posedge clk) begin
        if (exp_125) begin
          exp_135_reg <= exp_18;
        end
      end
      assign exp_135 = exp_135_reg;
      assign exp_342 = exp_126 + exp_341;
  assign exp_341 = $signed(exp_340);
  assign exp_340 = exp_339 + exp_338;
  assign exp_339 = 0;
  assign exp_338 = exp_134[11:0];
  assign exp_11 = exp_4 & exp_2;
  assign exp_13 = 2;
  assign exp_267 = 0;

  reg [31:0] exp_255_reg;
  always@(*) begin
    case (exp_209)
      0:exp_255_reg <= exp_241;
      1:exp_255_reg <= exp_249;
      2:exp_255_reg <= exp_251;
      3:exp_255_reg <= exp_253;
      default:exp_255_reg <= exp_254;
    endcase
  end
  assign exp_255 = exp_255_reg;
  assign exp_254 = 0;
  assign exp_241 = exp_240;
  assign exp_240 = exp_239 + exp_238;
  assign exp_239 = 0;
  assign exp_238 = exp_127[7:0];
  assign exp_249 = exp_241 << exp_248;
  assign exp_248 = 8;
  assign exp_251 = exp_241 << exp_250;
  assign exp_250 = 16;
  assign exp_253 = exp_241 << exp_252;
  assign exp_252 = 24;

  reg [31:0] exp_259_reg;
  always@(*) begin
    case (exp_212)
      0:exp_259_reg <= exp_245;
      1:exp_259_reg <= exp_257;
      default:exp_259_reg <= exp_258;
    endcase
  end
  assign exp_259 = exp_259_reg;
  assign exp_258 = 0;
  assign exp_245 = exp_244;
  assign exp_244 = exp_243 + exp_242;
  assign exp_243 = 0;
  assign exp_242 = exp_127[15:0];
  assign exp_257 = exp_245 << exp_256;
  assign exp_256 = 16;
  assign exp_261 = exp_260 + exp_247;
  assign exp_260 = 0;
  assign exp_247 = exp_246 + exp_127;
  assign exp_246 = 0;
  assign exp_262 = 0;
  assign exp_263 = 0;
  assign exp_264 = 0;
  assign exp_265 = 0;
  assign exp_266 = 0;

  reg [3:0] exp_286_reg;
  always@(*) begin
    case (exp_140)
      0:exp_286_reg <= exp_273;
      1:exp_286_reg <= exp_278;
      2:exp_286_reg <= exp_279;
      3:exp_286_reg <= exp_280;
      4:exp_286_reg <= exp_281;
      5:exp_286_reg <= exp_282;
      6:exp_286_reg <= exp_283;
      7:exp_286_reg <= exp_284;
      default:exp_286_reg <= exp_285;
    endcase
  end
  assign exp_286 = exp_286_reg;
  assign exp_285 = 0;
  assign exp_273 = exp_269 << exp_272;
  assign exp_269 = 1;
  assign exp_272 = exp_271 + exp_270;
  assign exp_271 = 0;
  assign exp_270 = exp_206[1:0];
  assign exp_278 = exp_274 << exp_277;
  assign exp_274 = 3;
  assign exp_277 = exp_276 + exp_275;
  assign exp_276 = 0;
  assign exp_275 = exp_206[1:1];
  assign exp_279 = 15;
  assign exp_280 = 0;
  assign exp_281 = 0;
  assign exp_282 = 0;
  assign exp_283 = 0;
  assign exp_284 = 0;
  assign data_out = exp_268;
  assign address = exp_206;
  assign byte_enable = exp_286;
  assign data_valid = exp_287;
  assign write_read = exp_156;

endmodule
