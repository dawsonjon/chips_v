
module test(clk, stdout_ready_in, spare_ready_in, stdout_valid_out, stdout_out, spare_valid_out, spare_out);
  input [0:0] stdout_ready_in;
  input [0:0] spare_ready_in;
  input [0:0] clk;
  output [0:0] stdout_valid_out;
  output [31:0] stdout_out;
  output [0:0] spare_valid_out;
  output [31:0] spare_out;
  wire [0:0] exp_193;
  wire [0:0] exp_177;
  wire [0:0] exp_185;
  wire [0:0] exp_5;
  wire [0:0] exp_221;
  wire [0:0] exp_505;
  wire [0:0] exp_370;
  wire [6:0] exp_355;
  wire [31:0] exp_353;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [19:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_235;
  wire [32:0] exp_837;
  wire [0:0] exp_833;
  wire [0:0] exp_530;
  wire [0:0] exp_508;
  wire [0:0] exp_366;
  wire [6:0] exp_365;
  wire [0:0] exp_368;
  wire [6:0] exp_367;
  wire [0:0] exp_529;
  wire [0:0] exp_374;
  wire [6:0] exp_373;
  wire [0:0] exp_528;
  wire [0:0] exp_527;
  wire [0:0] exp_526;
  wire [2:0] exp_356;
  wire [0:0] exp_525;
  wire [0:0] exp_509;
  wire [31:0] exp_345;
  wire [31:0] exp_283;
  wire [0:0] exp_279;
  wire [4:0] exp_259;
  wire [0:0] exp_278;
  wire [0:0] exp_282;
  wire [31:0] exp_275;
  wire [0:0] exp_256;
  wire [0:0] exp_828;
  wire [0:0] exp_827;
  wire [0:0] exp_826;
  wire [0:0] exp_825;
  wire [4:0] exp_238;
  wire [4:0] exp_820;
  wire [0:0] exp_819;
  wire [0:0] exp_412;
  wire [0:0] exp_411;
  wire [0:0] exp_410;
  wire [0:0] exp_409;
  wire [0:0] exp_408;
  wire [0:0] exp_407;
  wire [0:0] exp_358;
  wire [4:0] exp_357;
  wire [0:0] exp_360;
  wire [5:0] exp_359;
  wire [0:0] exp_362;
  wire [5:0] exp_361;
  wire [0:0] exp_364;
  wire [4:0] exp_363;
  wire [0:0] exp_814;
  wire [0:0] exp_813;
  wire [0:0] exp_599;
  wire [0:0] exp_573;
  wire [0:0] exp_571;
  wire [6:0] exp_569;
  wire [5:0] exp_570;
  wire [0:0] exp_572;
  wire [0:0] exp_598;
  wire [2:0] exp_568;
  wire [0:0] exp_812;
  wire [0:0] exp_810;
  wire [0:0] exp_803;
  wire [2:0] exp_718;
  wire [2:0] exp_725;
  wire [0:0] exp_720;
  wire [2:0] exp_719;
  wire [0:0] exp_724;
  wire [2:0] exp_722;
  wire [0:0] exp_721;
  wire [0:0] exp_723;
  wire [0:0] exp_714;
  wire [0:0] exp_713;
  wire [0:0] exp_712;
  wire [2:0] exp_802;
  wire [0:0] exp_811;
  wire [0:0] exp_621;
  wire [5:0] exp_605;
  wire [5:0] exp_612;
  wire [0:0] exp_607;
  wire [5:0] exp_606;
  wire [0:0] exp_611;
  wire [5:0] exp_609;
  wire [0:0] exp_608;
  wire [0:0] exp_610;
  wire [5:0] exp_620;
  wire [0:0] exp_233;
  wire [0:0] exp_232;
  wire [0:0] exp_230;
  wire [0:0] exp_229;
  wire [0:0] exp_227;
  wire [0:0] exp_228;
  wire [0:0] exp_226;
  wire [0:0] exp_838;
  wire [0:0] exp_225;
  wire [0:0] exp_224;
  wire [0:0] exp_842;
  wire [0:0] exp_841;
  wire [0:0] exp_840;
  wire [0:0] exp_839;
  wire [0:0] exp_220;
  wire [0:0] exp_211;
  wire [0:0] exp_206;
  wire [0:0] exp_203;
  wire [31:0] exp_1;
  wire [31:0] exp_217;
  wire [31:0] exp_424;
  wire [31:0] exp_423;
  wire [31:0] exp_422;
  wire [31:0] exp_421;
  wire [11:0] exp_420;
  wire [11:0] exp_419;
  wire [11:0] exp_418;
  wire [0:0] exp_372;
  wire [5:0] exp_371;
  wire [0:0] exp_417;
  wire [11:0] exp_413;
  wire [11:0] exp_416;
  wire [6:0] exp_414;
  wire [4:0] exp_415;
  wire [31:0] exp_202;
  wire [0:0] exp_205;
  wire [31:0] exp_204;
  wire [0:0] exp_210;
  wire [0:0] exp_189;
  wire [0:0] exp_184;
  wire [0:0] exp_181;
  wire [31:0] exp_180;
  wire [0:0] exp_183;
  wire [31:0] exp_182;
  wire [0:0] exp_188;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [31:0] exp_146;
  wire [0:0] exp_149;
  wire [31:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [21:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_222;
  wire [0:0] exp_507;
  wire [0:0] exp_506;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_167;
  wire [0:0] exp_176;
  wire [0:0] exp_191;
  wire [0:0] exp_198;
  wire [0:0] exp_213;
  wire [0:0] exp_816;
  wire [0:0] exp_815;
  wire [0:0] exp_231;
  wire [0:0] exp_274;
  wire [31:0] exp_246;
  wire [0:0] exp_245;
  wire [1:0] exp_254;
  wire [4:0] exp_241;
  wire [0:0] exp_244;
  wire [0:0] exp_822;
  wire [0:0] exp_821;
  wire [4:0] exp_240;
  wire [31:0] exp_242;
  wire [31:0] exp_818;
  wire [0:0] exp_817;
  wire [31:0] exp_455;
  wire [0:0] exp_454;
  wire [31:0] exp_406;
  wire [2:0] exp_349;
  wire [2:0] exp_340;
  wire [0:0] exp_337;
  wire [0:0] exp_271;
  wire [6:0] exp_261;
  wire [6:0] exp_270;
  wire [0:0] exp_273;
  wire [6:0] exp_272;
  wire [0:0] exp_339;
  wire [2:0] exp_327;
  wire [0:0] exp_269;
  wire [4:0] exp_268;
  wire [0:0] exp_326;
  wire [2:0] exp_314;
  wire [0:0] exp_267;
  wire [5:0] exp_266;
  wire [0:0] exp_313;
  wire [2:0] exp_263;
  wire [0:0] exp_312;
  wire [0:0] exp_325;
  wire [0:0] exp_338;
  wire [0:0] exp_344;
  wire [0:0] exp_405;
  wire [31:0] exp_385;
  wire [0:0] exp_351;
  wire [0:0] exp_343;
  wire [0:0] exp_329;
  wire [0:0] exp_316;
  wire [0:0] exp_302;
  wire [0:0] exp_300;
  wire [0:0] exp_301;
  wire [0:0] exp_265;
  wire [4:0] exp_264;
  wire [0:0] exp_315;
  wire [0:0] exp_328;
  wire [0:0] exp_342;
  wire [0:0] exp_341;
  wire [0:0] exp_384;
  wire [31:0] exp_382;
  wire [31:0] exp_347;
  wire [31:0] exp_333;
  wire [0:0] exp_330;
  wire [0:0] exp_332;
  wire [31:0] exp_322;
  wire [0:0] exp_321;
  wire [31:0] exp_308;
  wire [0:0] exp_307;
  wire [31:0] exp_306;
  wire [31:0] exp_304;
  wire [19:0] exp_303;
  wire [3:0] exp_305;
  wire [31:0] exp_320;
  wire [31:0] exp_318;
  wire [19:0] exp_317;
  wire [3:0] exp_319;
  wire [31:0] exp_331;
  wire [31:0] exp_348;
  wire [31:0] exp_336;
  wire [0:0] exp_334;
  wire [0:0] exp_335;
  wire [31:0] exp_324;
  wire [0:0] exp_323;
  wire [31:0] exp_311;
  wire [0:0] exp_310;
  wire [31:0] exp_295;
  wire [0:0] exp_294;
  wire [31:0] exp_289;
  wire [0:0] exp_285;
  wire [4:0] exp_260;
  wire [0:0] exp_284;
  wire [0:0] exp_288;
  wire [31:0] exp_277;
  wire [0:0] exp_257;
  wire [0:0] exp_832;
  wire [0:0] exp_831;
  wire [0:0] exp_830;
  wire [0:0] exp_829;
  wire [4:0] exp_239;
  wire [0:0] exp_276;
  wire [31:0] exp_253;
  wire [0:0] exp_252;
  wire [1:0] exp_255;
  wire [4:0] exp_248;
  wire [0:0] exp_251;
  wire [0:0] exp_824;
  wire [0:0] exp_823;
  wire [4:0] exp_247;
  wire [31:0] exp_249;
  wire [31:0] exp_258;
  wire [31:0] exp_287;
  wire [0:0] exp_286;
  wire [31:0] exp_293;
  wire [31:0] exp_290;
  wire [31:0] exp_292;
  wire [11:0] exp_291;
  wire [31:0] exp_309;
  wire [31:0] exp_237;
  wire [0:0] exp_236;
  wire [31:0] exp_383;
  wire [31:0] exp_387;
  wire [31:0] exp_386;
  wire [5:0] exp_381;
  wire [5:0] exp_380;
  wire [5:0] exp_379;
  wire [4:0] exp_350;
  wire [4:0] exp_299;
  wire [0:0] exp_298;
  wire [4:0] exp_297;
  wire [4:0] exp_262;
  wire [31:0] exp_403;
  wire [1:0] exp_389;
  wire [0:0] exp_388;
  wire [31:0] exp_404;
  wire [1:0] exp_395;
  wire [0:0] exp_394;
  wire [31:0] exp_391;
  wire [31:0] exp_390;
  wire [31:0] exp_393;
  wire [31:0] exp_392;
  wire [31:0] exp_396;
  wire [31:0] exp_400;
  wire [32:0] exp_399;
  wire [32:0] exp_397;
  wire [0:0] exp_378;
  wire [0:0] exp_352;
  wire [0:0] exp_296;
  wire [0:0] exp_377;
  wire [0:0] exp_376;
  wire [0:0] exp_375;
  wire [32:0] exp_398;
  wire [31:0] exp_401;
  wire [31:0] exp_402;
  wire [31:0] exp_453;
  wire [0:0] exp_452;
  wire [31:0] exp_443;
  wire [7:0] exp_442;
  wire [7:0] exp_441;
  wire [7:0] exp_436;
  wire [1:0] exp_427;
  wire [1:0] exp_426;
  wire [1:0] exp_425;
  wire [0:0] exp_435;
  wire [7:0] exp_431;
  wire [31:0] exp_219;
  wire [31:0] exp_209;
  wire [0:0] exp_208;
  wire [31:0] exp_187;
  wire [0:0] exp_186;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [19:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_223;
  wire [3:0] exp_504;
  wire [0:0] exp_503;
  wire [3:0] exp_491;
  wire [3:0] exp_487;
  wire [1:0] exp_490;
  wire [1:0] exp_489;
  wire [1:0] exp_488;
  wire [3:0] exp_496;
  wire [3:0] exp_492;
  wire [0:0] exp_495;
  wire [0:0] exp_494;
  wire [0:0] exp_493;
  wire [3:0] exp_497;
  wire [3:0] exp_498;
  wire [3:0] exp_499;
  wire [3:0] exp_500;
  wire [3:0] exp_501;
  wire [3:0] exp_502;
  wire [19:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_218;
  wire [31:0] exp_486;
  wire [0:0] exp_485;
  wire [31:0] exp_473;
  wire [0:0] exp_472;
  wire [31:0] exp_459;
  wire [7:0] exp_458;
  wire [7:0] exp_457;
  wire [7:0] exp_456;
  wire [31:0] exp_346;
  wire [31:0] exp_467;
  wire [3:0] exp_466;
  wire [31:0] exp_469;
  wire [4:0] exp_468;
  wire [31:0] exp_471;
  wire [4:0] exp_470;
  wire [31:0] exp_477;
  wire [0:0] exp_430;
  wire [0:0] exp_429;
  wire [0:0] exp_428;
  wire [0:0] exp_476;
  wire [31:0] exp_463;
  wire [15:0] exp_462;
  wire [15:0] exp_461;
  wire [15:0] exp_460;
  wire [31:0] exp_475;
  wire [4:0] exp_474;
  wire [31:0] exp_479;
  wire [31:0] exp_478;
  wire [31:0] exp_465;
  wire [31:0] exp_464;
  wire [31:0] exp_480;
  wire [31:0] exp_481;
  wire [31:0] exp_482;
  wire [31:0] exp_483;
  wire [31:0] exp_484;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [19:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [19:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [19:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [19:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [19:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [19:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [19:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [19:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [19:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [19:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [19:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [19:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_172;
  wire [0:0] exp_168;
  wire [31:0] exp_139;
  wire [0:0] exp_171;
  wire [31:0] exp_169;
  wire [63:0] exp_157;
  wire [63:0] exp_164;
  wire [0:0] exp_159;
  wire [63:0] exp_158;
  wire [0:0] exp_163;
  wire [63:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [31:0] exp_170;
  wire [31:0] exp_175;
  wire [31:0] exp_194;
  wire [31:0] exp_197;
  wire [31:0] exp_216;
  wire [7:0] exp_432;
  wire [7:0] exp_433;
  wire [7:0] exp_434;
  wire [31:0] exp_446;
  wire [15:0] exp_445;
  wire [15:0] exp_444;
  wire [15:0] exp_440;
  wire [0:0] exp_439;
  wire [15:0] exp_437;
  wire [15:0] exp_438;
  wire [31:0] exp_447;
  wire [31:0] exp_448;
  wire [31:0] exp_449;
  wire [31:0] exp_450;
  wire [31:0] exp_451;
  wire [31:0] exp_809;
  wire [0:0] exp_808;
  wire [31:0] exp_805;
  wire [0:0] exp_576;
  wire [0:0] exp_575;
  wire [0:0] exp_574;
  wire [0:0] exp_804;
  wire [31:0] exp_800;
  wire [63:0] exp_799;
  wire [0:0] exp_796;
  wire [0:0] exp_779;
  wire [0:0] exp_756;
  wire [0:0] exp_753;
  wire [0:0] exp_751;
  wire [0:0] exp_733;
  wire [0:0] exp_732;
  wire [0:0] exp_731;
  wire [31:0] exp_729;
  wire [0:0] exp_728;
  wire [0:0] exp_727;
  wire [0:0] exp_716;
  wire [0:0] exp_715;
  wire [0:0] exp_579;
  wire [0:0] exp_578;
  wire [0:0] exp_577;
  wire [0:0] exp_582;
  wire [0:0] exp_581;
  wire [1:0] exp_580;
  wire [0:0] exp_752;
  wire [0:0] exp_736;
  wire [0:0] exp_735;
  wire [0:0] exp_734;
  wire [31:0] exp_730;
  wire [0:0] exp_717;
  wire [0:0] exp_738;
  wire [0:0] exp_737;
  wire [0:0] exp_758;
  wire [1:0] exp_757;
  wire [0:0] exp_781;
  wire [1:0] exp_780;
  wire [0:0] exp_798;
  wire [63:0] exp_795;
  wire [63:0] exp_794;
  wire [63:0] exp_790;
  wire [63:0] exp_786;
  wire [63:0] exp_782;
  wire [31:0] exp_775;
  wire [31:0] exp_762;
  wire [31:0] exp_760;
  wire [15:0] exp_759;
  wire [31:0] exp_754;
  wire [31:0] exp_744;
  wire [31:0] exp_743;
  wire [31:0] exp_742;
  wire [0:0] exp_739;
  wire [0:0] exp_741;
  wire [31:0] exp_740;
  wire [15:0] exp_761;
  wire [31:0] exp_755;
  wire [31:0] exp_750;
  wire [31:0] exp_749;
  wire [31:0] exp_748;
  wire [0:0] exp_745;
  wire [0:0] exp_747;
  wire [31:0] exp_746;
  wire [63:0] exp_785;
  wire [63:0] exp_783;
  wire [31:0] exp_776;
  wire [31:0] exp_766;
  wire [31:0] exp_764;
  wire [15:0] exp_763;
  wire [15:0] exp_765;
  wire [4:0] exp_784;
  wire [63:0] exp_789;
  wire [63:0] exp_787;
  wire [31:0] exp_777;
  wire [31:0] exp_770;
  wire [31:0] exp_768;
  wire [15:0] exp_767;
  wire [15:0] exp_769;
  wire [4:0] exp_788;
  wire [63:0] exp_793;
  wire [63:0] exp_791;
  wire [31:0] exp_778;
  wire [31:0] exp_774;
  wire [31:0] exp_772;
  wire [15:0] exp_771;
  wire [15:0] exp_773;
  wire [5:0] exp_792;
  wire [63:0] exp_797;
  wire [31:0] exp_801;
  wire [31:0] exp_807;
  wire [0:0] exp_600;
  wire [0:0] exp_806;
  wire [31:0] exp_710;
  wire [31:0] exp_704;
  wire [0:0] exp_700;
  wire [0:0] exp_699;
  wire [31:0] exp_648;
  wire [31:0] exp_645;
  wire [31:0] exp_644;
  wire [31:0] exp_643;
  wire [0:0] exp_640;
  wire [0:0] exp_631;
  wire [0:0] exp_630;
  wire [0:0] exp_629;
  wire [31:0] exp_625;
  wire [0:0] exp_623;
  wire [0:0] exp_622;
  wire [0:0] exp_602;
  wire [0:0] exp_601;
  wire [0:0] exp_642;
  wire [31:0] exp_641;
  wire [0:0] exp_633;
  wire [0:0] exp_632;
  wire [0:0] exp_698;
  wire [0:0] exp_703;
  wire [31:0] exp_691;
  wire [31:0] exp_690;
  wire [31:0] exp_689;
  wire [0:0] exp_686;
  wire [0:0] exp_650;
  wire [0:0] exp_646;
  wire [0:0] exp_628;
  wire [0:0] exp_627;
  wire [0:0] exp_626;
  wire [31:0] exp_624;
  wire [0:0] exp_688;
  wire [31:0] exp_684;
  wire [31:0] exp_654;
  wire [31:0] exp_681;
  wire [0:0] exp_615;
  wire [1:0] exp_614;
  wire [0:0] exp_680;
  wire [31:0] exp_673;
  wire [0:0] exp_663;
  wire [0:0] exp_662;
  wire [32:0] exp_661;
  wire [32:0] exp_660;
  wire [32:0] exp_659;
  wire [31:0] exp_657;
  wire [31:0] exp_652;
  wire [32:0] exp_678;
  wire [0:0] exp_677;
  wire [32:0] exp_665;
  wire [0:0] exp_664;
  wire [0:0] exp_676;
  wire [0:0] exp_651;
  wire [0:0] exp_658;
  wire [31:0] exp_656;
  wire [31:0] exp_683;
  wire [0:0] exp_682;
  wire [31:0] exp_675;
  wire [0:0] exp_674;
  wire [31:0] exp_647;
  wire [31:0] exp_639;
  wire [31:0] exp_638;
  wire [31:0] exp_637;
  wire [0:0] exp_634;
  wire [0:0] exp_636;
  wire [31:0] exp_635;
  wire [0:0] exp_655;
  wire [0:0] exp_672;
  wire [31:0] exp_667;
  wire [0:0] exp_666;
  wire [31:0] exp_671;
  wire [31:0] exp_669;
  wire [0:0] exp_668;
  wire [0:0] exp_670;
  wire [0:0] exp_679;
  wire [0:0] exp_653;
  wire [0:0] exp_617;
  wire [5:0] exp_616;
  wire [31:0] exp_687;
  wire [31:0] exp_702;
  wire [0:0] exp_701;
  wire [0:0] exp_619;
  wire [5:0] exp_618;
  wire [31:0] exp_711;
  wire [31:0] exp_709;
  wire [0:0] exp_707;
  wire [0:0] exp_706;
  wire [0:0] exp_705;
  wire [0:0] exp_708;
  wire [31:0] exp_697;
  wire [31:0] exp_696;
  wire [31:0] exp_695;
  wire [0:0] exp_692;
  wire [0:0] exp_649;
  wire [0:0] exp_694;
  wire [31:0] exp_685;
  wire [31:0] exp_693;
  wire [31:0] exp_281;
  wire [0:0] exp_280;
  wire [0:0] exp_510;
  wire [0:0] exp_523;
  wire [0:0] exp_524;
  wire [0:0] exp_511;
  wire [0:0] exp_512;
  wire [0:0] exp_517;
  wire [31:0] exp_514;
  wire [31:0] exp_513;
  wire [31:0] exp_516;
  wire [31:0] exp_515;
  wire [0:0] exp_522;
  wire [31:0] exp_519;
  wire [31:0] exp_518;
  wire [31:0] exp_521;
  wire [31:0] exp_520;
  wire [0:0] exp_836;
  wire [31:0] exp_835;
  wire [2:0] exp_834;
  wire [32:0] exp_567;
  wire [0:0] exp_566;
  wire [31:0] exp_557;
  wire [31:0] exp_556;
  wire [0:0] exp_555;
  wire [31:0] exp_542;
  wire [12:0] exp_541;
  wire [12:0] exp_540;
  wire [12:0] exp_539;
  wire [11:0] exp_538;
  wire [7:0] exp_537;
  wire [1:0] exp_536;
  wire [0:0] exp_531;
  wire [0:0] exp_532;
  wire [5:0] exp_533;
  wire [3:0] exp_534;
  wire [0:0] exp_535;
  wire [31:0] exp_554;
  wire [20:0] exp_553;
  wire [20:0] exp_552;
  wire [20:0] exp_551;
  wire [19:0] exp_550;
  wire [9:0] exp_549;
  wire [8:0] exp_548;
  wire [0:0] exp_543;
  wire [7:0] exp_544;
  wire [0:0] exp_545;
  wire [9:0] exp_546;
  wire [0:0] exp_547;
  wire [31:0] exp_354;
  wire [32:0] exp_565;
  wire [32:0] exp_564;
  wire [31:0] exp_562;
  wire [31:0] exp_561;
  wire [11:0] exp_560;
  wire [11:0] exp_559;
  wire [11:0] exp_558;
  wire [32:0] exp_563;
  wire [0:0] exp_234;
  wire [0:0] exp_80;
  wire [19:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_369;
  wire [0:0] exp_178;
  wire [31:0] exp_174;
  wire [0:0] exp_215;
  wire [0:0] exp_199;
  wire [0:0] exp_207;
  wire [0:0] exp_200;
  wire [31:0] exp_196;

  assign exp_193 = exp_177 & exp_178;
  assign exp_177 = exp_185;
  assign exp_185 = exp_5 & exp_184;
  assign exp_5 = exp_221;
  assign exp_221 = exp_505;
  assign exp_505 = exp_370 | exp_372;
  assign exp_370 = exp_355 == exp_369;
  assign exp_355 = exp_353[6:0];

      reg [31:0] exp_353_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_353_reg <= exp_96;
        end
      end
      assign exp_353 = exp_353_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};

  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_235;

      reg [31:0] exp_235_reg = 0;
      always@(posedge clk) begin
        if (exp_234) begin
          exp_235_reg <= exp_837;
        end
      end
      assign exp_235 = exp_235_reg;
    
  reg [32:0] exp_837_reg;
  always@(*) begin
    case (exp_833)
      0:exp_837_reg <= exp_835;
      1:exp_837_reg <= exp_567;
      default:exp_837_reg <= exp_836;
    endcase
  end
  assign exp_837 = exp_837_reg;
  assign exp_833 = exp_530 & exp_233;
  assign exp_530 = exp_508 | exp_529;
  assign exp_508 = exp_366 | exp_368;
  assign exp_366 = exp_355 == exp_365;
  assign exp_365 = 111;
  assign exp_368 = exp_355 == exp_367;
  assign exp_367 = 103;

  reg [0:0] exp_529_reg;
  always@(*) begin
    case (exp_374)
      0:exp_529_reg <= exp_527;
      1:exp_529_reg <= exp_526;
      default:exp_529_reg <= exp_528;
    endcase
  end
  assign exp_529 = exp_529_reg;
  assign exp_374 = exp_355 == exp_373;
  assign exp_373 = 99;
  assign exp_528 = 0;
  assign exp_527 = 0;

  reg [0:0] exp_526_reg;
  always@(*) begin
    case (exp_356)
      0:exp_526_reg <= exp_509;
      1:exp_526_reg <= exp_510;
      2:exp_526_reg <= exp_523;
      3:exp_526_reg <= exp_524;
      4:exp_526_reg <= exp_511;
      5:exp_526_reg <= exp_512;
      6:exp_526_reg <= exp_517;
      7:exp_526_reg <= exp_522;
      default:exp_526_reg <= exp_525;
    endcase
  end
  assign exp_526 = exp_526_reg;
  assign exp_356 = exp_353[14:12];
  assign exp_525 = 0;
  assign exp_509 = exp_345 == exp_346;

      reg [31:0] exp_345_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_345_reg <= exp_283;
        end
      end
      assign exp_345 = exp_345_reg;
    
  reg [31:0] exp_283_reg;
  always@(*) begin
    case (exp_279)
      0:exp_283_reg <= exp_275;
      1:exp_283_reg <= exp_281;
      default:exp_283_reg <= exp_282;
    endcase
  end
  assign exp_283 = exp_283_reg;
  assign exp_279 = exp_259 == exp_278;
  assign exp_259 = exp_96[19:15];
  assign exp_278 = 0;
  assign exp_282 = 0;

  reg [31:0] exp_275_reg;
  always@(*) begin
    case (exp_256)
      0:exp_275_reg <= exp_246;
      1:exp_275_reg <= exp_258;
      default:exp_275_reg <= exp_274;
    endcase
  end
  assign exp_275 = exp_275_reg;
  assign exp_256 = exp_828;
  assign exp_828 = exp_827 & exp_225;
  assign exp_827 = exp_826 & exp_233;
  assign exp_826 = exp_825 & exp_819;
  assign exp_825 = exp_238 == exp_820;
  assign exp_238 = exp_96[19:15];
  assign exp_820 = exp_353[11:7];
  assign exp_819 = exp_412 | exp_814;
  assign exp_412 = exp_411 | exp_370;
  assign exp_411 = exp_410 | exp_364;
  assign exp_410 = exp_409 | exp_362;
  assign exp_409 = exp_408 | exp_368;
  assign exp_408 = exp_407 | exp_366;
  assign exp_407 = exp_358 | exp_360;
  assign exp_358 = exp_355 == exp_357;
  assign exp_357 = 19;
  assign exp_360 = exp_355 == exp_359;
  assign exp_359 = 51;
  assign exp_362 = exp_355 == exp_361;
  assign exp_361 = 55;
  assign exp_364 = exp_355 == exp_363;
  assign exp_363 = 23;
  assign exp_814 = exp_813 & exp_573;

  reg [0:0] exp_813_reg;
  always@(*) begin
    case (exp_599)
      0:exp_813_reg <= exp_810;
      1:exp_813_reg <= exp_811;
      default:exp_813_reg <= exp_812;
    endcase
  end
  assign exp_813 = exp_813_reg;
  assign exp_599 = exp_573 & exp_598;
  assign exp_573 = exp_571 & exp_572;
  assign exp_571 = exp_569 == exp_570;
  assign exp_569 = exp_353[6:0];
  assign exp_570 = 51;
  assign exp_572 = exp_353[25:25];
  assign exp_598 = exp_568[2:2];
  assign exp_568 = exp_353[14:12];
  assign exp_812 = 0;
  assign exp_810 = exp_803 & exp_573;
  assign exp_803 = exp_718 == exp_802;

      reg [2:0] exp_718_reg = 0;
      always@(posedge clk) begin
        if (exp_714) begin
          exp_718_reg <= exp_725;
        end
      end
      assign exp_718 = exp_718_reg;
    
  reg [2:0] exp_725_reg;
  always@(*) begin
    case (exp_720)
      0:exp_725_reg <= exp_722;
      1:exp_725_reg <= exp_723;
      default:exp_725_reg <= exp_724;
    endcase
  end
  assign exp_725 = exp_725_reg;
  assign exp_720 = exp_718 == exp_719;
  assign exp_719 = 4;
  assign exp_724 = 0;
  assign exp_722 = exp_718 + exp_721;
  assign exp_721 = 1;
  assign exp_723 = 0;
  assign exp_714 = exp_573 & exp_713;
  assign exp_713 = ~exp_712;
  assign exp_712 = exp_568[2:2];
  assign exp_802 = 4;
  assign exp_811 = exp_621 & exp_573;
  assign exp_621 = exp_605 == exp_620;

      reg [5:0] exp_605_reg = 0;
      always@(posedge clk) begin
        if (exp_599) begin
          exp_605_reg <= exp_612;
        end
      end
      assign exp_605 = exp_605_reg;
    
  reg [5:0] exp_612_reg;
  always@(*) begin
    case (exp_607)
      0:exp_612_reg <= exp_609;
      1:exp_612_reg <= exp_610;
      default:exp_612_reg <= exp_611;
    endcase
  end
  assign exp_612 = exp_612_reg;
  assign exp_607 = exp_605 == exp_606;
  assign exp_606 = 37;
  assign exp_611 = 0;
  assign exp_609 = exp_605 + exp_608;
  assign exp_608 = 1;
  assign exp_610 = 0;
  assign exp_620 = 37;

      reg [0:0] exp_233_reg = 0;
      always@(posedge clk) begin
        if (exp_225) begin
          exp_233_reg <= exp_232;
        end
      end
      assign exp_233 = exp_233_reg;
      assign exp_232 = exp_230 & exp_231;

      reg [0:0] exp_230_reg = 0;
      always@(posedge clk) begin
        if (exp_225) begin
          exp_230_reg <= exp_229;
        end
      end
      assign exp_230 = exp_230_reg;
      assign exp_229 = exp_227 & exp_228;
  assign exp_227 = 1;
  assign exp_228 = ~exp_226;
  assign exp_226 = exp_838;
  assign exp_838 = exp_233 & exp_530;
  assign exp_225 = ~exp_224;
  assign exp_224 = exp_842;
  assign exp_842 = exp_233 & exp_841;
  assign exp_841 = exp_840 | exp_816;
  assign exp_840 = exp_221 & exp_839;
  assign exp_839 = ~exp_220;
  assign exp_220 = exp_211;

  reg [0:0] exp_211_reg;
  always@(*) begin
    case (exp_206)
      0:exp_211_reg <= exp_189;
      1:exp_211_reg <= exp_198;
      default:exp_211_reg <= exp_210;
    endcase
  end
  assign exp_211 = exp_211_reg;
  assign exp_206 = exp_203 & exp_205;
  assign exp_203 = exp_1 >= exp_202;
  assign exp_1 = exp_217;
  assign exp_217 = exp_424;
  assign exp_424 = exp_423 + exp_422;
  assign exp_423 = 0;
  assign exp_422 = exp_345 + exp_421;
  assign exp_421 = $signed(exp_420);
  assign exp_420 = exp_419 + exp_418;
  assign exp_419 = 0;

  reg [11:0] exp_418_reg;
  always@(*) begin
    case (exp_372)
      0:exp_418_reg <= exp_413;
      1:exp_418_reg <= exp_416;
      default:exp_418_reg <= exp_417;
    endcase
  end
  assign exp_418 = exp_418_reg;
  assign exp_372 = exp_355 == exp_371;
  assign exp_371 = 35;
  assign exp_417 = 0;
  assign exp_413 = exp_353[31:20];
  assign exp_416 = {exp_414, exp_415};  assign exp_414 = exp_353[31:25];
  assign exp_415 = exp_353[11:7];
  assign exp_202 = 2147483660;
  assign exp_205 = exp_1 <= exp_204;
  assign exp_204 = 2147483660;
  assign exp_210 = 0;

  reg [0:0] exp_189_reg;
  always@(*) begin
    case (exp_184)
      0:exp_189_reg <= exp_155;
      1:exp_189_reg <= exp_176;
      default:exp_189_reg <= exp_188;
    endcase
  end
  assign exp_189 = exp_189_reg;
  assign exp_184 = exp_181 & exp_183;
  assign exp_181 = exp_1 >= exp_180;
  assign exp_180 = 2147483656;
  assign exp_183 = exp_1 <= exp_182;
  assign exp_182 = 2147483656;
  assign exp_188 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 2147483648;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 2147483652;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 4194300;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_222;
  assign exp_222 = exp_507;
  assign exp_507 = exp_506 + exp_372;
  assign exp_506 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_167;
  assign exp_167 = 1;
  assign exp_176 = exp_191;
  assign exp_191 = stdout_ready_in;
  assign exp_198 = exp_213;
  assign exp_213 = spare_ready_in;
  assign exp_816 = exp_573 & exp_815;
  assign exp_815 = ~exp_813;
  assign exp_231 = ~exp_226;
  assign exp_274 = 0;

  //Create RAM
  reg [31:0] exp_246_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_244) begin
      exp_246_ram[exp_240] <= exp_242;
    end
  end
  assign exp_246 = exp_246_ram[exp_241];
  assign exp_245 = exp_254;
  assign exp_254 = 1;
  assign exp_241 = exp_238;
  assign exp_244 = exp_822;
  assign exp_822 = exp_821 & exp_225;
  assign exp_821 = exp_819 & exp_233;
  assign exp_240 = exp_820;
  assign exp_242 = exp_818;

  reg [31:0] exp_818_reg;
  always@(*) begin
    case (exp_814)
      0:exp_818_reg <= exp_455;
      1:exp_818_reg <= exp_809;
      default:exp_818_reg <= exp_817;
    endcase
  end
  assign exp_818 = exp_818_reg;
  assign exp_817 = 0;

  reg [31:0] exp_455_reg;
  always@(*) begin
    case (exp_370)
      0:exp_455_reg <= exp_406;
      1:exp_455_reg <= exp_453;
      default:exp_455_reg <= exp_454;
    endcase
  end
  assign exp_455 = exp_455_reg;
  assign exp_454 = 0;

  reg [31:0] exp_406_reg;
  always@(*) begin
    case (exp_349)
      0:exp_406_reg <= exp_385;
      1:exp_406_reg <= exp_387;
      2:exp_406_reg <= exp_403;
      3:exp_406_reg <= exp_404;
      4:exp_406_reg <= exp_396;
      5:exp_406_reg <= exp_400;
      6:exp_406_reg <= exp_401;
      7:exp_406_reg <= exp_402;
      default:exp_406_reg <= exp_405;
    endcase
  end
  assign exp_406 = exp_406_reg;

      reg [2:0] exp_349_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_349_reg <= exp_340;
        end
      end
      assign exp_349 = exp_349_reg;
    
  reg [2:0] exp_340_reg;
  always@(*) begin
    case (exp_337)
      0:exp_340_reg <= exp_327;
      1:exp_340_reg <= exp_338;
      default:exp_340_reg <= exp_339;
    endcase
  end
  assign exp_340 = exp_340_reg;
  assign exp_337 = exp_271 | exp_273;
  assign exp_271 = exp_261 == exp_270;
  assign exp_261 = exp_96[6:0];
  assign exp_270 = 111;
  assign exp_273 = exp_261 == exp_272;
  assign exp_272 = 103;
  assign exp_339 = 0;

  reg [2:0] exp_327_reg;
  always@(*) begin
    case (exp_269)
      0:exp_327_reg <= exp_314;
      1:exp_327_reg <= exp_325;
      default:exp_327_reg <= exp_326;
    endcase
  end
  assign exp_327 = exp_327_reg;
  assign exp_269 = exp_261 == exp_268;
  assign exp_268 = 23;
  assign exp_326 = 0;

  reg [2:0] exp_314_reg;
  always@(*) begin
    case (exp_267)
      0:exp_314_reg <= exp_263;
      1:exp_314_reg <= exp_312;
      default:exp_314_reg <= exp_313;
    endcase
  end
  assign exp_314 = exp_314_reg;
  assign exp_267 = exp_261 == exp_266;
  assign exp_266 = 55;
  assign exp_313 = 0;
  assign exp_263 = exp_96[14:12];
  assign exp_312 = 0;
  assign exp_325 = 0;
  assign exp_338 = 0;
  assign exp_344 = exp_225 & exp_230;
  assign exp_405 = 0;

  reg [31:0] exp_385_reg;
  always@(*) begin
    case (exp_351)
      0:exp_385_reg <= exp_382;
      1:exp_385_reg <= exp_383;
      default:exp_385_reg <= exp_384;
    endcase
  end
  assign exp_385 = exp_385_reg;

      reg [0:0] exp_351_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_351_reg <= exp_343;
        end
      end
      assign exp_351 = exp_351_reg;
      assign exp_343 = exp_329 & exp_342;
  assign exp_329 = exp_316 & exp_328;
  assign exp_316 = exp_302 & exp_315;
  assign exp_302 = exp_300 & exp_301;
  assign exp_300 = exp_96[30:30];
  assign exp_301 = ~exp_265;
  assign exp_265 = exp_261 == exp_264;
  assign exp_264 = 19;
  assign exp_315 = ~exp_267;
  assign exp_328 = ~exp_269;
  assign exp_342 = ~exp_341;
  assign exp_341 = exp_271 | exp_273;
  assign exp_384 = 0;
  assign exp_382 = exp_347 + exp_348;

      reg [31:0] exp_347_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_347_reg <= exp_333;
        end
      end
      assign exp_347 = exp_347_reg;
    
  reg [31:0] exp_333_reg;
  always@(*) begin
    case (exp_330)
      0:exp_333_reg <= exp_322;
      1:exp_333_reg <= exp_331;
      default:exp_333_reg <= exp_332;
    endcase
  end
  assign exp_333 = exp_333_reg;
  assign exp_330 = exp_271 | exp_273;
  assign exp_332 = 0;

  reg [31:0] exp_322_reg;
  always@(*) begin
    case (exp_269)
      0:exp_322_reg <= exp_308;
      1:exp_322_reg <= exp_320;
      default:exp_322_reg <= exp_321;
    endcase
  end
  assign exp_322 = exp_322_reg;
  assign exp_321 = 0;

  reg [31:0] exp_308_reg;
  always@(*) begin
    case (exp_267)
      0:exp_308_reg <= exp_283;
      1:exp_308_reg <= exp_306;
      default:exp_308_reg <= exp_307;
    endcase
  end
  assign exp_308 = exp_308_reg;
  assign exp_307 = 0;
  assign exp_306 = exp_304 << exp_305;
  assign exp_304 = exp_303;
  assign exp_303 = exp_96[31:12];
  assign exp_305 = 12;
  assign exp_320 = exp_318 << exp_319;
  assign exp_318 = exp_317;
  assign exp_317 = exp_96[31:12];
  assign exp_319 = 12;
  assign exp_331 = 4;

      reg [31:0] exp_348_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_348_reg <= exp_336;
        end
      end
      assign exp_348 = exp_348_reg;
    
  reg [31:0] exp_336_reg;
  always@(*) begin
    case (exp_334)
      0:exp_336_reg <= exp_324;
      1:exp_336_reg <= exp_237;
      default:exp_336_reg <= exp_335;
    endcase
  end
  assign exp_336 = exp_336_reg;
  assign exp_334 = exp_271 | exp_273;
  assign exp_335 = 0;

  reg [31:0] exp_324_reg;
  always@(*) begin
    case (exp_269)
      0:exp_324_reg <= exp_311;
      1:exp_324_reg <= exp_237;
      default:exp_324_reg <= exp_323;
    endcase
  end
  assign exp_324 = exp_324_reg;
  assign exp_323 = 0;

  reg [31:0] exp_311_reg;
  always@(*) begin
    case (exp_267)
      0:exp_311_reg <= exp_295;
      1:exp_311_reg <= exp_309;
      default:exp_311_reg <= exp_310;
    endcase
  end
  assign exp_311 = exp_311_reg;
  assign exp_310 = 0;

  reg [31:0] exp_295_reg;
  always@(*) begin
    case (exp_265)
      0:exp_295_reg <= exp_289;
      1:exp_295_reg <= exp_293;
      default:exp_295_reg <= exp_294;
    endcase
  end
  assign exp_295 = exp_295_reg;
  assign exp_294 = 0;

  reg [31:0] exp_289_reg;
  always@(*) begin
    case (exp_285)
      0:exp_289_reg <= exp_277;
      1:exp_289_reg <= exp_287;
      default:exp_289_reg <= exp_288;
    endcase
  end
  assign exp_289 = exp_289_reg;
  assign exp_285 = exp_260 == exp_284;
  assign exp_260 = exp_96[24:20];
  assign exp_284 = 0;
  assign exp_288 = 0;

  reg [31:0] exp_277_reg;
  always@(*) begin
    case (exp_257)
      0:exp_277_reg <= exp_253;
      1:exp_277_reg <= exp_258;
      default:exp_277_reg <= exp_276;
    endcase
  end
  assign exp_277 = exp_277_reg;
  assign exp_257 = exp_832;
  assign exp_832 = exp_831 & exp_225;
  assign exp_831 = exp_830 & exp_233;
  assign exp_830 = exp_829 & exp_819;
  assign exp_829 = exp_239 == exp_820;
  assign exp_239 = exp_96[24:20];
  assign exp_276 = 0;

  //Create RAM
  reg [31:0] exp_253_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_251) begin
      exp_253_ram[exp_247] <= exp_249;
    end
  end
  assign exp_253 = exp_253_ram[exp_248];
  assign exp_252 = exp_255;
  assign exp_255 = 1;
  assign exp_248 = exp_239;
  assign exp_251 = exp_824;
  assign exp_824 = exp_823 & exp_225;
  assign exp_823 = exp_819 & exp_233;
  assign exp_247 = exp_820;
  assign exp_249 = exp_818;
  assign exp_258 = exp_818;
  assign exp_287 = $signed(exp_286);
  assign exp_286 = 0;
  assign exp_293 = exp_290 + exp_292;
  assign exp_290 = 0;
  assign exp_292 = $signed(exp_291);
  assign exp_291 = exp_96[31:20];
  assign exp_309 = 0;

      reg [31:0] exp_237_reg = 0;
      always@(posedge clk) begin
        if (exp_236) begin
          exp_237_reg <= exp_235;
        end
      end
      assign exp_237 = exp_237_reg;
      assign exp_236 = exp_227 & exp_225;
  assign exp_383 = exp_347 - exp_348;
  assign exp_387 = exp_347 << exp_386;
  assign exp_386 = $signed(exp_381);
  assign exp_381 = exp_380 + exp_379;
  assign exp_380 = 0;
  assign exp_379 = exp_350;

      reg [4:0] exp_350_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_350_reg <= exp_299;
        end
      end
      assign exp_350 = exp_350_reg;
    
  reg [4:0] exp_299_reg;
  always@(*) begin
    case (exp_265)
      0:exp_299_reg <= exp_297;
      1:exp_299_reg <= exp_262;
      default:exp_299_reg <= exp_298;
    endcase
  end
  assign exp_299 = exp_299_reg;
  assign exp_298 = 0;
  assign exp_297 = exp_295[4:0];
  assign exp_262 = exp_96[24:20];
  assign exp_403 = $signed(exp_389);
  assign exp_389 = exp_388;
  assign exp_388 = $signed(exp_347) < $signed(exp_348);
  assign exp_404 = $signed(exp_395);
  assign exp_395 = exp_394;
  assign exp_394 = exp_391 < exp_393;
  assign exp_391 = exp_390 + exp_347;
  assign exp_390 = 0;
  assign exp_393 = exp_392 + exp_348;
  assign exp_392 = 0;
  assign exp_396 = exp_347 ^ exp_348;
  assign exp_400 = exp_399[31:0];
  assign exp_399 = $signed(exp_397) >>> $signed(exp_398);
  assign exp_397 = {exp_378, exp_347};
  reg [0:0] exp_378_reg;
  always@(*) begin
    case (exp_352)
      0:exp_378_reg <= exp_376;
      1:exp_378_reg <= exp_375;
      default:exp_378_reg <= exp_377;
    endcase
  end
  assign exp_378 = exp_378_reg;

      reg [0:0] exp_352_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_352_reg <= exp_296;
        end
      end
      assign exp_352 = exp_352_reg;
      assign exp_296 = exp_96[30:30];
  assign exp_377 = 0;
  assign exp_376 = 0;
  assign exp_375 = exp_347[31:31];
  assign exp_398 = $signed(exp_381);
  assign exp_401 = exp_347 | exp_348;
  assign exp_402 = exp_347 & exp_348;

  reg [31:0] exp_453_reg;
  always@(*) begin
    case (exp_356)
      0:exp_453_reg <= exp_443;
      1:exp_453_reg <= exp_446;
      2:exp_453_reg <= exp_219;
      3:exp_453_reg <= exp_447;
      4:exp_453_reg <= exp_448;
      5:exp_453_reg <= exp_449;
      6:exp_453_reg <= exp_450;
      7:exp_453_reg <= exp_451;
      default:exp_453_reg <= exp_452;
    endcase
  end
  assign exp_453 = exp_453_reg;
  assign exp_452 = 0;
  assign exp_443 = $signed(exp_442);
  assign exp_442 = exp_441 + exp_436;
  assign exp_441 = 0;

  reg [7:0] exp_436_reg;
  always@(*) begin
    case (exp_427)
      0:exp_436_reg <= exp_431;
      1:exp_436_reg <= exp_432;
      2:exp_436_reg <= exp_433;
      3:exp_436_reg <= exp_434;
      default:exp_436_reg <= exp_435;
    endcase
  end
  assign exp_436 = exp_436_reg;
  assign exp_427 = exp_426 + exp_425;
  assign exp_426 = 0;
  assign exp_425 = exp_424[1:0];
  assign exp_435 = 0;
  assign exp_431 = exp_219[7:0];
  assign exp_219 = exp_209;

  reg [31:0] exp_209_reg;
  always@(*) begin
    case (exp_206)
      0:exp_209_reg <= exp_187;
      1:exp_209_reg <= exp_197;
      default:exp_209_reg <= exp_208;
    endcase
  end
  assign exp_209 = exp_209_reg;
  assign exp_208 = 0;

  reg [31:0] exp_187_reg;
  always@(*) begin
    case (exp_184)
      0:exp_187_reg <= exp_153;
      1:exp_187_reg <= exp_175;
      default:exp_187_reg <= exp_186;
    endcase
  end
  assign exp_187 = exp_187_reg;
  assign exp_186 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [1048575:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 0;
    exp_54_ram[32] = 255;
    exp_54_ram[33] = 3;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 0;
    exp_54_ram[36] = 0;
    exp_54_ram[37] = 0;
    exp_54_ram[38] = 0;
    exp_54_ram[39] = 0;
    exp_54_ram[40] = 0;
    exp_54_ram[41] = 0;
    exp_54_ram[42] = 0;
    exp_54_ram[43] = 254;
    exp_54_ram[44] = 128;
    exp_54_ram[45] = 0;
    exp_54_ram[46] = 253;
    exp_54_ram[47] = 12;
    exp_54_ram[48] = 255;
    exp_54_ram[49] = 108;
    exp_54_ram[50] = 111;
    exp_54_ram[51] = 33;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_223;
  assign exp_223 = exp_504;

  reg [3:0] exp_504_reg;
  always@(*) begin
    case (exp_356)
      0:exp_504_reg <= exp_491;
      1:exp_504_reg <= exp_496;
      2:exp_504_reg <= exp_497;
      3:exp_504_reg <= exp_498;
      4:exp_504_reg <= exp_499;
      5:exp_504_reg <= exp_500;
      6:exp_504_reg <= exp_501;
      7:exp_504_reg <= exp_502;
      default:exp_504_reg <= exp_503;
    endcase
  end
  assign exp_504 = exp_504_reg;
  assign exp_503 = 0;
  assign exp_491 = exp_487 << exp_490;
  assign exp_487 = 1;
  assign exp_490 = exp_489 + exp_488;
  assign exp_489 = 0;
  assign exp_488 = exp_424[1:0];
  assign exp_496 = exp_492 << exp_495;
  assign exp_492 = 3;
  assign exp_495 = exp_494 + exp_493;
  assign exp_494 = 0;
  assign exp_493 = exp_424[1:1];
  assign exp_497 = 15;
  assign exp_498 = 0;
  assign exp_499 = 0;
  assign exp_500 = 0;
  assign exp_501 = 0;
  assign exp_502 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_218;
  assign exp_218 = exp_486;

  reg [31:0] exp_486_reg;
  always@(*) begin
    case (exp_356)
      0:exp_486_reg <= exp_473;
      1:exp_486_reg <= exp_477;
      2:exp_486_reg <= exp_479;
      3:exp_486_reg <= exp_480;
      4:exp_486_reg <= exp_481;
      5:exp_486_reg <= exp_482;
      6:exp_486_reg <= exp_483;
      7:exp_486_reg <= exp_484;
      default:exp_486_reg <= exp_485;
    endcase
  end
  assign exp_486 = exp_486_reg;
  assign exp_485 = 0;

  reg [31:0] exp_473_reg;
  always@(*) begin
    case (exp_427)
      0:exp_473_reg <= exp_459;
      1:exp_473_reg <= exp_467;
      2:exp_473_reg <= exp_469;
      3:exp_473_reg <= exp_471;
      default:exp_473_reg <= exp_472;
    endcase
  end
  assign exp_473 = exp_473_reg;
  assign exp_472 = 0;
  assign exp_459 = exp_458;
  assign exp_458 = exp_457 + exp_456;
  assign exp_457 = 0;
  assign exp_456 = exp_346[7:0];

      reg [31:0] exp_346_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_346_reg <= exp_289;
        end
      end
      assign exp_346 = exp_346_reg;
      assign exp_467 = exp_459 << exp_466;
  assign exp_466 = 8;
  assign exp_469 = exp_459 << exp_468;
  assign exp_468 = 16;
  assign exp_471 = exp_459 << exp_470;
  assign exp_470 = 24;

  reg [31:0] exp_477_reg;
  always@(*) begin
    case (exp_430)
      0:exp_477_reg <= exp_463;
      1:exp_477_reg <= exp_475;
      default:exp_477_reg <= exp_476;
    endcase
  end
  assign exp_477 = exp_477_reg;
  assign exp_430 = exp_429 + exp_428;
  assign exp_429 = 0;
  assign exp_428 = exp_424[1:1];
  assign exp_476 = 0;
  assign exp_463 = exp_462;
  assign exp_462 = exp_461 + exp_460;
  assign exp_461 = 0;
  assign exp_460 = exp_346[15:0];
  assign exp_475 = exp_463 << exp_474;
  assign exp_474 = 16;
  assign exp_479 = exp_478 + exp_465;
  assign exp_478 = 0;
  assign exp_465 = exp_464 + exp_346;
  assign exp_464 = 0;
  assign exp_480 = 0;
  assign exp_481 = 0;
  assign exp_482 = 0;
  assign exp_483 = 0;
  assign exp_484 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [1048575:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 16;
    exp_47_ram[32] = 193;
    exp_47_ram[33] = 128;
    exp_47_ram[34] = 0;
    exp_47_ram[35] = 5;
    exp_47_ram[36] = 0;
    exp_47_ram[37] = 167;
    exp_47_ram[38] = 7;
    exp_47_ram[39] = 7;
    exp_47_ram[40] = 0;
    exp_47_ram[41] = 21;
    exp_47_ram[42] = 229;
    exp_47_ram[43] = 159;
    exp_47_ram[44] = 0;
    exp_47_ram[45] = 133;
    exp_47_ram[46] = 95;
    exp_47_ram[47] = 64;
    exp_47_ram[48] = 31;
    exp_47_ram[49] = 108;
    exp_47_ram[50] = 87;
    exp_47_ram[51] = 100;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [1048575:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 1;
    exp_40_ram[32] = 1;
    exp_40_ram[33] = 0;
    exp_40_ram[34] = 0;
    exp_40_ram[35] = 7;
    exp_40_ram[36] = 5;
    exp_40_ram[37] = 135;
    exp_40_ram[38] = 71;
    exp_40_ram[39] = 20;
    exp_40_ram[40] = 128;
    exp_40_ram[41] = 5;
    exp_40_ram[42] = 160;
    exp_40_ram[43] = 240;
    exp_40_ram[44] = 5;
    exp_40_ram[45] = 133;
    exp_40_ram[46] = 240;
    exp_40_ram[47] = 5;
    exp_40_ram[48] = 240;
    exp_40_ram[49] = 101;
    exp_40_ram[50] = 32;
    exp_40_ram[51] = 108;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [1048575:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 55;
    exp_33_ram[32] = 19;
    exp_33_ram[33] = 239;
    exp_33_ram[34] = 111;
    exp_33_ram[35] = 147;
    exp_33_ram[36] = 19;
    exp_33_ram[37] = 51;
    exp_33_ram[38] = 3;
    exp_33_ram[39] = 99;
    exp_33_ram[40] = 103;
    exp_33_ram[41] = 19;
    exp_33_ram[42] = 35;
    exp_33_ram[43] = 111;
    exp_33_ram[44] = 183;
    exp_33_ram[45] = 147;
    exp_33_ram[46] = 111;
    exp_33_ram[47] = 19;
    exp_33_ram[48] = 111;
    exp_33_ram[49] = 72;
    exp_33_ram[50] = 111;
    exp_33_ram[51] = 114;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_172;

  reg [31:0] exp_172_reg;
  always@(*) begin
    case (exp_168)
      0:exp_172_reg <= exp_169;
      1:exp_172_reg <= exp_170;
      default:exp_172_reg <= exp_171;
    endcase
  end
  assign exp_172 = exp_172_reg;
  assign exp_168 = exp_139[2:2];
  assign exp_139 = exp_1;
  assign exp_171 = 0;
  assign exp_169 = exp_157[31:0];

      reg [63:0] exp_157_reg = 0;
      always@(posedge clk) begin
        if (exp_156) begin
          exp_157_reg <= exp_164;
        end
      end
      assign exp_157 = exp_157_reg;
    
  reg [63:0] exp_164_reg;
  always@(*) begin
    case (exp_159)
      0:exp_164_reg <= exp_161;
      1:exp_164_reg <= exp_162;
      default:exp_164_reg <= exp_163;
    endcase
  end
  assign exp_164 = exp_164_reg;
  assign exp_159 = exp_157 == exp_158;
  assign exp_158 = 18446744073709551616;
  assign exp_163 = 0;
  assign exp_161 = exp_157 + exp_160;
  assign exp_160 = 1;
  assign exp_162 = 0;
  assign exp_156 = 1;
  assign exp_170 = exp_157[63:32];
  assign exp_175 = exp_194;
  assign exp_194 = 0;
  assign exp_197 = exp_216;
  assign exp_216 = 0;
  assign exp_432 = exp_219[15:8];
  assign exp_433 = exp_219[23:16];
  assign exp_434 = exp_219[31:24];
  assign exp_446 = $signed(exp_445);
  assign exp_445 = exp_444 + exp_440;
  assign exp_444 = 0;

  reg [15:0] exp_440_reg;
  always@(*) begin
    case (exp_430)
      0:exp_440_reg <= exp_437;
      1:exp_440_reg <= exp_438;
      default:exp_440_reg <= exp_439;
    endcase
  end
  assign exp_440 = exp_440_reg;
  assign exp_439 = 0;
  assign exp_437 = exp_219[15:0];
  assign exp_438 = exp_219[31:16];
  assign exp_447 = 0;
  assign exp_448 = exp_436;
  assign exp_449 = exp_440;
  assign exp_450 = 0;
  assign exp_451 = 0;

  reg [31:0] exp_809_reg;
  always@(*) begin
    case (exp_599)
      0:exp_809_reg <= exp_805;
      1:exp_809_reg <= exp_807;
      default:exp_809_reg <= exp_808;
    endcase
  end
  assign exp_809 = exp_809_reg;
  assign exp_808 = 0;

  reg [31:0] exp_805_reg;
  always@(*) begin
    case (exp_576)
      0:exp_805_reg <= exp_800;
      1:exp_805_reg <= exp_801;
      default:exp_805_reg <= exp_804;
    endcase
  end
  assign exp_805 = exp_805_reg;
  assign exp_576 = exp_575 & exp_573;
  assign exp_575 = exp_568 == exp_574;
  assign exp_574 = 0;
  assign exp_804 = 0;
  assign exp_800 = exp_799[63:32];

  reg [63:0] exp_799_reg;
  always@(*) begin
    case (exp_796)
      0:exp_799_reg <= exp_795;
      1:exp_799_reg <= exp_797;
      default:exp_799_reg <= exp_798;
    endcase
  end
  assign exp_799 = exp_799_reg;

      reg [0:0] exp_796_reg = 0;
      always@(posedge clk) begin
        if (exp_781) begin
          exp_796_reg <= exp_779;
        end
      end
      assign exp_796 = exp_796_reg;
    
      reg [0:0] exp_779_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_779_reg <= exp_756;
        end
      end
      assign exp_779 = exp_779_reg;
    
      reg [0:0] exp_756_reg = 0;
      always@(posedge clk) begin
        if (exp_738) begin
          exp_756_reg <= exp_753;
        end
      end
      assign exp_756 = exp_756_reg;
      assign exp_753 = exp_751 ^ exp_752;
  assign exp_751 = exp_733 & exp_716;
  assign exp_733 = exp_732 + exp_731;
  assign exp_732 = 0;
  assign exp_731 = exp_729[31:31];

      reg [31:0] exp_729_reg = 0;
      always@(posedge clk) begin
        if (exp_728) begin
          exp_729_reg <= exp_347;
        end
      end
      assign exp_729 = exp_729_reg;
      assign exp_728 = exp_718 == exp_727;
  assign exp_727 = 0;
  assign exp_716 = exp_715 | exp_582;
  assign exp_715 = exp_576 | exp_579;
  assign exp_579 = exp_578 & exp_573;
  assign exp_578 = exp_568 == exp_577;
  assign exp_577 = 1;
  assign exp_582 = exp_581 & exp_573;
  assign exp_581 = exp_568 == exp_580;
  assign exp_580 = 2;
  assign exp_752 = exp_736 & exp_717;
  assign exp_736 = exp_735 + exp_734;
  assign exp_735 = 0;
  assign exp_734 = exp_730[31:31];

      reg [31:0] exp_730_reg = 0;
      always@(posedge clk) begin
        if (exp_728) begin
          exp_730_reg <= exp_348;
        end
      end
      assign exp_730 = exp_730_reg;
      assign exp_717 = exp_576 | exp_579;
  assign exp_738 = exp_718 == exp_737;
  assign exp_737 = 1;
  assign exp_758 = exp_718 == exp_757;
  assign exp_757 = 2;
  assign exp_781 = exp_718 == exp_780;
  assign exp_780 = 3;
  assign exp_798 = 0;

      reg [63:0] exp_795_reg = 0;
      always@(posedge clk) begin
        if (exp_781) begin
          exp_795_reg <= exp_794;
        end
      end
      assign exp_795 = exp_795_reg;
      assign exp_794 = exp_790 + exp_793;
  assign exp_790 = exp_786 + exp_789;
  assign exp_786 = exp_782 + exp_785;
  assign exp_782 = exp_775;

      reg [31:0] exp_775_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_775_reg <= exp_762;
        end
      end
      assign exp_775 = exp_775_reg;
      assign exp_762 = exp_760 * exp_761;
  assign exp_760 = exp_759;
  assign exp_759 = exp_754[15:0];

      reg [31:0] exp_754_reg = 0;
      always@(posedge clk) begin
        if (exp_738) begin
          exp_754_reg <= exp_744;
        end
      end
      assign exp_754 = exp_754_reg;
      assign exp_744 = exp_743 + exp_742;
  assign exp_743 = 0;

  reg [31:0] exp_742_reg;
  always@(*) begin
    case (exp_739)
      0:exp_742_reg <= exp_729;
      1:exp_742_reg <= exp_740;
      default:exp_742_reg <= exp_741;
    endcase
  end
  assign exp_742 = exp_742_reg;
  assign exp_739 = exp_733 & exp_716;
  assign exp_741 = 0;
  assign exp_740 = -exp_729;
  assign exp_761 = exp_755[15:0];

      reg [31:0] exp_755_reg = 0;
      always@(posedge clk) begin
        if (exp_738) begin
          exp_755_reg <= exp_750;
        end
      end
      assign exp_755 = exp_755_reg;
      assign exp_750 = exp_749 + exp_748;
  assign exp_749 = 0;

  reg [31:0] exp_748_reg;
  always@(*) begin
    case (exp_745)
      0:exp_748_reg <= exp_730;
      1:exp_748_reg <= exp_746;
      default:exp_748_reg <= exp_747;
    endcase
  end
  assign exp_748 = exp_748_reg;
  assign exp_745 = exp_736 & exp_717;
  assign exp_747 = 0;
  assign exp_746 = -exp_730;
  assign exp_785 = exp_783 << exp_784;
  assign exp_783 = exp_776;

      reg [31:0] exp_776_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_776_reg <= exp_766;
        end
      end
      assign exp_776 = exp_776_reg;
      assign exp_766 = exp_764 * exp_765;
  assign exp_764 = exp_763;
  assign exp_763 = exp_754[15:0];
  assign exp_765 = exp_755[31:16];
  assign exp_784 = 16;
  assign exp_789 = exp_787 << exp_788;
  assign exp_787 = exp_777;

      reg [31:0] exp_777_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_777_reg <= exp_770;
        end
      end
      assign exp_777 = exp_777_reg;
      assign exp_770 = exp_768 * exp_769;
  assign exp_768 = exp_767;
  assign exp_767 = exp_754[31:16];
  assign exp_769 = exp_755[15:0];
  assign exp_788 = 16;
  assign exp_793 = exp_791 << exp_792;
  assign exp_791 = exp_778;

      reg [31:0] exp_778_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_778_reg <= exp_774;
        end
      end
      assign exp_778 = exp_778_reg;
      assign exp_774 = exp_772 * exp_773;
  assign exp_772 = exp_771;
  assign exp_771 = exp_754[31:16];
  assign exp_773 = exp_755[31:16];
  assign exp_792 = 32;
  assign exp_797 = -exp_795;
  assign exp_801 = exp_799[31:0];

  reg [31:0] exp_807_reg;
  always@(*) begin
    case (exp_600)
      0:exp_807_reg <= exp_710;
      1:exp_807_reg <= exp_711;
      default:exp_807_reg <= exp_806;
    endcase
  end
  assign exp_807 = exp_807_reg;
  assign exp_600 = exp_568[1:1];
  assign exp_806 = 0;

      reg [31:0] exp_710_reg = 0;
      always@(posedge clk) begin
        if (exp_619) begin
          exp_710_reg <= exp_704;
        end
      end
      assign exp_710 = exp_710_reg;
    
  reg [31:0] exp_704_reg;
  always@(*) begin
    case (exp_700)
      0:exp_704_reg <= exp_691;
      1:exp_704_reg <= exp_702;
      default:exp_704_reg <= exp_703;
    endcase
  end
  assign exp_704 = exp_704_reg;
  assign exp_700 = exp_699 & exp_602;
  assign exp_699 = exp_648 == exp_698;

      reg [31:0] exp_648_reg = 0;
      always@(posedge clk) begin
        if (exp_633) begin
          exp_648_reg <= exp_645;
        end
      end
      assign exp_648 = exp_648_reg;
      assign exp_645 = exp_644 + exp_643;
  assign exp_644 = 0;

  reg [31:0] exp_643_reg;
  always@(*) begin
    case (exp_640)
      0:exp_643_reg <= exp_625;
      1:exp_643_reg <= exp_641;
      default:exp_643_reg <= exp_642;
    endcase
  end
  assign exp_643 = exp_643_reg;
  assign exp_640 = exp_631 & exp_602;
  assign exp_631 = exp_630 + exp_629;
  assign exp_630 = 0;
  assign exp_629 = exp_625[31:31];

      reg [31:0] exp_625_reg = 0;
      always@(posedge clk) begin
        if (exp_623) begin
          exp_625_reg <= exp_348;
        end
      end
      assign exp_625 = exp_625_reg;
      assign exp_623 = exp_605 == exp_622;
  assign exp_622 = 0;
  assign exp_602 = ~exp_601;
  assign exp_601 = exp_568[0:0];
  assign exp_642 = 0;
  assign exp_641 = -exp_625;
  assign exp_633 = exp_605 == exp_632;
  assign exp_632 = 1;
  assign exp_698 = 0;
  assign exp_703 = 0;
  assign exp_691 = exp_690 + exp_689;
  assign exp_690 = 0;

  reg [31:0] exp_689_reg;
  always@(*) begin
    case (exp_686)
      0:exp_689_reg <= exp_684;
      1:exp_689_reg <= exp_687;
      default:exp_689_reg <= exp_688;
    endcase
  end
  assign exp_689 = exp_689_reg;
  assign exp_686 = exp_650 & exp_602;

      reg [0:0] exp_650_reg = 0;
      always@(posedge clk) begin
        if (exp_633) begin
          exp_650_reg <= exp_646;
        end
      end
      assign exp_650 = exp_650_reg;
      assign exp_646 = exp_628 ^ exp_631;
  assign exp_628 = exp_627 + exp_626;
  assign exp_627 = 0;
  assign exp_626 = exp_624[31:31];

      reg [31:0] exp_624_reg = 0;
      always@(posedge clk) begin
        if (exp_623) begin
          exp_624_reg <= exp_347;
        end
      end
      assign exp_624 = exp_624_reg;
      assign exp_688 = 0;

      reg [31:0] exp_684_reg = 0;
      always@(posedge clk) begin
        if (exp_617) begin
          exp_684_reg <= exp_654;
        end
      end
      assign exp_684 = exp_684_reg;
    
      reg [31:0] exp_654_reg = 0;
      always@(posedge clk) begin
        if (exp_653) begin
          exp_654_reg <= exp_681;
        end
      end
      assign exp_654 = exp_654_reg;
    
  reg [31:0] exp_681_reg;
  always@(*) begin
    case (exp_615)
      0:exp_681_reg <= exp_673;
      1:exp_681_reg <= exp_679;
      default:exp_681_reg <= exp_680;
    endcase
  end
  assign exp_681 = exp_681_reg;
  assign exp_615 = exp_605 == exp_614;
  assign exp_614 = 2;
  assign exp_680 = 0;

  reg [31:0] exp_673_reg;
  always@(*) begin
    case (exp_663)
      0:exp_673_reg <= exp_667;
      1:exp_673_reg <= exp_671;
      default:exp_673_reg <= exp_672;
    endcase
  end
  assign exp_673 = exp_673_reg;
  assign exp_663 = ~exp_662;
  assign exp_662 = exp_661[32:32];
  assign exp_661 = exp_660 - exp_648;
  assign exp_660 = exp_659;
  assign exp_659 = {exp_657, exp_658};  assign exp_657 = exp_652[31:0];

      reg [31:0] exp_652_reg = 0;
      always@(posedge clk) begin
        if (exp_651) begin
          exp_652_reg <= exp_678;
        end
      end
      assign exp_652 = exp_652_reg;
    
  reg [32:0] exp_678_reg;
  always@(*) begin
    case (exp_615)
      0:exp_678_reg <= exp_665;
      1:exp_678_reg <= exp_676;
      default:exp_678_reg <= exp_677;
    endcase
  end
  assign exp_678 = exp_678_reg;
  assign exp_677 = 0;

  reg [32:0] exp_665_reg;
  always@(*) begin
    case (exp_663)
      0:exp_665_reg <= exp_659;
      1:exp_665_reg <= exp_661;
      default:exp_665_reg <= exp_664;
    endcase
  end
  assign exp_665 = exp_665_reg;
  assign exp_664 = 0;
  assign exp_676 = 0;
  assign exp_651 = 1;
  assign exp_658 = exp_656[31:31];

      reg [31:0] exp_656_reg = 0;
      always@(posedge clk) begin
        if (exp_655) begin
          exp_656_reg <= exp_683;
        end
      end
      assign exp_656 = exp_656_reg;
    
  reg [31:0] exp_683_reg;
  always@(*) begin
    case (exp_615)
      0:exp_683_reg <= exp_675;
      1:exp_683_reg <= exp_647;
      default:exp_683_reg <= exp_682;
    endcase
  end
  assign exp_683 = exp_683_reg;
  assign exp_682 = 0;
  assign exp_675 = exp_656 << exp_674;
  assign exp_674 = 1;

      reg [31:0] exp_647_reg = 0;
      always@(posedge clk) begin
        if (exp_633) begin
          exp_647_reg <= exp_639;
        end
      end
      assign exp_647 = exp_647_reg;
      assign exp_639 = exp_638 + exp_637;
  assign exp_638 = 0;

  reg [31:0] exp_637_reg;
  always@(*) begin
    case (exp_634)
      0:exp_637_reg <= exp_624;
      1:exp_637_reg <= exp_635;
      default:exp_637_reg <= exp_636;
    endcase
  end
  assign exp_637 = exp_637_reg;
  assign exp_634 = exp_628 & exp_602;
  assign exp_636 = 0;
  assign exp_635 = -exp_624;
  assign exp_655 = 1;
  assign exp_672 = 0;
  assign exp_667 = exp_654 << exp_666;
  assign exp_666 = 1;
  assign exp_671 = exp_669 | exp_670;
  assign exp_669 = exp_654 << exp_668;
  assign exp_668 = 1;
  assign exp_670 = 1;
  assign exp_679 = 0;
  assign exp_653 = 1;
  assign exp_617 = exp_605 == exp_616;
  assign exp_616 = 35;
  assign exp_687 = -exp_684;
  assign exp_702 = $signed(exp_701);
  assign exp_701 = -1;
  assign exp_619 = exp_605 == exp_618;
  assign exp_618 = 36;

      reg [31:0] exp_711_reg = 0;
      always@(posedge clk) begin
        if (exp_619) begin
          exp_711_reg <= exp_709;
        end
      end
      assign exp_711 = exp_711_reg;
    
  reg [31:0] exp_709_reg;
  always@(*) begin
    case (exp_707)
      0:exp_709_reg <= exp_697;
      1:exp_709_reg <= exp_624;
      default:exp_709_reg <= exp_708;
    endcase
  end
  assign exp_709 = exp_709_reg;
  assign exp_707 = exp_706 & exp_602;
  assign exp_706 = exp_648 == exp_705;
  assign exp_705 = 0;
  assign exp_708 = 0;
  assign exp_697 = exp_696 + exp_695;
  assign exp_696 = 0;

  reg [31:0] exp_695_reg;
  always@(*) begin
    case (exp_692)
      0:exp_695_reg <= exp_685;
      1:exp_695_reg <= exp_693;
      default:exp_695_reg <= exp_694;
    endcase
  end
  assign exp_695 = exp_695_reg;
  assign exp_692 = exp_649 & exp_602;

      reg [0:0] exp_649_reg = 0;
      always@(posedge clk) begin
        if (exp_633) begin
          exp_649_reg <= exp_628;
        end
      end
      assign exp_649 = exp_649_reg;
      assign exp_694 = 0;

      reg [31:0] exp_685_reg = 0;
      always@(posedge clk) begin
        if (exp_617) begin
          exp_685_reg <= exp_652;
        end
      end
      assign exp_685 = exp_685_reg;
      assign exp_693 = -exp_685;
  assign exp_281 = $signed(exp_280);
  assign exp_280 = 0;
  assign exp_510 = exp_345 != exp_346;
  assign exp_523 = 0;
  assign exp_524 = 0;
  assign exp_511 = $signed(exp_345) < $signed(exp_346);
  assign exp_512 = $signed(exp_345) >= $signed(exp_346);
  assign exp_517 = exp_514 < exp_516;
  assign exp_514 = exp_513 + exp_345;
  assign exp_513 = 0;
  assign exp_516 = exp_515 + exp_346;
  assign exp_515 = 0;
  assign exp_522 = exp_519 >= exp_521;
  assign exp_519 = exp_518 + exp_345;
  assign exp_518 = 0;
  assign exp_521 = exp_520 + exp_346;
  assign exp_520 = 0;
  assign exp_836 = 0;
  assign exp_835 = exp_235 + exp_834;
  assign exp_834 = 4;

  reg [32:0] exp_567_reg;
  always@(*) begin
    case (exp_368)
      0:exp_567_reg <= exp_557;
      1:exp_567_reg <= exp_565;
      default:exp_567_reg <= exp_566;
    endcase
  end
  assign exp_567 = exp_567_reg;
  assign exp_566 = 0;
  assign exp_557 = exp_556 + exp_354;

  reg [31:0] exp_556_reg;
  always@(*) begin
    case (exp_366)
      0:exp_556_reg <= exp_542;
      1:exp_556_reg <= exp_554;
      default:exp_556_reg <= exp_555;
    endcase
  end
  assign exp_556 = exp_556_reg;
  assign exp_555 = 0;
  assign exp_542 = $signed(exp_541);
  assign exp_541 = exp_540 + exp_539;
  assign exp_540 = 0;
  assign exp_539 = {exp_538, exp_535};  assign exp_538 = {exp_537, exp_534};  assign exp_537 = {exp_536, exp_533};  assign exp_536 = {exp_531, exp_532};  assign exp_531 = exp_353[31:31];
  assign exp_532 = exp_353[7:7];
  assign exp_533 = exp_353[30:25];
  assign exp_534 = exp_353[11:8];
  assign exp_535 = 0;
  assign exp_554 = $signed(exp_553);
  assign exp_553 = exp_552 + exp_551;
  assign exp_552 = 0;
  assign exp_551 = {exp_550, exp_547};  assign exp_550 = {exp_549, exp_546};  assign exp_549 = {exp_548, exp_545};  assign exp_548 = {exp_543, exp_544};  assign exp_543 = exp_353[31:31];
  assign exp_544 = exp_353[19:12];
  assign exp_545 = exp_353[20:20];
  assign exp_546 = exp_353[30:21];
  assign exp_547 = 0;

      reg [31:0] exp_354_reg = 0;
      always@(posedge clk) begin
        if (exp_344) begin
          exp_354_reg <= exp_237;
        end
      end
      assign exp_354 = exp_354_reg;
      assign exp_565 = exp_564 & exp_563;
  assign exp_564 = $signed(exp_562);
  assign exp_562 = exp_345 + exp_561;
  assign exp_561 = $signed(exp_560);
  assign exp_560 = exp_559 + exp_558;
  assign exp_559 = 0;
  assign exp_558 = exp_353[31:20];
  assign exp_563 = 4294967294;
  assign exp_234 = exp_227 & exp_225;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_236;
  assign exp_369 = 3;
  assign exp_178 = exp_6;
  assign exp_174 = exp_2;
  assign exp_215 = exp_199 & exp_200;
  assign exp_199 = exp_207;
  assign exp_207 = exp_5 & exp_206;
  assign exp_200 = exp_6;
  assign exp_196 = exp_2;
  assign stdout_valid_out = exp_193;
  assign stdout_out = exp_174;
  assign spare_valid_out = exp_215;
  assign spare_out = exp_196;

endmodule