
module hello_world(clk, stdin_valid_in, stdin_in, stdout_ready_in, stdin_ready_out, stdout_valid_out, stdout_out);
  input [0:0] stdin_valid_in;
  input [31:0] stdin_in;
  input [0:0] stdout_ready_in;
  input [0:0] clk;
  output [0:0] stdin_ready_out;
  output [0:0] stdout_valid_out;
  output [31:0] stdout_out;
  wire [0:0] exp_223;
  wire [0:0] exp_206;
  wire [0:0] exp_214;
  wire [0:0] exp_5;
  wire [0:0] exp_228;
  wire [0:0] exp_575;
  wire [0:0] exp_512;
  wire [0:0] exp_377;
  wire [6:0] exp_362;
  wire [31:0] exp_360;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [10:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_242;
  wire [32:0] exp_845;
  wire [0:0] exp_841;
  wire [0:0] exp_537;
  wire [0:0] exp_515;
  wire [0:0] exp_373;
  wire [6:0] exp_372;
  wire [0:0] exp_375;
  wire [6:0] exp_374;
  wire [0:0] exp_536;
  wire [0:0] exp_381;
  wire [6:0] exp_380;
  wire [0:0] exp_535;
  wire [0:0] exp_534;
  wire [0:0] exp_533;
  wire [2:0] exp_363;
  wire [0:0] exp_532;
  wire [0:0] exp_516;
  wire [31:0] exp_352;
  wire [31:0] exp_290;
  wire [0:0] exp_286;
  wire [4:0] exp_266;
  wire [0:0] exp_285;
  wire [0:0] exp_289;
  wire [31:0] exp_282;
  wire [0:0] exp_263;
  wire [0:0] exp_836;
  wire [0:0] exp_835;
  wire [0:0] exp_834;
  wire [0:0] exp_833;
  wire [4:0] exp_245;
  wire [4:0] exp_828;
  wire [0:0] exp_827;
  wire [0:0] exp_419;
  wire [0:0] exp_418;
  wire [0:0] exp_417;
  wire [0:0] exp_416;
  wire [0:0] exp_415;
  wire [0:0] exp_414;
  wire [0:0] exp_365;
  wire [4:0] exp_364;
  wire [0:0] exp_367;
  wire [5:0] exp_366;
  wire [0:0] exp_369;
  wire [5:0] exp_368;
  wire [0:0] exp_371;
  wire [4:0] exp_370;
  wire [0:0] exp_822;
  wire [0:0] exp_821;
  wire [0:0] exp_607;
  wire [0:0] exp_581;
  wire [0:0] exp_579;
  wire [6:0] exp_577;
  wire [5:0] exp_578;
  wire [0:0] exp_580;
  wire [0:0] exp_606;
  wire [2:0] exp_576;
  wire [0:0] exp_820;
  wire [0:0] exp_818;
  wire [0:0] exp_811;
  wire [2:0] exp_726;
  wire [2:0] exp_733;
  wire [0:0] exp_728;
  wire [2:0] exp_727;
  wire [0:0] exp_732;
  wire [2:0] exp_730;
  wire [0:0] exp_729;
  wire [0:0] exp_731;
  wire [0:0] exp_722;
  wire [0:0] exp_721;
  wire [0:0] exp_720;
  wire [2:0] exp_810;
  wire [0:0] exp_819;
  wire [0:0] exp_629;
  wire [5:0] exp_613;
  wire [5:0] exp_620;
  wire [0:0] exp_615;
  wire [5:0] exp_614;
  wire [0:0] exp_619;
  wire [5:0] exp_617;
  wire [0:0] exp_616;
  wire [0:0] exp_618;
  wire [5:0] exp_628;
  wire [0:0] exp_240;
  wire [0:0] exp_239;
  wire [0:0] exp_237;
  wire [0:0] exp_236;
  wire [0:0] exp_234;
  wire [0:0] exp_235;
  wire [0:0] exp_233;
  wire [0:0] exp_846;
  wire [0:0] exp_232;
  wire [0:0] exp_231;
  wire [0:0] exp_850;
  wire [0:0] exp_849;
  wire [0:0] exp_848;
  wire [0:0] exp_847;
  wire [0:0] exp_227;
  wire [0:0] exp_218;
  wire [0:0] exp_213;
  wire [0:0] exp_210;
  wire [31:0] exp_1;
  wire [31:0] exp_224;
  wire [31:0] exp_431;
  wire [31:0] exp_430;
  wire [31:0] exp_429;
  wire [31:0] exp_428;
  wire [11:0] exp_427;
  wire [11:0] exp_426;
  wire [11:0] exp_425;
  wire [0:0] exp_379;
  wire [5:0] exp_378;
  wire [0:0] exp_424;
  wire [11:0] exp_420;
  wire [11:0] exp_423;
  wire [6:0] exp_421;
  wire [4:0] exp_422;
  wire [31:0] exp_209;
  wire [0:0] exp_212;
  wire [31:0] exp_211;
  wire [0:0] exp_217;
  wire [0:0] exp_196;
  wire [0:0] exp_191;
  wire [0:0] exp_188;
  wire [31:0] exp_187;
  wire [0:0] exp_190;
  wire [31:0] exp_189;
  wire [0:0] exp_195;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [31:0] exp_146;
  wire [0:0] exp_149;
  wire [31:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [12:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_229;
  wire [0:0] exp_514;
  wire [0:0] exp_513;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_176;
  wire [0:0] exp_183;
  wire [0:0] exp_198;
  wire [0:0] exp_205;
  wire [0:0] exp_221;
  wire [0:0] exp_824;
  wire [0:0] exp_823;
  wire [0:0] exp_238;
  wire [0:0] exp_281;
  wire [31:0] exp_253;
  wire [0:0] exp_252;
  wire [1:0] exp_261;
  wire [4:0] exp_248;
  wire [0:0] exp_251;
  wire [0:0] exp_830;
  wire [0:0] exp_829;
  wire [4:0] exp_247;
  wire [31:0] exp_249;
  wire [31:0] exp_826;
  wire [0:0] exp_825;
  wire [31:0] exp_462;
  wire [0:0] exp_461;
  wire [31:0] exp_413;
  wire [2:0] exp_356;
  wire [2:0] exp_347;
  wire [0:0] exp_344;
  wire [0:0] exp_278;
  wire [6:0] exp_268;
  wire [6:0] exp_277;
  wire [0:0] exp_280;
  wire [6:0] exp_279;
  wire [0:0] exp_346;
  wire [2:0] exp_334;
  wire [0:0] exp_276;
  wire [4:0] exp_275;
  wire [0:0] exp_333;
  wire [2:0] exp_321;
  wire [0:0] exp_274;
  wire [5:0] exp_273;
  wire [0:0] exp_320;
  wire [2:0] exp_270;
  wire [0:0] exp_319;
  wire [0:0] exp_332;
  wire [0:0] exp_345;
  wire [0:0] exp_351;
  wire [0:0] exp_412;
  wire [31:0] exp_392;
  wire [0:0] exp_358;
  wire [0:0] exp_350;
  wire [0:0] exp_336;
  wire [0:0] exp_323;
  wire [0:0] exp_309;
  wire [0:0] exp_307;
  wire [0:0] exp_308;
  wire [0:0] exp_272;
  wire [4:0] exp_271;
  wire [0:0] exp_322;
  wire [0:0] exp_335;
  wire [0:0] exp_349;
  wire [0:0] exp_348;
  wire [0:0] exp_391;
  wire [31:0] exp_389;
  wire [31:0] exp_354;
  wire [31:0] exp_340;
  wire [0:0] exp_337;
  wire [0:0] exp_339;
  wire [31:0] exp_329;
  wire [0:0] exp_328;
  wire [31:0] exp_315;
  wire [0:0] exp_314;
  wire [31:0] exp_313;
  wire [31:0] exp_311;
  wire [19:0] exp_310;
  wire [3:0] exp_312;
  wire [31:0] exp_327;
  wire [31:0] exp_325;
  wire [19:0] exp_324;
  wire [3:0] exp_326;
  wire [31:0] exp_338;
  wire [31:0] exp_355;
  wire [31:0] exp_343;
  wire [0:0] exp_341;
  wire [0:0] exp_342;
  wire [31:0] exp_331;
  wire [0:0] exp_330;
  wire [31:0] exp_318;
  wire [0:0] exp_317;
  wire [31:0] exp_302;
  wire [0:0] exp_301;
  wire [31:0] exp_296;
  wire [0:0] exp_292;
  wire [4:0] exp_267;
  wire [0:0] exp_291;
  wire [0:0] exp_295;
  wire [31:0] exp_284;
  wire [0:0] exp_264;
  wire [0:0] exp_840;
  wire [0:0] exp_839;
  wire [0:0] exp_838;
  wire [0:0] exp_837;
  wire [4:0] exp_246;
  wire [0:0] exp_283;
  wire [31:0] exp_260;
  wire [0:0] exp_259;
  wire [1:0] exp_262;
  wire [4:0] exp_255;
  wire [0:0] exp_258;
  wire [0:0] exp_832;
  wire [0:0] exp_831;
  wire [4:0] exp_254;
  wire [31:0] exp_256;
  wire [31:0] exp_265;
  wire [31:0] exp_294;
  wire [0:0] exp_293;
  wire [31:0] exp_300;
  wire [31:0] exp_297;
  wire [31:0] exp_299;
  wire [11:0] exp_298;
  wire [31:0] exp_316;
  wire [31:0] exp_244;
  wire [0:0] exp_243;
  wire [31:0] exp_390;
  wire [31:0] exp_394;
  wire [31:0] exp_393;
  wire [5:0] exp_388;
  wire [5:0] exp_387;
  wire [5:0] exp_386;
  wire [4:0] exp_357;
  wire [4:0] exp_306;
  wire [0:0] exp_305;
  wire [4:0] exp_304;
  wire [4:0] exp_269;
  wire [31:0] exp_410;
  wire [1:0] exp_396;
  wire [0:0] exp_395;
  wire [31:0] exp_411;
  wire [1:0] exp_402;
  wire [0:0] exp_401;
  wire [31:0] exp_398;
  wire [31:0] exp_397;
  wire [31:0] exp_400;
  wire [31:0] exp_399;
  wire [31:0] exp_403;
  wire [31:0] exp_407;
  wire [32:0] exp_406;
  wire [32:0] exp_404;
  wire [0:0] exp_385;
  wire [0:0] exp_359;
  wire [0:0] exp_303;
  wire [0:0] exp_384;
  wire [0:0] exp_383;
  wire [0:0] exp_382;
  wire [32:0] exp_405;
  wire [31:0] exp_408;
  wire [31:0] exp_409;
  wire [31:0] exp_460;
  wire [0:0] exp_459;
  wire [31:0] exp_450;
  wire [7:0] exp_449;
  wire [7:0] exp_448;
  wire [7:0] exp_443;
  wire [1:0] exp_434;
  wire [1:0] exp_433;
  wire [1:0] exp_432;
  wire [0:0] exp_442;
  wire [7:0] exp_438;
  wire [31:0] exp_226;
  wire [31:0] exp_216;
  wire [0:0] exp_215;
  wire [31:0] exp_194;
  wire [0:0] exp_193;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [10:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_230;
  wire [3:0] exp_511;
  wire [0:0] exp_510;
  wire [3:0] exp_498;
  wire [3:0] exp_494;
  wire [1:0] exp_497;
  wire [1:0] exp_496;
  wire [1:0] exp_495;
  wire [3:0] exp_503;
  wire [3:0] exp_499;
  wire [0:0] exp_502;
  wire [0:0] exp_501;
  wire [0:0] exp_500;
  wire [3:0] exp_504;
  wire [3:0] exp_505;
  wire [3:0] exp_506;
  wire [3:0] exp_507;
  wire [3:0] exp_508;
  wire [3:0] exp_509;
  wire [10:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_225;
  wire [31:0] exp_493;
  wire [0:0] exp_492;
  wire [31:0] exp_480;
  wire [0:0] exp_479;
  wire [31:0] exp_466;
  wire [7:0] exp_465;
  wire [7:0] exp_464;
  wire [7:0] exp_463;
  wire [31:0] exp_353;
  wire [31:0] exp_474;
  wire [3:0] exp_473;
  wire [31:0] exp_476;
  wire [4:0] exp_475;
  wire [31:0] exp_478;
  wire [4:0] exp_477;
  wire [31:0] exp_484;
  wire [0:0] exp_437;
  wire [0:0] exp_436;
  wire [0:0] exp_435;
  wire [0:0] exp_483;
  wire [31:0] exp_470;
  wire [15:0] exp_469;
  wire [15:0] exp_468;
  wire [15:0] exp_467;
  wire [31:0] exp_482;
  wire [4:0] exp_481;
  wire [31:0] exp_486;
  wire [31:0] exp_485;
  wire [31:0] exp_472;
  wire [31:0] exp_471;
  wire [31:0] exp_487;
  wire [31:0] exp_488;
  wire [31:0] exp_489;
  wire [31:0] exp_490;
  wire [31:0] exp_491;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [10:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [10:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [10:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [10:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [10:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [10:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [10:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [10:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [10:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [10:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [10:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [10:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_179;
  wire [0:0] exp_177;
  wire [31:0] exp_139;
  wire [0:0] exp_178;
  wire [31:0] exp_157;
  wire [31:0] exp_164;
  wire [0:0] exp_159;
  wire [31:0] exp_158;
  wire [0:0] exp_163;
  wire [31:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [31:0] exp_167;
  wire [31:0] exp_174;
  wire [0:0] exp_169;
  wire [31:0] exp_168;
  wire [0:0] exp_173;
  wire [31:0] exp_171;
  wire [0:0] exp_170;
  wire [0:0] exp_172;
  wire [0:0] exp_166;
  wire [0:0] exp_165;
  wire [31:0] exp_182;
  wire [31:0] exp_201;
  wire [31:0] exp_204;
  wire [31:0] exp_219;
  wire [7:0] exp_439;
  wire [7:0] exp_440;
  wire [7:0] exp_441;
  wire [31:0] exp_453;
  wire [15:0] exp_452;
  wire [15:0] exp_451;
  wire [15:0] exp_447;
  wire [0:0] exp_446;
  wire [15:0] exp_444;
  wire [15:0] exp_445;
  wire [31:0] exp_454;
  wire [31:0] exp_455;
  wire [31:0] exp_456;
  wire [31:0] exp_457;
  wire [31:0] exp_458;
  wire [31:0] exp_817;
  wire [0:0] exp_816;
  wire [31:0] exp_813;
  wire [0:0] exp_584;
  wire [0:0] exp_583;
  wire [0:0] exp_582;
  wire [0:0] exp_812;
  wire [31:0] exp_808;
  wire [63:0] exp_807;
  wire [0:0] exp_804;
  wire [0:0] exp_787;
  wire [0:0] exp_764;
  wire [0:0] exp_761;
  wire [0:0] exp_759;
  wire [0:0] exp_741;
  wire [0:0] exp_740;
  wire [0:0] exp_739;
  wire [31:0] exp_737;
  wire [0:0] exp_736;
  wire [0:0] exp_735;
  wire [0:0] exp_724;
  wire [0:0] exp_723;
  wire [0:0] exp_587;
  wire [0:0] exp_586;
  wire [0:0] exp_585;
  wire [0:0] exp_590;
  wire [0:0] exp_589;
  wire [1:0] exp_588;
  wire [0:0] exp_760;
  wire [0:0] exp_744;
  wire [0:0] exp_743;
  wire [0:0] exp_742;
  wire [31:0] exp_738;
  wire [0:0] exp_725;
  wire [0:0] exp_746;
  wire [0:0] exp_745;
  wire [0:0] exp_766;
  wire [1:0] exp_765;
  wire [0:0] exp_789;
  wire [1:0] exp_788;
  wire [0:0] exp_806;
  wire [63:0] exp_803;
  wire [63:0] exp_802;
  wire [63:0] exp_798;
  wire [63:0] exp_794;
  wire [63:0] exp_790;
  wire [31:0] exp_783;
  wire [31:0] exp_770;
  wire [31:0] exp_768;
  wire [15:0] exp_767;
  wire [31:0] exp_762;
  wire [31:0] exp_752;
  wire [31:0] exp_751;
  wire [31:0] exp_750;
  wire [0:0] exp_747;
  wire [0:0] exp_749;
  wire [31:0] exp_748;
  wire [15:0] exp_769;
  wire [31:0] exp_763;
  wire [31:0] exp_758;
  wire [31:0] exp_757;
  wire [31:0] exp_756;
  wire [0:0] exp_753;
  wire [0:0] exp_755;
  wire [31:0] exp_754;
  wire [63:0] exp_793;
  wire [63:0] exp_791;
  wire [31:0] exp_784;
  wire [31:0] exp_774;
  wire [31:0] exp_772;
  wire [15:0] exp_771;
  wire [15:0] exp_773;
  wire [4:0] exp_792;
  wire [63:0] exp_797;
  wire [63:0] exp_795;
  wire [31:0] exp_785;
  wire [31:0] exp_778;
  wire [31:0] exp_776;
  wire [15:0] exp_775;
  wire [15:0] exp_777;
  wire [4:0] exp_796;
  wire [63:0] exp_801;
  wire [63:0] exp_799;
  wire [31:0] exp_786;
  wire [31:0] exp_782;
  wire [31:0] exp_780;
  wire [15:0] exp_779;
  wire [15:0] exp_781;
  wire [5:0] exp_800;
  wire [63:0] exp_805;
  wire [31:0] exp_809;
  wire [31:0] exp_815;
  wire [0:0] exp_608;
  wire [0:0] exp_814;
  wire [31:0] exp_718;
  wire [31:0] exp_712;
  wire [0:0] exp_708;
  wire [0:0] exp_707;
  wire [31:0] exp_656;
  wire [31:0] exp_653;
  wire [31:0] exp_652;
  wire [31:0] exp_651;
  wire [0:0] exp_648;
  wire [0:0] exp_639;
  wire [0:0] exp_638;
  wire [0:0] exp_637;
  wire [31:0] exp_633;
  wire [0:0] exp_631;
  wire [0:0] exp_630;
  wire [0:0] exp_610;
  wire [0:0] exp_609;
  wire [0:0] exp_650;
  wire [31:0] exp_649;
  wire [0:0] exp_641;
  wire [0:0] exp_640;
  wire [0:0] exp_706;
  wire [0:0] exp_711;
  wire [31:0] exp_699;
  wire [31:0] exp_698;
  wire [31:0] exp_697;
  wire [0:0] exp_694;
  wire [0:0] exp_658;
  wire [0:0] exp_654;
  wire [0:0] exp_636;
  wire [0:0] exp_635;
  wire [0:0] exp_634;
  wire [31:0] exp_632;
  wire [0:0] exp_696;
  wire [31:0] exp_692;
  wire [31:0] exp_662;
  wire [31:0] exp_689;
  wire [0:0] exp_623;
  wire [1:0] exp_622;
  wire [0:0] exp_688;
  wire [31:0] exp_681;
  wire [0:0] exp_671;
  wire [0:0] exp_670;
  wire [32:0] exp_669;
  wire [32:0] exp_668;
  wire [32:0] exp_667;
  wire [31:0] exp_665;
  wire [31:0] exp_660;
  wire [32:0] exp_686;
  wire [0:0] exp_685;
  wire [32:0] exp_673;
  wire [0:0] exp_672;
  wire [0:0] exp_684;
  wire [0:0] exp_659;
  wire [0:0] exp_666;
  wire [31:0] exp_664;
  wire [31:0] exp_691;
  wire [0:0] exp_690;
  wire [31:0] exp_683;
  wire [0:0] exp_682;
  wire [31:0] exp_655;
  wire [31:0] exp_647;
  wire [31:0] exp_646;
  wire [31:0] exp_645;
  wire [0:0] exp_642;
  wire [0:0] exp_644;
  wire [31:0] exp_643;
  wire [0:0] exp_663;
  wire [0:0] exp_680;
  wire [31:0] exp_675;
  wire [0:0] exp_674;
  wire [31:0] exp_679;
  wire [31:0] exp_677;
  wire [0:0] exp_676;
  wire [0:0] exp_678;
  wire [0:0] exp_687;
  wire [0:0] exp_661;
  wire [0:0] exp_625;
  wire [5:0] exp_624;
  wire [31:0] exp_695;
  wire [31:0] exp_710;
  wire [0:0] exp_709;
  wire [0:0] exp_627;
  wire [5:0] exp_626;
  wire [31:0] exp_719;
  wire [31:0] exp_717;
  wire [0:0] exp_715;
  wire [0:0] exp_714;
  wire [0:0] exp_713;
  wire [0:0] exp_716;
  wire [31:0] exp_705;
  wire [31:0] exp_704;
  wire [31:0] exp_703;
  wire [0:0] exp_700;
  wire [0:0] exp_657;
  wire [0:0] exp_702;
  wire [31:0] exp_693;
  wire [31:0] exp_701;
  wire [31:0] exp_288;
  wire [0:0] exp_287;
  wire [0:0] exp_517;
  wire [0:0] exp_530;
  wire [0:0] exp_531;
  wire [0:0] exp_518;
  wire [0:0] exp_519;
  wire [0:0] exp_524;
  wire [31:0] exp_521;
  wire [31:0] exp_520;
  wire [31:0] exp_523;
  wire [31:0] exp_522;
  wire [0:0] exp_529;
  wire [31:0] exp_526;
  wire [31:0] exp_525;
  wire [31:0] exp_528;
  wire [31:0] exp_527;
  wire [0:0] exp_844;
  wire [31:0] exp_843;
  wire [2:0] exp_842;
  wire [32:0] exp_574;
  wire [0:0] exp_573;
  wire [31:0] exp_564;
  wire [31:0] exp_563;
  wire [0:0] exp_562;
  wire [31:0] exp_549;
  wire [12:0] exp_548;
  wire [12:0] exp_547;
  wire [12:0] exp_546;
  wire [11:0] exp_545;
  wire [7:0] exp_544;
  wire [1:0] exp_543;
  wire [0:0] exp_538;
  wire [0:0] exp_539;
  wire [5:0] exp_540;
  wire [3:0] exp_541;
  wire [0:0] exp_542;
  wire [31:0] exp_561;
  wire [20:0] exp_560;
  wire [20:0] exp_559;
  wire [20:0] exp_558;
  wire [19:0] exp_557;
  wire [9:0] exp_556;
  wire [8:0] exp_555;
  wire [0:0] exp_550;
  wire [7:0] exp_551;
  wire [0:0] exp_552;
  wire [9:0] exp_553;
  wire [0:0] exp_554;
  wire [31:0] exp_361;
  wire [32:0] exp_572;
  wire [32:0] exp_571;
  wire [31:0] exp_569;
  wire [31:0] exp_568;
  wire [11:0] exp_567;
  wire [11:0] exp_566;
  wire [11:0] exp_565;
  wire [32:0] exp_570;
  wire [0:0] exp_241;
  wire [0:0] exp_80;
  wire [10:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_376;
  wire [0:0] exp_222;
  wire [0:0] exp_207;
  wire [0:0] exp_200;
  wire [0:0] exp_184;
  wire [0:0] exp_192;
  wire [0:0] exp_185;
  wire [31:0] exp_181;

  assign exp_223 = exp_206 & exp_222;
  assign exp_206 = exp_214;
  assign exp_214 = exp_5 & exp_213;
  assign exp_5 = exp_228;
  assign exp_228 = exp_575;
  assign exp_575 = exp_512 & exp_240;
  assign exp_512 = exp_377 | exp_379;
  assign exp_377 = exp_362 == exp_376;
  assign exp_362 = exp_360[6:0];

      reg [31:0] exp_360_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_360_reg <= exp_96;
        end
      end
      assign exp_360 = exp_360_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_242;

      reg [31:0] exp_242_reg = 0;
      always@(posedge clk) begin
        if (exp_241) begin
          exp_242_reg <= exp_845;
        end
      end
      assign exp_242 = exp_242_reg;
    
  reg [32:0] exp_845_reg;
  always@(*) begin
    case (exp_841)
      0:exp_845_reg <= exp_843;
      1:exp_845_reg <= exp_574;
      default:exp_845_reg <= exp_844;
    endcase
  end
  assign exp_845 = exp_845_reg;
  assign exp_841 = exp_537 & exp_240;
  assign exp_537 = exp_515 | exp_536;
  assign exp_515 = exp_373 | exp_375;
  assign exp_373 = exp_362 == exp_372;
  assign exp_372 = 111;
  assign exp_375 = exp_362 == exp_374;
  assign exp_374 = 103;

  reg [0:0] exp_536_reg;
  always@(*) begin
    case (exp_381)
      0:exp_536_reg <= exp_534;
      1:exp_536_reg <= exp_533;
      default:exp_536_reg <= exp_535;
    endcase
  end
  assign exp_536 = exp_536_reg;
  assign exp_381 = exp_362 == exp_380;
  assign exp_380 = 99;
  assign exp_535 = 0;
  assign exp_534 = 0;

  reg [0:0] exp_533_reg;
  always@(*) begin
    case (exp_363)
      0:exp_533_reg <= exp_516;
      1:exp_533_reg <= exp_517;
      2:exp_533_reg <= exp_530;
      3:exp_533_reg <= exp_531;
      4:exp_533_reg <= exp_518;
      5:exp_533_reg <= exp_519;
      6:exp_533_reg <= exp_524;
      7:exp_533_reg <= exp_529;
      default:exp_533_reg <= exp_532;
    endcase
  end
  assign exp_533 = exp_533_reg;
  assign exp_363 = exp_360[14:12];
  assign exp_532 = 0;
  assign exp_516 = exp_352 == exp_353;

      reg [31:0] exp_352_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_352_reg <= exp_290;
        end
      end
      assign exp_352 = exp_352_reg;
    
  reg [31:0] exp_290_reg;
  always@(*) begin
    case (exp_286)
      0:exp_290_reg <= exp_282;
      1:exp_290_reg <= exp_288;
      default:exp_290_reg <= exp_289;
    endcase
  end
  assign exp_290 = exp_290_reg;
  assign exp_286 = exp_266 == exp_285;
  assign exp_266 = exp_96[19:15];
  assign exp_285 = 0;
  assign exp_289 = 0;

  reg [31:0] exp_282_reg;
  always@(*) begin
    case (exp_263)
      0:exp_282_reg <= exp_253;
      1:exp_282_reg <= exp_265;
      default:exp_282_reg <= exp_281;
    endcase
  end
  assign exp_282 = exp_282_reg;
  assign exp_263 = exp_836;
  assign exp_836 = exp_835 & exp_232;
  assign exp_835 = exp_834 & exp_240;
  assign exp_834 = exp_833 & exp_827;
  assign exp_833 = exp_245 == exp_828;
  assign exp_245 = exp_96[19:15];
  assign exp_828 = exp_360[11:7];
  assign exp_827 = exp_419 | exp_822;
  assign exp_419 = exp_418 | exp_377;
  assign exp_418 = exp_417 | exp_371;
  assign exp_417 = exp_416 | exp_369;
  assign exp_416 = exp_415 | exp_375;
  assign exp_415 = exp_414 | exp_373;
  assign exp_414 = exp_365 | exp_367;
  assign exp_365 = exp_362 == exp_364;
  assign exp_364 = 19;
  assign exp_367 = exp_362 == exp_366;
  assign exp_366 = 51;
  assign exp_369 = exp_362 == exp_368;
  assign exp_368 = 55;
  assign exp_371 = exp_362 == exp_370;
  assign exp_370 = 23;
  assign exp_822 = exp_821 & exp_581;

  reg [0:0] exp_821_reg;
  always@(*) begin
    case (exp_607)
      0:exp_821_reg <= exp_818;
      1:exp_821_reg <= exp_819;
      default:exp_821_reg <= exp_820;
    endcase
  end
  assign exp_821 = exp_821_reg;
  assign exp_607 = exp_581 & exp_606;
  assign exp_581 = exp_579 & exp_580;
  assign exp_579 = exp_577 == exp_578;
  assign exp_577 = exp_360[6:0];
  assign exp_578 = 51;
  assign exp_580 = exp_360[25:25];
  assign exp_606 = exp_576[2:2];
  assign exp_576 = exp_360[14:12];
  assign exp_820 = 0;
  assign exp_818 = exp_811 & exp_581;
  assign exp_811 = exp_726 == exp_810;

      reg [2:0] exp_726_reg = 0;
      always@(posedge clk) begin
        if (exp_722) begin
          exp_726_reg <= exp_733;
        end
      end
      assign exp_726 = exp_726_reg;
    
  reg [2:0] exp_733_reg;
  always@(*) begin
    case (exp_728)
      0:exp_733_reg <= exp_730;
      1:exp_733_reg <= exp_731;
      default:exp_733_reg <= exp_732;
    endcase
  end
  assign exp_733 = exp_733_reg;
  assign exp_728 = exp_726 == exp_727;
  assign exp_727 = 4;
  assign exp_732 = 0;
  assign exp_730 = exp_726 + exp_729;
  assign exp_729 = 1;
  assign exp_731 = 0;
  assign exp_722 = exp_581 & exp_721;
  assign exp_721 = ~exp_720;
  assign exp_720 = exp_576[2:2];
  assign exp_810 = 4;
  assign exp_819 = exp_629 & exp_581;
  assign exp_629 = exp_613 == exp_628;

      reg [5:0] exp_613_reg = 0;
      always@(posedge clk) begin
        if (exp_607) begin
          exp_613_reg <= exp_620;
        end
      end
      assign exp_613 = exp_613_reg;
    
  reg [5:0] exp_620_reg;
  always@(*) begin
    case (exp_615)
      0:exp_620_reg <= exp_617;
      1:exp_620_reg <= exp_618;
      default:exp_620_reg <= exp_619;
    endcase
  end
  assign exp_620 = exp_620_reg;
  assign exp_615 = exp_613 == exp_614;
  assign exp_614 = 37;
  assign exp_619 = 0;
  assign exp_617 = exp_613 + exp_616;
  assign exp_616 = 1;
  assign exp_618 = 0;
  assign exp_628 = 37;

      reg [0:0] exp_240_reg = 0;
      always@(posedge clk) begin
        if (exp_232) begin
          exp_240_reg <= exp_239;
        end
      end
      assign exp_240 = exp_240_reg;
      assign exp_239 = exp_237 & exp_238;

      reg [0:0] exp_237_reg = 0;
      always@(posedge clk) begin
        if (exp_232) begin
          exp_237_reg <= exp_236;
        end
      end
      assign exp_237 = exp_237_reg;
      assign exp_236 = exp_234 & exp_235;
  assign exp_234 = 1;
  assign exp_235 = ~exp_233;
  assign exp_233 = exp_846;
  assign exp_846 = exp_240 & exp_537;
  assign exp_232 = ~exp_231;
  assign exp_231 = exp_850;
  assign exp_850 = exp_240 & exp_849;
  assign exp_849 = exp_848 | exp_824;
  assign exp_848 = exp_228 & exp_847;
  assign exp_847 = ~exp_227;
  assign exp_227 = exp_218;

  reg [0:0] exp_218_reg;
  always@(*) begin
    case (exp_213)
      0:exp_218_reg <= exp_196;
      1:exp_218_reg <= exp_205;
      default:exp_218_reg <= exp_217;
    endcase
  end
  assign exp_218 = exp_218_reg;
  assign exp_213 = exp_210 & exp_212;
  assign exp_210 = exp_1 >= exp_209;
  assign exp_1 = exp_224;
  assign exp_224 = exp_431;
  assign exp_431 = exp_430 + exp_429;
  assign exp_430 = 0;
  assign exp_429 = exp_352 + exp_428;
  assign exp_428 = $signed(exp_427);
  assign exp_427 = exp_426 + exp_425;
  assign exp_426 = 0;

  reg [11:0] exp_425_reg;
  always@(*) begin
    case (exp_379)
      0:exp_425_reg <= exp_420;
      1:exp_425_reg <= exp_423;
      default:exp_425_reg <= exp_424;
    endcase
  end
  assign exp_425 = exp_425_reg;
  assign exp_379 = exp_362 == exp_378;
  assign exp_378 = 35;
  assign exp_424 = 0;
  assign exp_420 = exp_360[31:20];
  assign exp_423 = {exp_421, exp_422};  assign exp_421 = exp_360[31:25];
  assign exp_422 = exp_360[11:7];
  assign exp_209 = 2147483660;
  assign exp_212 = exp_1 <= exp_211;
  assign exp_211 = 2147483660;
  assign exp_217 = 0;

  reg [0:0] exp_196_reg;
  always@(*) begin
    case (exp_191)
      0:exp_196_reg <= exp_155;
      1:exp_196_reg <= exp_183;
      default:exp_196_reg <= exp_195;
    endcase
  end
  assign exp_196 = exp_196_reg;
  assign exp_191 = exp_188 & exp_190;
  assign exp_188 = exp_1 >= exp_187;
  assign exp_187 = 2147483656;
  assign exp_190 = exp_1 <= exp_189;
  assign exp_189 = 2147483656;
  assign exp_195 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 2147483648;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 2147483652;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 8188;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_229;
  assign exp_229 = exp_514;
  assign exp_514 = exp_513 + exp_379;
  assign exp_513 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_176;
  assign exp_176 = 1;
  assign exp_183 = exp_198;
  assign exp_198 = stdout_ready_in;
  assign exp_205 = exp_221;
  assign exp_221 = stdin_valid_in;
  assign exp_824 = exp_581 & exp_823;
  assign exp_823 = ~exp_821;
  assign exp_238 = ~exp_233;
  assign exp_281 = 0;

  //Create RAM
  reg [31:0] exp_253_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_251) begin
      exp_253_ram[exp_247] <= exp_249;
    end
  end
  assign exp_253 = exp_253_ram[exp_248];
  assign exp_252 = exp_261;
  assign exp_261 = 1;
  assign exp_248 = exp_245;
  assign exp_251 = exp_830;
  assign exp_830 = exp_829 & exp_232;
  assign exp_829 = exp_827 & exp_240;
  assign exp_247 = exp_828;
  assign exp_249 = exp_826;

  reg [31:0] exp_826_reg;
  always@(*) begin
    case (exp_822)
      0:exp_826_reg <= exp_462;
      1:exp_826_reg <= exp_817;
      default:exp_826_reg <= exp_825;
    endcase
  end
  assign exp_826 = exp_826_reg;
  assign exp_825 = 0;

  reg [31:0] exp_462_reg;
  always@(*) begin
    case (exp_377)
      0:exp_462_reg <= exp_413;
      1:exp_462_reg <= exp_460;
      default:exp_462_reg <= exp_461;
    endcase
  end
  assign exp_462 = exp_462_reg;
  assign exp_461 = 0;

  reg [31:0] exp_413_reg;
  always@(*) begin
    case (exp_356)
      0:exp_413_reg <= exp_392;
      1:exp_413_reg <= exp_394;
      2:exp_413_reg <= exp_410;
      3:exp_413_reg <= exp_411;
      4:exp_413_reg <= exp_403;
      5:exp_413_reg <= exp_407;
      6:exp_413_reg <= exp_408;
      7:exp_413_reg <= exp_409;
      default:exp_413_reg <= exp_412;
    endcase
  end
  assign exp_413 = exp_413_reg;

      reg [2:0] exp_356_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_356_reg <= exp_347;
        end
      end
      assign exp_356 = exp_356_reg;
    
  reg [2:0] exp_347_reg;
  always@(*) begin
    case (exp_344)
      0:exp_347_reg <= exp_334;
      1:exp_347_reg <= exp_345;
      default:exp_347_reg <= exp_346;
    endcase
  end
  assign exp_347 = exp_347_reg;
  assign exp_344 = exp_278 | exp_280;
  assign exp_278 = exp_268 == exp_277;
  assign exp_268 = exp_96[6:0];
  assign exp_277 = 111;
  assign exp_280 = exp_268 == exp_279;
  assign exp_279 = 103;
  assign exp_346 = 0;

  reg [2:0] exp_334_reg;
  always@(*) begin
    case (exp_276)
      0:exp_334_reg <= exp_321;
      1:exp_334_reg <= exp_332;
      default:exp_334_reg <= exp_333;
    endcase
  end
  assign exp_334 = exp_334_reg;
  assign exp_276 = exp_268 == exp_275;
  assign exp_275 = 23;
  assign exp_333 = 0;

  reg [2:0] exp_321_reg;
  always@(*) begin
    case (exp_274)
      0:exp_321_reg <= exp_270;
      1:exp_321_reg <= exp_319;
      default:exp_321_reg <= exp_320;
    endcase
  end
  assign exp_321 = exp_321_reg;
  assign exp_274 = exp_268 == exp_273;
  assign exp_273 = 55;
  assign exp_320 = 0;
  assign exp_270 = exp_96[14:12];
  assign exp_319 = 0;
  assign exp_332 = 0;
  assign exp_345 = 0;
  assign exp_351 = exp_232 & exp_237;
  assign exp_412 = 0;

  reg [31:0] exp_392_reg;
  always@(*) begin
    case (exp_358)
      0:exp_392_reg <= exp_389;
      1:exp_392_reg <= exp_390;
      default:exp_392_reg <= exp_391;
    endcase
  end
  assign exp_392 = exp_392_reg;

      reg [0:0] exp_358_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_358_reg <= exp_350;
        end
      end
      assign exp_358 = exp_358_reg;
      assign exp_350 = exp_336 & exp_349;
  assign exp_336 = exp_323 & exp_335;
  assign exp_323 = exp_309 & exp_322;
  assign exp_309 = exp_307 & exp_308;
  assign exp_307 = exp_96[30:30];
  assign exp_308 = ~exp_272;
  assign exp_272 = exp_268 == exp_271;
  assign exp_271 = 19;
  assign exp_322 = ~exp_274;
  assign exp_335 = ~exp_276;
  assign exp_349 = ~exp_348;
  assign exp_348 = exp_278 | exp_280;
  assign exp_391 = 0;
  assign exp_389 = exp_354 + exp_355;

      reg [31:0] exp_354_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_354_reg <= exp_340;
        end
      end
      assign exp_354 = exp_354_reg;
    
  reg [31:0] exp_340_reg;
  always@(*) begin
    case (exp_337)
      0:exp_340_reg <= exp_329;
      1:exp_340_reg <= exp_338;
      default:exp_340_reg <= exp_339;
    endcase
  end
  assign exp_340 = exp_340_reg;
  assign exp_337 = exp_278 | exp_280;
  assign exp_339 = 0;

  reg [31:0] exp_329_reg;
  always@(*) begin
    case (exp_276)
      0:exp_329_reg <= exp_315;
      1:exp_329_reg <= exp_327;
      default:exp_329_reg <= exp_328;
    endcase
  end
  assign exp_329 = exp_329_reg;
  assign exp_328 = 0;

  reg [31:0] exp_315_reg;
  always@(*) begin
    case (exp_274)
      0:exp_315_reg <= exp_290;
      1:exp_315_reg <= exp_313;
      default:exp_315_reg <= exp_314;
    endcase
  end
  assign exp_315 = exp_315_reg;
  assign exp_314 = 0;
  assign exp_313 = exp_311 << exp_312;
  assign exp_311 = exp_310;
  assign exp_310 = exp_96[31:12];
  assign exp_312 = 12;
  assign exp_327 = exp_325 << exp_326;
  assign exp_325 = exp_324;
  assign exp_324 = exp_96[31:12];
  assign exp_326 = 12;
  assign exp_338 = 4;

      reg [31:0] exp_355_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_355_reg <= exp_343;
        end
      end
      assign exp_355 = exp_355_reg;
    
  reg [31:0] exp_343_reg;
  always@(*) begin
    case (exp_341)
      0:exp_343_reg <= exp_331;
      1:exp_343_reg <= exp_244;
      default:exp_343_reg <= exp_342;
    endcase
  end
  assign exp_343 = exp_343_reg;
  assign exp_341 = exp_278 | exp_280;
  assign exp_342 = 0;

  reg [31:0] exp_331_reg;
  always@(*) begin
    case (exp_276)
      0:exp_331_reg <= exp_318;
      1:exp_331_reg <= exp_244;
      default:exp_331_reg <= exp_330;
    endcase
  end
  assign exp_331 = exp_331_reg;
  assign exp_330 = 0;

  reg [31:0] exp_318_reg;
  always@(*) begin
    case (exp_274)
      0:exp_318_reg <= exp_302;
      1:exp_318_reg <= exp_316;
      default:exp_318_reg <= exp_317;
    endcase
  end
  assign exp_318 = exp_318_reg;
  assign exp_317 = 0;

  reg [31:0] exp_302_reg;
  always@(*) begin
    case (exp_272)
      0:exp_302_reg <= exp_296;
      1:exp_302_reg <= exp_300;
      default:exp_302_reg <= exp_301;
    endcase
  end
  assign exp_302 = exp_302_reg;
  assign exp_301 = 0;

  reg [31:0] exp_296_reg;
  always@(*) begin
    case (exp_292)
      0:exp_296_reg <= exp_284;
      1:exp_296_reg <= exp_294;
      default:exp_296_reg <= exp_295;
    endcase
  end
  assign exp_296 = exp_296_reg;
  assign exp_292 = exp_267 == exp_291;
  assign exp_267 = exp_96[24:20];
  assign exp_291 = 0;
  assign exp_295 = 0;

  reg [31:0] exp_284_reg;
  always@(*) begin
    case (exp_264)
      0:exp_284_reg <= exp_260;
      1:exp_284_reg <= exp_265;
      default:exp_284_reg <= exp_283;
    endcase
  end
  assign exp_284 = exp_284_reg;
  assign exp_264 = exp_840;
  assign exp_840 = exp_839 & exp_232;
  assign exp_839 = exp_838 & exp_240;
  assign exp_838 = exp_837 & exp_827;
  assign exp_837 = exp_246 == exp_828;
  assign exp_246 = exp_96[24:20];
  assign exp_283 = 0;

  //Create RAM
  reg [31:0] exp_260_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_258) begin
      exp_260_ram[exp_254] <= exp_256;
    end
  end
  assign exp_260 = exp_260_ram[exp_255];
  assign exp_259 = exp_262;
  assign exp_262 = 1;
  assign exp_255 = exp_246;
  assign exp_258 = exp_832;
  assign exp_832 = exp_831 & exp_232;
  assign exp_831 = exp_827 & exp_240;
  assign exp_254 = exp_828;
  assign exp_256 = exp_826;
  assign exp_265 = exp_826;
  assign exp_294 = $signed(exp_293);
  assign exp_293 = 0;
  assign exp_300 = exp_297 + exp_299;
  assign exp_297 = 0;
  assign exp_299 = $signed(exp_298);
  assign exp_298 = exp_96[31:20];
  assign exp_316 = 0;

      reg [31:0] exp_244_reg = 0;
      always@(posedge clk) begin
        if (exp_243) begin
          exp_244_reg <= exp_242;
        end
      end
      assign exp_244 = exp_244_reg;
      assign exp_243 = exp_234 & exp_232;
  assign exp_390 = exp_354 - exp_355;
  assign exp_394 = exp_354 << exp_393;
  assign exp_393 = $signed(exp_388);
  assign exp_388 = exp_387 + exp_386;
  assign exp_387 = 0;
  assign exp_386 = exp_357;

      reg [4:0] exp_357_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_357_reg <= exp_306;
        end
      end
      assign exp_357 = exp_357_reg;
    
  reg [4:0] exp_306_reg;
  always@(*) begin
    case (exp_272)
      0:exp_306_reg <= exp_304;
      1:exp_306_reg <= exp_269;
      default:exp_306_reg <= exp_305;
    endcase
  end
  assign exp_306 = exp_306_reg;
  assign exp_305 = 0;
  assign exp_304 = exp_302[4:0];
  assign exp_269 = exp_96[24:20];
  assign exp_410 = $signed(exp_396);
  assign exp_396 = exp_395;
  assign exp_395 = $signed(exp_354) < $signed(exp_355);
  assign exp_411 = $signed(exp_402);
  assign exp_402 = exp_401;
  assign exp_401 = exp_398 < exp_400;
  assign exp_398 = exp_397 + exp_354;
  assign exp_397 = 0;
  assign exp_400 = exp_399 + exp_355;
  assign exp_399 = 0;
  assign exp_403 = exp_354 ^ exp_355;
  assign exp_407 = exp_406[31:0];
  assign exp_406 = $signed(exp_404) >>> $signed(exp_405);
  assign exp_404 = {exp_385, exp_354};
  reg [0:0] exp_385_reg;
  always@(*) begin
    case (exp_359)
      0:exp_385_reg <= exp_383;
      1:exp_385_reg <= exp_382;
      default:exp_385_reg <= exp_384;
    endcase
  end
  assign exp_385 = exp_385_reg;

      reg [0:0] exp_359_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_359_reg <= exp_303;
        end
      end
      assign exp_359 = exp_359_reg;
      assign exp_303 = exp_96[30:30];
  assign exp_384 = 0;
  assign exp_383 = 0;
  assign exp_382 = exp_354[31:31];
  assign exp_405 = $signed(exp_388);
  assign exp_408 = exp_354 | exp_355;
  assign exp_409 = exp_354 & exp_355;

  reg [31:0] exp_460_reg;
  always@(*) begin
    case (exp_363)
      0:exp_460_reg <= exp_450;
      1:exp_460_reg <= exp_453;
      2:exp_460_reg <= exp_226;
      3:exp_460_reg <= exp_454;
      4:exp_460_reg <= exp_455;
      5:exp_460_reg <= exp_456;
      6:exp_460_reg <= exp_457;
      7:exp_460_reg <= exp_458;
      default:exp_460_reg <= exp_459;
    endcase
  end
  assign exp_460 = exp_460_reg;
  assign exp_459 = 0;
  assign exp_450 = $signed(exp_449);
  assign exp_449 = exp_448 + exp_443;
  assign exp_448 = 0;

  reg [7:0] exp_443_reg;
  always@(*) begin
    case (exp_434)
      0:exp_443_reg <= exp_438;
      1:exp_443_reg <= exp_439;
      2:exp_443_reg <= exp_440;
      3:exp_443_reg <= exp_441;
      default:exp_443_reg <= exp_442;
    endcase
  end
  assign exp_443 = exp_443_reg;
  assign exp_434 = exp_433 + exp_432;
  assign exp_433 = 0;
  assign exp_432 = exp_431[1:0];
  assign exp_442 = 0;
  assign exp_438 = exp_226[7:0];
  assign exp_226 = exp_216;

  reg [31:0] exp_216_reg;
  always@(*) begin
    case (exp_213)
      0:exp_216_reg <= exp_194;
      1:exp_216_reg <= exp_204;
      default:exp_216_reg <= exp_215;
    endcase
  end
  assign exp_216 = exp_216_reg;
  assign exp_215 = 0;

  reg [31:0] exp_194_reg;
  always@(*) begin
    case (exp_191)
      0:exp_194_reg <= exp_153;
      1:exp_194_reg <= exp_182;
      default:exp_194_reg <= exp_193;
    endcase
  end
  assign exp_194 = exp_194_reg;
  assign exp_193 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 0;
    exp_54_ram[32] = 252;
    exp_54_ram[33] = 47;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 108;
    exp_54_ram[36] = 111;
    exp_54_ram[37] = 33;
    exp_54_ram[38] = 0;
    exp_54_ram[39] = 253;
    exp_54_ram[40] = 2;
    exp_54_ram[41] = 3;
    exp_54_ram[42] = 252;
    exp_54_ram[43] = 252;
    exp_54_ram[44] = 253;
    exp_54_ram[45] = 254;
    exp_54_ram[46] = 253;
    exp_54_ram[47] = 254;
    exp_54_ram[48] = 0;
    exp_54_ram[49] = 253;
    exp_54_ram[50] = 0;
    exp_54_ram[51] = 2;
    exp_54_ram[52] = 3;
    exp_54_ram[53] = 0;
    exp_54_ram[54] = 254;
    exp_54_ram[55] = 0;
    exp_54_ram[56] = 2;
    exp_54_ram[57] = 0;
    exp_54_ram[58] = 254;
    exp_54_ram[59] = 254;
    exp_54_ram[60] = 254;
    exp_54_ram[61] = 254;
    exp_54_ram[62] = 0;
    exp_54_ram[63] = 1;
    exp_54_ram[64] = 2;
    exp_54_ram[65] = 0;
    exp_54_ram[66] = 254;
    exp_54_ram[67] = 0;
    exp_54_ram[68] = 0;
    exp_54_ram[69] = 2;
    exp_54_ram[70] = 0;
    exp_54_ram[71] = 254;
    exp_54_ram[72] = 254;
    exp_54_ram[73] = 254;
    exp_54_ram[74] = 254;
    exp_54_ram[75] = 254;
    exp_54_ram[76] = 0;
    exp_54_ram[77] = 254;
    exp_54_ram[78] = 0;
    exp_54_ram[79] = 31;
    exp_54_ram[80] = 0;
    exp_54_ram[81] = 1;
    exp_54_ram[82] = 1;
    exp_54_ram[83] = 2;
    exp_54_ram[84] = 0;
    exp_54_ram[85] = 253;
    exp_54_ram[86] = 2;
    exp_54_ram[87] = 3;
    exp_54_ram[88] = 252;
    exp_54_ram[89] = 252;
    exp_54_ram[90] = 253;
    exp_54_ram[91] = 254;
    exp_54_ram[92] = 1;
    exp_54_ram[93] = 254;
    exp_54_ram[94] = 0;
    exp_54_ram[95] = 254;
    exp_54_ram[96] = 254;
    exp_54_ram[97] = 0;
    exp_54_ram[98] = 0;
    exp_54_ram[99] = 253;
    exp_54_ram[100] = 255;
    exp_54_ram[101] = 252;
    exp_54_ram[102] = 252;
    exp_54_ram[103] = 254;
    exp_54_ram[104] = 253;
    exp_54_ram[105] = 64;
    exp_54_ram[106] = 0;
    exp_54_ram[107] = 2;
    exp_54_ram[108] = 3;
    exp_54_ram[109] = 0;
    exp_54_ram[110] = 254;
    exp_54_ram[111] = 0;
    exp_54_ram[112] = 2;
    exp_54_ram[113] = 0;
    exp_54_ram[114] = 254;
    exp_54_ram[115] = 254;
    exp_54_ram[116] = 2;
    exp_54_ram[117] = 0;
    exp_54_ram[118] = 254;
    exp_54_ram[119] = 3;
    exp_54_ram[120] = 0;
    exp_54_ram[121] = 0;
    exp_54_ram[122] = 0;
    exp_54_ram[123] = 0;
    exp_54_ram[124] = 0;
    exp_54_ram[125] = 15;
    exp_54_ram[126] = 0;
    exp_54_ram[127] = 1;
    exp_54_ram[128] = 2;
    exp_54_ram[129] = 0;
    exp_54_ram[130] = 253;
    exp_54_ram[131] = 2;
    exp_54_ram[132] = 2;
    exp_54_ram[133] = 3;
    exp_54_ram[134] = 252;
    exp_54_ram[135] = 254;
    exp_54_ram[136] = 4;
    exp_54_ram[137] = 254;
    exp_54_ram[138] = 0;
    exp_54_ram[139] = 0;
    exp_54_ram[140] = 0;
    exp_54_ram[141] = 0;
    exp_54_ram[142] = 0;
    exp_54_ram[143] = 253;
    exp_54_ram[144] = 0;
    exp_54_ram[145] = 0;
    exp_54_ram[146] = 253;
    exp_54_ram[147] = 0;
    exp_54_ram[148] = 0;
    exp_54_ram[149] = 0;
    exp_54_ram[150] = 253;
    exp_54_ram[151] = 254;
    exp_54_ram[152] = 253;
    exp_54_ram[153] = 0;
    exp_54_ram[154] = 0;
    exp_54_ram[155] = 0;
    exp_54_ram[156] = 244;
    exp_54_ram[157] = 0;
    exp_54_ram[158] = 250;
    exp_54_ram[159] = 254;
    exp_54_ram[160] = 0;
    exp_54_ram[161] = 2;
    exp_54_ram[162] = 2;
    exp_54_ram[163] = 3;
    exp_54_ram[164] = 0;
    exp_54_ram[165] = 252;
    exp_54_ram[166] = 2;
    exp_54_ram[167] = 2;
    exp_54_ram[168] = 4;
    exp_54_ram[169] = 252;
    exp_54_ram[170] = 252;
    exp_54_ram[171] = 252;
    exp_54_ram[172] = 252;
    exp_54_ram[173] = 252;
    exp_54_ram[174] = 252;
    exp_54_ram[175] = 253;
    exp_54_ram[176] = 253;
    exp_54_ram[177] = 253;
    exp_54_ram[178] = 254;
    exp_54_ram[179] = 252;
    exp_54_ram[180] = 0;
    exp_54_ram[181] = 8;
    exp_54_ram[182] = 252;
    exp_54_ram[183] = 0;
    exp_54_ram[184] = 8;
    exp_54_ram[185] = 252;
    exp_54_ram[186] = 254;
    exp_54_ram[187] = 3;
    exp_54_ram[188] = 253;
    exp_54_ram[189] = 0;
    exp_54_ram[190] = 252;
    exp_54_ram[191] = 253;
    exp_54_ram[192] = 253;
    exp_54_ram[193] = 0;
    exp_54_ram[194] = 253;
    exp_54_ram[195] = 2;
    exp_54_ram[196] = 0;
    exp_54_ram[197] = 254;
    exp_54_ram[198] = 0;
    exp_54_ram[199] = 254;
    exp_54_ram[200] = 254;
    exp_54_ram[201] = 252;
    exp_54_ram[202] = 252;
    exp_54_ram[203] = 4;
    exp_54_ram[204] = 252;
    exp_54_ram[205] = 255;
    exp_54_ram[206] = 252;
    exp_54_ram[207] = 252;
    exp_54_ram[208] = 252;
    exp_54_ram[209] = 0;
    exp_54_ram[210] = 0;
    exp_54_ram[211] = 253;
    exp_54_ram[212] = 0;
    exp_54_ram[213] = 252;
    exp_54_ram[214] = 253;
    exp_54_ram[215] = 253;
    exp_54_ram[216] = 0;
    exp_54_ram[217] = 253;
    exp_54_ram[218] = 0;
    exp_54_ram[219] = 252;
    exp_54_ram[220] = 252;
    exp_54_ram[221] = 252;
    exp_54_ram[222] = 0;
    exp_54_ram[223] = 4;
    exp_54_ram[224] = 2;
    exp_54_ram[225] = 253;
    exp_54_ram[226] = 0;
    exp_54_ram[227] = 252;
    exp_54_ram[228] = 253;
    exp_54_ram[229] = 253;
    exp_54_ram[230] = 0;
    exp_54_ram[231] = 253;
    exp_54_ram[232] = 2;
    exp_54_ram[233] = 0;
    exp_54_ram[234] = 253;
    exp_54_ram[235] = 254;
    exp_54_ram[236] = 64;
    exp_54_ram[237] = 252;
    exp_54_ram[238] = 252;
    exp_54_ram[239] = 253;
    exp_54_ram[240] = 0;
    exp_54_ram[241] = 3;
    exp_54_ram[242] = 3;
    exp_54_ram[243] = 4;
    exp_54_ram[244] = 0;
    exp_54_ram[245] = 253;
    exp_54_ram[246] = 2;
    exp_54_ram[247] = 2;
    exp_54_ram[248] = 3;
    exp_54_ram[249] = 254;
    exp_54_ram[250] = 254;
    exp_54_ram[251] = 254;
    exp_54_ram[252] = 254;
    exp_54_ram[253] = 252;
    exp_54_ram[254] = 252;
    exp_54_ram[255] = 0;
    exp_54_ram[256] = 253;
    exp_54_ram[257] = 252;
    exp_54_ram[258] = 0;
    exp_54_ram[259] = 0;
    exp_54_ram[260] = 10;
    exp_54_ram[261] = 0;
    exp_54_ram[262] = 4;
    exp_54_ram[263] = 0;
    exp_54_ram[264] = 0;
    exp_54_ram[265] = 4;
    exp_54_ram[266] = 253;
    exp_54_ram[267] = 0;
    exp_54_ram[268] = 0;
    exp_54_ram[269] = 0;
    exp_54_ram[270] = 2;
    exp_54_ram[271] = 0;
    exp_54_ram[272] = 255;
    exp_54_ram[273] = 0;
    exp_54_ram[274] = 2;
    exp_54_ram[275] = 253;
    exp_54_ram[276] = 0;
    exp_54_ram[277] = 252;
    exp_54_ram[278] = 253;
    exp_54_ram[279] = 0;
    exp_54_ram[280] = 3;
    exp_54_ram[281] = 0;
    exp_54_ram[282] = 253;
    exp_54_ram[283] = 0;
    exp_54_ram[284] = 2;
    exp_54_ram[285] = 253;
    exp_54_ram[286] = 1;
    exp_54_ram[287] = 252;
    exp_54_ram[288] = 2;
    exp_54_ram[289] = 253;
    exp_54_ram[290] = 0;
    exp_54_ram[291] = 252;
    exp_54_ram[292] = 253;
    exp_54_ram[293] = 0;
    exp_54_ram[294] = 3;
    exp_54_ram[295] = 0;
    exp_54_ram[296] = 0;
    exp_54_ram[297] = 0;
    exp_54_ram[298] = 0;
    exp_54_ram[299] = 253;
    exp_54_ram[300] = 0;
    exp_54_ram[301] = 0;
    exp_54_ram[302] = 253;
    exp_54_ram[303] = 1;
    exp_54_ram[304] = 252;
    exp_54_ram[305] = 0;
    exp_54_ram[306] = 1;
    exp_54_ram[307] = 20;
    exp_54_ram[308] = 0;
    exp_54_ram[309] = 64;
    exp_54_ram[310] = 4;
    exp_54_ram[311] = 253;
    exp_54_ram[312] = 4;
    exp_54_ram[313] = 253;
    exp_54_ram[314] = 0;
    exp_54_ram[315] = 0;
    exp_54_ram[316] = 253;
    exp_54_ram[317] = 0;
    exp_54_ram[318] = 2;
    exp_54_ram[319] = 253;
    exp_54_ram[320] = 255;
    exp_54_ram[321] = 252;
    exp_54_ram[322] = 253;
    exp_54_ram[323] = 0;
    exp_54_ram[324] = 253;
    exp_54_ram[325] = 1;
    exp_54_ram[326] = 0;
    exp_54_ram[327] = 253;
    exp_54_ram[328] = 255;
    exp_54_ram[329] = 252;
    exp_54_ram[330] = 253;
    exp_54_ram[331] = 1;
    exp_54_ram[332] = 2;
    exp_54_ram[333] = 0;
    exp_54_ram[334] = 2;
    exp_54_ram[335] = 2;
    exp_54_ram[336] = 253;
    exp_54_ram[337] = 1;
    exp_54_ram[338] = 2;
    exp_54_ram[339] = 253;
    exp_54_ram[340] = 0;
    exp_54_ram[341] = 252;
    exp_54_ram[342] = 253;
    exp_54_ram[343] = 0;
    exp_54_ram[344] = 7;
    exp_54_ram[345] = 0;
    exp_54_ram[346] = 7;
    exp_54_ram[347] = 253;
    exp_54_ram[348] = 1;
    exp_54_ram[349] = 2;
    exp_54_ram[350] = 0;
    exp_54_ram[351] = 2;
    exp_54_ram[352] = 2;
    exp_54_ram[353] = 253;
    exp_54_ram[354] = 1;
    exp_54_ram[355] = 2;
    exp_54_ram[356] = 253;
    exp_54_ram[357] = 0;
    exp_54_ram[358] = 252;
    exp_54_ram[359] = 253;
    exp_54_ram[360] = 0;
    exp_54_ram[361] = 5;
    exp_54_ram[362] = 0;
    exp_54_ram[363] = 3;
    exp_54_ram[364] = 253;
    exp_54_ram[365] = 0;
    exp_54_ram[366] = 2;
    exp_54_ram[367] = 253;
    exp_54_ram[368] = 1;
    exp_54_ram[369] = 2;
    exp_54_ram[370] = 253;
    exp_54_ram[371] = 0;
    exp_54_ram[372] = 252;
    exp_54_ram[373] = 253;
    exp_54_ram[374] = 0;
    exp_54_ram[375] = 6;
    exp_54_ram[376] = 0;
    exp_54_ram[377] = 253;
    exp_54_ram[378] = 1;
    exp_54_ram[379] = 2;
    exp_54_ram[380] = 253;
    exp_54_ram[381] = 0;
    exp_54_ram[382] = 252;
    exp_54_ram[383] = 253;
    exp_54_ram[384] = 0;
    exp_54_ram[385] = 3;
    exp_54_ram[386] = 0;
    exp_54_ram[387] = 253;
    exp_54_ram[388] = 1;
    exp_54_ram[389] = 8;
    exp_54_ram[390] = 253;
    exp_54_ram[391] = 2;
    exp_54_ram[392] = 253;
    exp_54_ram[393] = 0;
    exp_54_ram[394] = 252;
    exp_54_ram[395] = 253;
    exp_54_ram[396] = 0;
    exp_54_ram[397] = 2;
    exp_54_ram[398] = 0;
    exp_54_ram[399] = 5;
    exp_54_ram[400] = 0;
    exp_54_ram[401] = 0;
    exp_54_ram[402] = 2;
    exp_54_ram[403] = 253;
    exp_54_ram[404] = 0;
    exp_54_ram[405] = 252;
    exp_54_ram[406] = 253;
    exp_54_ram[407] = 0;
    exp_54_ram[408] = 2;
    exp_54_ram[409] = 0;
    exp_54_ram[410] = 2;
    exp_54_ram[411] = 0;
    exp_54_ram[412] = 0;
    exp_54_ram[413] = 2;
    exp_54_ram[414] = 253;
    exp_54_ram[415] = 0;
    exp_54_ram[416] = 252;
    exp_54_ram[417] = 253;
    exp_54_ram[418] = 0;
    exp_54_ram[419] = 2;
    exp_54_ram[420] = 0;
    exp_54_ram[421] = 0;
    exp_54_ram[422] = 0;
    exp_54_ram[423] = 253;
    exp_54_ram[424] = 253;
    exp_54_ram[425] = 254;
    exp_54_ram[426] = 254;
    exp_54_ram[427] = 254;
    exp_54_ram[428] = 254;
    exp_54_ram[429] = 190;
    exp_54_ram[430] = 0;
    exp_54_ram[431] = 0;
    exp_54_ram[432] = 2;
    exp_54_ram[433] = 2;
    exp_54_ram[434] = 3;
    exp_54_ram[435] = 0;
    exp_54_ram[436] = 249;
    exp_54_ram[437] = 6;
    exp_54_ram[438] = 6;
    exp_54_ram[439] = 7;
    exp_54_ram[440] = 250;
    exp_54_ram[441] = 250;
    exp_54_ram[442] = 250;
    exp_54_ram[443] = 250;
    exp_54_ram[444] = 250;
    exp_54_ram[445] = 251;
    exp_54_ram[446] = 251;
    exp_54_ram[447] = 250;
    exp_54_ram[448] = 254;
    exp_54_ram[449] = 250;
    exp_54_ram[450] = 0;
    exp_54_ram[451] = 0;
    exp_54_ram[452] = 254;
    exp_54_ram[453] = 0;
    exp_54_ram[454] = 0;
    exp_54_ram[455] = 64;
    exp_54_ram[456] = 0;
    exp_54_ram[457] = 250;
    exp_54_ram[458] = 8;
    exp_54_ram[459] = 250;
    exp_54_ram[460] = 250;
    exp_54_ram[461] = 2;
    exp_54_ram[462] = 254;
    exp_54_ram[463] = 254;
    exp_54_ram[464] = 0;
    exp_54_ram[465] = 0;
    exp_54_ram[466] = 254;
    exp_54_ram[467] = 3;
    exp_54_ram[468] = 15;
    exp_54_ram[469] = 3;
    exp_54_ram[470] = 0;
    exp_54_ram[471] = 2;
    exp_54_ram[472] = 0;
    exp_54_ram[473] = 4;
    exp_54_ram[474] = 0;
    exp_54_ram[475] = 6;
    exp_54_ram[476] = 254;
    exp_54_ram[477] = 0;
    exp_54_ram[478] = 15;
    exp_54_ram[479] = 255;
    exp_54_ram[480] = 15;
    exp_54_ram[481] = 254;
    exp_54_ram[482] = 0;
    exp_54_ram[483] = 254;
    exp_54_ram[484] = 255;
    exp_54_ram[485] = 0;
    exp_54_ram[486] = 252;
    exp_54_ram[487] = 250;
    exp_54_ram[488] = 250;
    exp_54_ram[489] = 2;
    exp_54_ram[490] = 250;
    exp_54_ram[491] = 250;
    exp_54_ram[492] = 0;
    exp_54_ram[493] = 254;
    exp_54_ram[494] = 1;
    exp_54_ram[495] = 246;
    exp_54_ram[496] = 250;
    exp_54_ram[497] = 252;
    exp_54_ram[498] = 0;
    exp_54_ram[499] = 0;
    exp_54_ram[500] = 0;
    exp_54_ram[501] = 0;
    exp_54_ram[502] = 250;
    exp_54_ram[503] = 0;
    exp_54_ram[504] = 250;
    exp_54_ram[505] = 0;
    exp_54_ram[506] = 254;
    exp_54_ram[507] = 251;
    exp_54_ram[508] = 251;
    exp_54_ram[509] = 251;
    exp_54_ram[510] = 251;
    exp_54_ram[511] = 189;
    exp_54_ram[512] = 0;
    exp_54_ram[513] = 0;
    exp_54_ram[514] = 6;
    exp_54_ram[515] = 6;
    exp_54_ram[516] = 7;
    exp_54_ram[517] = 0;
    exp_54_ram[518] = 248;
    exp_54_ram[519] = 6;
    exp_54_ram[520] = 6;
    exp_54_ram[521] = 8;
    exp_54_ram[522] = 250;
    exp_54_ram[523] = 250;
    exp_54_ram[524] = 250;
    exp_54_ram[525] = 250;
    exp_54_ram[526] = 248;
    exp_54_ram[527] = 252;
    exp_54_ram[528] = 250;
    exp_54_ram[529] = 32;
    exp_54_ram[530] = 13;
    exp_54_ram[531] = 250;
    exp_54_ram[532] = 32;
    exp_54_ram[533] = 250;
    exp_54_ram[534] = 0;
    exp_54_ram[535] = 2;
    exp_54_ram[536] = 2;
    exp_54_ram[537] = 250;
    exp_54_ram[538] = 0;
    exp_54_ram[539] = 253;
    exp_54_ram[540] = 0;
    exp_54_ram[541] = 252;
    exp_54_ram[542] = 250;
    exp_54_ram[543] = 250;
    exp_54_ram[544] = 0;
    exp_54_ram[545] = 250;
    exp_54_ram[546] = 0;
    exp_54_ram[547] = 250;
    exp_54_ram[548] = 0;
    exp_54_ram[549] = 250;
    exp_54_ram[550] = 28;
    exp_54_ram[551] = 250;
    exp_54_ram[552] = 0;
    exp_54_ram[553] = 250;
    exp_54_ram[554] = 254;
    exp_54_ram[555] = 250;
    exp_54_ram[556] = 0;
    exp_54_ram[557] = 254;
    exp_54_ram[558] = 1;
    exp_54_ram[559] = 12;
    exp_54_ram[560] = 0;
    exp_54_ram[561] = 0;
    exp_54_ram[562] = 58;
    exp_54_ram[563] = 0;
    exp_54_ram[564] = 0;
    exp_54_ram[565] = 0;
    exp_54_ram[566] = 254;
    exp_54_ram[567] = 0;
    exp_54_ram[568] = 254;
    exp_54_ram[569] = 250;
    exp_54_ram[570] = 0;
    exp_54_ram[571] = 250;
    exp_54_ram[572] = 0;
    exp_54_ram[573] = 254;
    exp_54_ram[574] = 9;
    exp_54_ram[575] = 254;
    exp_54_ram[576] = 0;
    exp_54_ram[577] = 254;
    exp_54_ram[578] = 250;
    exp_54_ram[579] = 0;
    exp_54_ram[580] = 250;
    exp_54_ram[581] = 0;
    exp_54_ram[582] = 254;
    exp_54_ram[583] = 7;
    exp_54_ram[584] = 254;
    exp_54_ram[585] = 0;
    exp_54_ram[586] = 254;
    exp_54_ram[587] = 250;
    exp_54_ram[588] = 0;
    exp_54_ram[589] = 250;
    exp_54_ram[590] = 0;
    exp_54_ram[591] = 254;
    exp_54_ram[592] = 5;
    exp_54_ram[593] = 254;
    exp_54_ram[594] = 0;
    exp_54_ram[595] = 254;
    exp_54_ram[596] = 250;
    exp_54_ram[597] = 0;
    exp_54_ram[598] = 250;
    exp_54_ram[599] = 0;
    exp_54_ram[600] = 254;
    exp_54_ram[601] = 3;
    exp_54_ram[602] = 254;
    exp_54_ram[603] = 1;
    exp_54_ram[604] = 254;
    exp_54_ram[605] = 250;
    exp_54_ram[606] = 0;
    exp_54_ram[607] = 250;
    exp_54_ram[608] = 0;
    exp_54_ram[609] = 254;
    exp_54_ram[610] = 0;
    exp_54_ram[611] = 254;
    exp_54_ram[612] = 0;
    exp_54_ram[613] = 254;
    exp_54_ram[614] = 240;
    exp_54_ram[615] = 254;
    exp_54_ram[616] = 250;
    exp_54_ram[617] = 0;
    exp_54_ram[618] = 0;
    exp_54_ram[619] = 128;
    exp_54_ram[620] = 0;
    exp_54_ram[621] = 0;
    exp_54_ram[622] = 250;
    exp_54_ram[623] = 0;
    exp_54_ram[624] = 132;
    exp_54_ram[625] = 254;
    exp_54_ram[626] = 6;
    exp_54_ram[627] = 250;
    exp_54_ram[628] = 0;
    exp_54_ram[629] = 2;
    exp_54_ram[630] = 4;
    exp_54_ram[631] = 249;
    exp_54_ram[632] = 0;
    exp_54_ram[633] = 248;
    exp_54_ram[634] = 0;
    exp_54_ram[635] = 252;
    exp_54_ram[636] = 252;
    exp_54_ram[637] = 2;
    exp_54_ram[638] = 254;
    exp_54_ram[639] = 0;
    exp_54_ram[640] = 254;
    exp_54_ram[641] = 252;
    exp_54_ram[642] = 64;
    exp_54_ram[643] = 254;
    exp_54_ram[644] = 0;
    exp_54_ram[645] = 252;
    exp_54_ram[646] = 254;
    exp_54_ram[647] = 250;
    exp_54_ram[648] = 0;
    exp_54_ram[649] = 250;
    exp_54_ram[650] = 254;
    exp_54_ram[651] = 250;
    exp_54_ram[652] = 0;
    exp_54_ram[653] = 2;
    exp_54_ram[654] = 8;
    exp_54_ram[655] = 254;
    exp_54_ram[656] = 64;
    exp_54_ram[657] = 254;
    exp_54_ram[658] = 250;
    exp_54_ram[659] = 0;
    exp_54_ram[660] = 250;
    exp_54_ram[661] = 250;
    exp_54_ram[662] = 0;
    exp_54_ram[663] = 0;
    exp_54_ram[664] = 245;
    exp_54_ram[665] = 0;
    exp_54_ram[666] = 0;
    exp_54_ram[667] = 250;
    exp_54_ram[668] = 0;
    exp_54_ram[669] = 249;
    exp_54_ram[670] = 254;
    exp_54_ram[671] = 4;
    exp_54_ram[672] = 250;
    exp_54_ram[673] = 0;
    exp_54_ram[674] = 2;
    exp_54_ram[675] = 2;
    exp_54_ram[676] = 249;
    exp_54_ram[677] = 0;
    exp_54_ram[678] = 248;
    exp_54_ram[679] = 0;
    exp_54_ram[680] = 252;
    exp_54_ram[681] = 252;
    exp_54_ram[682] = 0;
    exp_54_ram[683] = 0;
    exp_54_ram[684] = 254;
    exp_54_ram[685] = 250;
    exp_54_ram[686] = 0;
    exp_54_ram[687] = 250;
    exp_54_ram[688] = 250;
    exp_54_ram[689] = 0;
    exp_54_ram[690] = 249;
    exp_54_ram[691] = 1;
    exp_54_ram[692] = 14;
    exp_54_ram[693] = 0;
    exp_54_ram[694] = 0;
    exp_54_ram[695] = 62;
    exp_54_ram[696] = 0;
    exp_54_ram[697] = 0;
    exp_54_ram[698] = 0;
    exp_54_ram[699] = 254;
    exp_54_ram[700] = 16;
    exp_54_ram[701] = 254;
    exp_54_ram[702] = 250;
    exp_54_ram[703] = 0;
    exp_54_ram[704] = 250;
    exp_54_ram[705] = 250;
    exp_54_ram[706] = 0;
    exp_54_ram[707] = 6;
    exp_54_ram[708] = 12;
    exp_54_ram[709] = 254;
    exp_54_ram[710] = 32;
    exp_54_ram[711] = 254;
    exp_54_ram[712] = 250;
    exp_54_ram[713] = 0;
    exp_54_ram[714] = 250;
    exp_54_ram[715] = 10;
    exp_54_ram[716] = 254;
    exp_54_ram[717] = 8;
    exp_54_ram[718] = 254;
    exp_54_ram[719] = 250;
    exp_54_ram[720] = 0;
    exp_54_ram[721] = 250;
    exp_54_ram[722] = 250;
    exp_54_ram[723] = 0;
    exp_54_ram[724] = 6;
    exp_54_ram[725] = 8;
    exp_54_ram[726] = 254;
    exp_54_ram[727] = 4;
    exp_54_ram[728] = 254;
    exp_54_ram[729] = 250;
    exp_54_ram[730] = 0;
    exp_54_ram[731] = 250;
    exp_54_ram[732] = 6;
    exp_54_ram[733] = 254;
    exp_54_ram[734] = 16;
    exp_54_ram[735] = 254;
    exp_54_ram[736] = 250;
    exp_54_ram[737] = 0;
    exp_54_ram[738] = 250;
    exp_54_ram[739] = 5;
    exp_54_ram[740] = 254;
    exp_54_ram[741] = 32;
    exp_54_ram[742] = 254;
    exp_54_ram[743] = 250;
    exp_54_ram[744] = 0;
    exp_54_ram[745] = 250;
    exp_54_ram[746] = 3;
    exp_54_ram[747] = 254;
    exp_54_ram[748] = 16;
    exp_54_ram[749] = 254;
    exp_54_ram[750] = 250;
    exp_54_ram[751] = 0;
    exp_54_ram[752] = 250;
    exp_54_ram[753] = 1;
    exp_54_ram[754] = 0;
    exp_54_ram[755] = 1;
    exp_54_ram[756] = 0;
    exp_54_ram[757] = 0;
    exp_54_ram[758] = 0;
    exp_54_ram[759] = 250;
    exp_54_ram[760] = 0;
    exp_54_ram[761] = 253;
    exp_54_ram[762] = 5;
    exp_54_ram[763] = 98;
    exp_54_ram[764] = 0;
    exp_54_ram[765] = 0;
    exp_54_ram[766] = 67;
    exp_54_ram[767] = 0;
    exp_54_ram[768] = 0;
    exp_54_ram[769] = 0;
    exp_54_ram[770] = 250;
    exp_54_ram[771] = 0;
    exp_54_ram[772] = 7;
    exp_54_ram[773] = 0;
    exp_54_ram[774] = 250;
    exp_54_ram[775] = 0;
    exp_54_ram[776] = 5;
    exp_54_ram[777] = 0;
    exp_54_ram[778] = 1;
    exp_54_ram[779] = 252;
    exp_54_ram[780] = 5;
    exp_54_ram[781] = 250;
    exp_54_ram[782] = 0;
    exp_54_ram[783] = 6;
    exp_54_ram[784] = 0;
    exp_54_ram[785] = 0;
    exp_54_ram[786] = 252;
    exp_54_ram[787] = 3;
    exp_54_ram[788] = 250;
    exp_54_ram[789] = 0;
    exp_54_ram[790] = 6;
    exp_54_ram[791] = 0;
    exp_54_ram[792] = 0;
    exp_54_ram[793] = 252;
    exp_54_ram[794] = 1;
    exp_54_ram[795] = 0;
    exp_54_ram[796] = 252;
    exp_54_ram[797] = 254;
    exp_54_ram[798] = 254;
    exp_54_ram[799] = 254;
    exp_54_ram[800] = 250;
    exp_54_ram[801] = 0;
    exp_54_ram[802] = 5;
    exp_54_ram[803] = 0;
    exp_54_ram[804] = 254;
    exp_54_ram[805] = 2;
    exp_54_ram[806] = 254;
    exp_54_ram[807] = 250;
    exp_54_ram[808] = 0;
    exp_54_ram[809] = 6;
    exp_54_ram[810] = 2;
    exp_54_ram[811] = 250;
    exp_54_ram[812] = 0;
    exp_54_ram[813] = 6;
    exp_54_ram[814] = 0;
    exp_54_ram[815] = 254;
    exp_54_ram[816] = 255;
    exp_54_ram[817] = 254;
    exp_54_ram[818] = 254;
    exp_54_ram[819] = 64;
    exp_54_ram[820] = 0;
    exp_54_ram[821] = 254;
    exp_54_ram[822] = 255;
    exp_54_ram[823] = 254;
    exp_54_ram[824] = 250;
    exp_54_ram[825] = 0;
    exp_54_ram[826] = 6;
    exp_54_ram[827] = 0;
    exp_54_ram[828] = 250;
    exp_54_ram[829] = 0;
    exp_54_ram[830] = 6;
    exp_54_ram[831] = 20;
    exp_54_ram[832] = 254;
    exp_54_ram[833] = 32;
    exp_54_ram[834] = 34;
    exp_54_ram[835] = 254;
    exp_54_ram[836] = 16;
    exp_54_ram[837] = 6;
    exp_54_ram[838] = 249;
    exp_54_ram[839] = 0;
    exp_54_ram[840] = 248;
    exp_54_ram[841] = 0;
    exp_54_ram[842] = 250;
    exp_54_ram[843] = 251;
    exp_54_ram[844] = 65;
    exp_54_ram[845] = 251;
    exp_54_ram[846] = 0;
    exp_54_ram[847] = 64;
    exp_54_ram[848] = 0;
    exp_54_ram[849] = 251;
    exp_54_ram[850] = 1;
    exp_54_ram[851] = 15;
    exp_54_ram[852] = 254;
    exp_54_ram[853] = 0;
    exp_54_ram[854] = 254;
    exp_54_ram[855] = 0;
    exp_54_ram[856] = 254;
    exp_54_ram[857] = 253;
    exp_54_ram[858] = 0;
    exp_54_ram[859] = 0;
    exp_54_ram[860] = 250;
    exp_54_ram[861] = 253;
    exp_54_ram[862] = 250;
    exp_54_ram[863] = 250;
    exp_54_ram[864] = 149;
    exp_54_ram[865] = 252;
    exp_54_ram[866] = 27;
    exp_54_ram[867] = 254;
    exp_54_ram[868] = 4;
    exp_54_ram[869] = 0;
    exp_54_ram[870] = 249;
    exp_54_ram[871] = 0;
    exp_54_ram[872] = 248;
    exp_54_ram[873] = 0;
    exp_54_ram[874] = 15;
    exp_54_ram[875] = 3;
    exp_54_ram[876] = 254;
    exp_54_ram[877] = 8;
    exp_54_ram[878] = 2;
    exp_54_ram[879] = 249;
    exp_54_ram[880] = 0;
    exp_54_ram[881] = 248;
    exp_54_ram[882] = 0;
    exp_54_ram[883] = 1;
    exp_54_ram[884] = 65;
    exp_54_ram[885] = 1;
    exp_54_ram[886] = 249;
    exp_54_ram[887] = 0;
    exp_54_ram[888] = 248;
    exp_54_ram[889] = 0;
    exp_54_ram[890] = 250;
    exp_54_ram[891] = 251;
    exp_54_ram[892] = 65;
    exp_54_ram[893] = 251;
    exp_54_ram[894] = 0;
    exp_54_ram[895] = 64;
    exp_54_ram[896] = 0;
    exp_54_ram[897] = 251;
    exp_54_ram[898] = 1;
    exp_54_ram[899] = 15;
    exp_54_ram[900] = 254;
    exp_54_ram[901] = 0;
    exp_54_ram[902] = 254;
    exp_54_ram[903] = 0;
    exp_54_ram[904] = 254;
    exp_54_ram[905] = 253;
    exp_54_ram[906] = 0;
    exp_54_ram[907] = 0;
    exp_54_ram[908] = 250;
    exp_54_ram[909] = 253;
    exp_54_ram[910] = 250;
    exp_54_ram[911] = 250;
    exp_54_ram[912] = 137;
    exp_54_ram[913] = 252;
    exp_54_ram[914] = 15;
    exp_54_ram[915] = 254;
    exp_54_ram[916] = 32;
    exp_54_ram[917] = 14;
    exp_54_ram[918] = 254;
    exp_54_ram[919] = 16;
    exp_54_ram[920] = 4;
    exp_54_ram[921] = 249;
    exp_54_ram[922] = 0;
    exp_54_ram[923] = 248;
    exp_54_ram[924] = 0;
    exp_54_ram[925] = 254;
    exp_54_ram[926] = 0;
    exp_54_ram[927] = 254;
    exp_54_ram[928] = 0;
    exp_54_ram[929] = 254;
    exp_54_ram[930] = 253;
    exp_54_ram[931] = 0;
    exp_54_ram[932] = 250;
    exp_54_ram[933] = 253;
    exp_54_ram[934] = 250;
    exp_54_ram[935] = 250;
    exp_54_ram[936] = 131;
    exp_54_ram[937] = 252;
    exp_54_ram[938] = 9;
    exp_54_ram[939] = 254;
    exp_54_ram[940] = 4;
    exp_54_ram[941] = 0;
    exp_54_ram[942] = 249;
    exp_54_ram[943] = 0;
    exp_54_ram[944] = 248;
    exp_54_ram[945] = 0;
    exp_54_ram[946] = 15;
    exp_54_ram[947] = 3;
    exp_54_ram[948] = 254;
    exp_54_ram[949] = 8;
    exp_54_ram[950] = 2;
    exp_54_ram[951] = 249;
    exp_54_ram[952] = 0;
    exp_54_ram[953] = 248;
    exp_54_ram[954] = 0;
    exp_54_ram[955] = 1;
    exp_54_ram[956] = 1;
    exp_54_ram[957] = 1;
    exp_54_ram[958] = 249;
    exp_54_ram[959] = 0;
    exp_54_ram[960] = 248;
    exp_54_ram[961] = 0;
    exp_54_ram[962] = 252;
    exp_54_ram[963] = 254;
    exp_54_ram[964] = 0;
    exp_54_ram[965] = 254;
    exp_54_ram[966] = 0;
    exp_54_ram[967] = 254;
    exp_54_ram[968] = 253;
    exp_54_ram[969] = 0;
    exp_54_ram[970] = 252;
    exp_54_ram[971] = 250;
    exp_54_ram[972] = 253;
    exp_54_ram[973] = 250;
    exp_54_ram[974] = 250;
    exp_54_ram[975] = 249;
    exp_54_ram[976] = 252;
    exp_54_ram[977] = 250;
    exp_54_ram[978] = 0;
    exp_54_ram[979] = 250;
    exp_54_ram[980] = 48;
    exp_54_ram[981] = 0;
    exp_54_ram[982] = 252;
    exp_54_ram[983] = 254;
    exp_54_ram[984] = 0;
    exp_54_ram[985] = 4;
    exp_54_ram[986] = 2;
    exp_54_ram[987] = 253;
    exp_54_ram[988] = 0;
    exp_54_ram[989] = 252;
    exp_54_ram[990] = 250;
    exp_54_ram[991] = 250;
    exp_54_ram[992] = 0;
    exp_54_ram[993] = 250;
    exp_54_ram[994] = 2;
    exp_54_ram[995] = 0;
    exp_54_ram[996] = 253;
    exp_54_ram[997] = 0;
    exp_54_ram[998] = 252;
    exp_54_ram[999] = 254;
    exp_54_ram[1000] = 252;
    exp_54_ram[1001] = 249;
    exp_54_ram[1002] = 0;
    exp_54_ram[1003] = 248;
    exp_54_ram[1004] = 0;
    exp_54_ram[1005] = 15;
    exp_54_ram[1006] = 253;
    exp_54_ram[1007] = 0;
    exp_54_ram[1008] = 252;
    exp_54_ram[1009] = 250;
    exp_54_ram[1010] = 250;
    exp_54_ram[1011] = 0;
    exp_54_ram[1012] = 250;
    exp_54_ram[1013] = 0;
    exp_54_ram[1014] = 254;
    exp_54_ram[1015] = 0;
    exp_54_ram[1016] = 4;
    exp_54_ram[1017] = 2;
    exp_54_ram[1018] = 253;
    exp_54_ram[1019] = 0;
    exp_54_ram[1020] = 252;
    exp_54_ram[1021] = 250;
    exp_54_ram[1022] = 250;
    exp_54_ram[1023] = 0;
    exp_54_ram[1024] = 250;
    exp_54_ram[1025] = 2;
    exp_54_ram[1026] = 0;
    exp_54_ram[1027] = 253;
    exp_54_ram[1028] = 0;
    exp_54_ram[1029] = 252;
    exp_54_ram[1030] = 254;
    exp_54_ram[1031] = 252;
    exp_54_ram[1032] = 250;
    exp_54_ram[1033] = 0;
    exp_54_ram[1034] = 250;
    exp_54_ram[1035] = 35;
    exp_54_ram[1036] = 249;
    exp_54_ram[1037] = 0;
    exp_54_ram[1038] = 248;
    exp_54_ram[1039] = 0;
    exp_54_ram[1040] = 252;
    exp_54_ram[1041] = 254;
    exp_54_ram[1042] = 0;
    exp_54_ram[1043] = 254;
    exp_54_ram[1044] = 0;
    exp_54_ram[1045] = 255;
    exp_54_ram[1046] = 0;
    exp_54_ram[1047] = 253;
    exp_54_ram[1048] = 143;
    exp_54_ram[1049] = 252;
    exp_54_ram[1050] = 254;
    exp_54_ram[1051] = 64;
    exp_54_ram[1052] = 0;
    exp_54_ram[1053] = 252;
    exp_54_ram[1054] = 254;
    exp_54_ram[1055] = 0;
    exp_54_ram[1056] = 0;
    exp_54_ram[1057] = 252;
    exp_54_ram[1058] = 254;
    exp_54_ram[1059] = 0;
    exp_54_ram[1060] = 6;
    exp_54_ram[1061] = 2;
    exp_54_ram[1062] = 253;
    exp_54_ram[1063] = 0;
    exp_54_ram[1064] = 252;
    exp_54_ram[1065] = 250;
    exp_54_ram[1066] = 250;
    exp_54_ram[1067] = 0;
    exp_54_ram[1068] = 250;
    exp_54_ram[1069] = 2;
    exp_54_ram[1070] = 0;
    exp_54_ram[1071] = 252;
    exp_54_ram[1072] = 0;
    exp_54_ram[1073] = 252;
    exp_54_ram[1074] = 254;
    exp_54_ram[1075] = 252;
    exp_54_ram[1076] = 3;
    exp_54_ram[1077] = 253;
    exp_54_ram[1078] = 0;
    exp_54_ram[1079] = 252;
    exp_54_ram[1080] = 0;
    exp_54_ram[1081] = 253;
    exp_54_ram[1082] = 0;
    exp_54_ram[1083] = 252;
    exp_54_ram[1084] = 250;
    exp_54_ram[1085] = 250;
    exp_54_ram[1086] = 0;
    exp_54_ram[1087] = 250;
    exp_54_ram[1088] = 0;
    exp_54_ram[1089] = 253;
    exp_54_ram[1090] = 0;
    exp_54_ram[1091] = 2;
    exp_54_ram[1092] = 254;
    exp_54_ram[1093] = 64;
    exp_54_ram[1094] = 250;
    exp_54_ram[1095] = 254;
    exp_54_ram[1096] = 255;
    exp_54_ram[1097] = 254;
    exp_54_ram[1098] = 250;
    exp_54_ram[1099] = 254;
    exp_54_ram[1100] = 0;
    exp_54_ram[1101] = 4;
    exp_54_ram[1102] = 2;
    exp_54_ram[1103] = 253;
    exp_54_ram[1104] = 0;
    exp_54_ram[1105] = 252;
    exp_54_ram[1106] = 250;
    exp_54_ram[1107] = 250;
    exp_54_ram[1108] = 0;
    exp_54_ram[1109] = 250;
    exp_54_ram[1110] = 2;
    exp_54_ram[1111] = 0;
    exp_54_ram[1112] = 252;
    exp_54_ram[1113] = 0;
    exp_54_ram[1114] = 252;
    exp_54_ram[1115] = 254;
    exp_54_ram[1116] = 252;
    exp_54_ram[1117] = 250;
    exp_54_ram[1118] = 0;
    exp_54_ram[1119] = 250;
    exp_54_ram[1120] = 13;
    exp_54_ram[1121] = 0;
    exp_54_ram[1122] = 254;
    exp_54_ram[1123] = 254;
    exp_54_ram[1124] = 2;
    exp_54_ram[1125] = 254;
    exp_54_ram[1126] = 249;
    exp_54_ram[1127] = 0;
    exp_54_ram[1128] = 248;
    exp_54_ram[1129] = 0;
    exp_54_ram[1130] = 0;
    exp_54_ram[1131] = 254;
    exp_54_ram[1132] = 0;
    exp_54_ram[1133] = 254;
    exp_54_ram[1134] = 0;
    exp_54_ram[1135] = 254;
    exp_54_ram[1136] = 1;
    exp_54_ram[1137] = 0;
    exp_54_ram[1138] = 250;
    exp_54_ram[1139] = 253;
    exp_54_ram[1140] = 250;
    exp_54_ram[1141] = 250;
    exp_54_ram[1142] = 207;
    exp_54_ram[1143] = 252;
    exp_54_ram[1144] = 250;
    exp_54_ram[1145] = 0;
    exp_54_ram[1146] = 250;
    exp_54_ram[1147] = 7;
    exp_54_ram[1148] = 253;
    exp_54_ram[1149] = 0;
    exp_54_ram[1150] = 252;
    exp_54_ram[1151] = 250;
    exp_54_ram[1152] = 250;
    exp_54_ram[1153] = 0;
    exp_54_ram[1154] = 250;
    exp_54_ram[1155] = 2;
    exp_54_ram[1156] = 0;
    exp_54_ram[1157] = 250;
    exp_54_ram[1158] = 0;
    exp_54_ram[1159] = 250;
    exp_54_ram[1160] = 3;
    exp_54_ram[1161] = 250;
    exp_54_ram[1162] = 0;
    exp_54_ram[1163] = 253;
    exp_54_ram[1164] = 0;
    exp_54_ram[1165] = 252;
    exp_54_ram[1166] = 250;
    exp_54_ram[1167] = 250;
    exp_54_ram[1168] = 0;
    exp_54_ram[1169] = 250;
    exp_54_ram[1170] = 0;
    exp_54_ram[1171] = 250;
    exp_54_ram[1172] = 0;
    exp_54_ram[1173] = 250;
    exp_54_ram[1174] = 0;
    exp_54_ram[1175] = 250;
    exp_54_ram[1176] = 0;
    exp_54_ram[1177] = 222;
    exp_54_ram[1178] = 253;
    exp_54_ram[1179] = 250;
    exp_54_ram[1180] = 0;
    exp_54_ram[1181] = 250;
    exp_54_ram[1182] = 255;
    exp_54_ram[1183] = 0;
    exp_54_ram[1184] = 253;
    exp_54_ram[1185] = 250;
    exp_54_ram[1186] = 250;
    exp_54_ram[1187] = 0;
    exp_54_ram[1188] = 250;
    exp_54_ram[1189] = 0;
    exp_54_ram[1190] = 0;
    exp_54_ram[1191] = 253;
    exp_54_ram[1192] = 0;
    exp_54_ram[1193] = 7;
    exp_54_ram[1194] = 7;
    exp_54_ram[1195] = 8;
    exp_54_ram[1196] = 0;
    exp_54_ram[1197] = 251;
    exp_54_ram[1198] = 2;
    exp_54_ram[1199] = 2;
    exp_54_ram[1200] = 3;
    exp_54_ram[1201] = 252;
    exp_54_ram[1202] = 0;
    exp_54_ram[1203] = 0;
    exp_54_ram[1204] = 0;
    exp_54_ram[1205] = 0;
    exp_54_ram[1206] = 0;
    exp_54_ram[1207] = 1;
    exp_54_ram[1208] = 1;
    exp_54_ram[1209] = 2;
    exp_54_ram[1210] = 252;
    exp_54_ram[1211] = 253;
    exp_54_ram[1212] = 254;
    exp_54_ram[1213] = 254;
    exp_54_ram[1214] = 254;
    exp_54_ram[1215] = 254;
    exp_54_ram[1216] = 253;
    exp_54_ram[1217] = 255;
    exp_54_ram[1218] = 0;
    exp_54_ram[1219] = 16;
    exp_54_ram[1220] = 208;
    exp_54_ram[1221] = 254;
    exp_54_ram[1222] = 254;
    exp_54_ram[1223] = 0;
    exp_54_ram[1224] = 2;
    exp_54_ram[1225] = 2;
    exp_54_ram[1226] = 5;
    exp_54_ram[1227] = 0;
    exp_54_ram[1228] = 254;
    exp_54_ram[1229] = 0;
    exp_54_ram[1230] = 0;
    exp_54_ram[1231] = 2;
    exp_54_ram[1232] = 0;
    exp_54_ram[1233] = 254;
    exp_54_ram[1234] = 254;
    exp_54_ram[1235] = 0;
    exp_54_ram[1236] = 58;
    exp_54_ram[1237] = 0;
    exp_54_ram[1238] = 0;
    exp_54_ram[1239] = 212;
    exp_54_ram[1240] = 0;
    exp_54_ram[1241] = 1;
    exp_54_ram[1242] = 1;
    exp_54_ram[1243] = 2;
    exp_54_ram[1244] = 0;
    exp_54_ram[1245] = 255;
    exp_54_ram[1246] = 0;
    exp_54_ram[1247] = 0;
    exp_54_ram[1248] = 1;
    exp_54_ram[1249] = 8;
    exp_54_ram[1250] = 242;
    exp_54_ram[1251] = 0;
    exp_54_ram[1252] = 0;
    exp_54_ram[1253] = 0;
    exp_54_ram[1254] = 1;
    exp_54_ram[1255] = 0;
    exp_54_ram[1256] = 128;
    exp_54_ram[1257] = 0;
    exp_54_ram[1258] = 0;
    exp_54_ram[1259] = 0;
    exp_54_ram[1260] = 0;
    exp_54_ram[1261] = 0;
    exp_54_ram[1262] = 0;
    exp_54_ram[1263] = 0;
    exp_54_ram[1264] = 0;
    exp_54_ram[1265] = 0;
    exp_54_ram[1266] = 0;
    exp_54_ram[1267] = 0;
    exp_54_ram[1268] = 0;
    exp_54_ram[1269] = 0;
    exp_54_ram[1270] = 0;
    exp_54_ram[1271] = 0;
    exp_54_ram[1272] = 0;
    exp_54_ram[1273] = 0;
    exp_54_ram[1274] = 0;
    exp_54_ram[1275] = 0;
    exp_54_ram[1276] = 0;
    exp_54_ram[1277] = 0;
    exp_54_ram[1278] = 0;
    exp_54_ram[1279] = 0;
    exp_54_ram[1280] = 0;
    exp_54_ram[1281] = 0;
    exp_54_ram[1282] = 0;
    exp_54_ram[1283] = 0;
    exp_54_ram[1284] = 0;
    exp_54_ram[1285] = 0;
    exp_54_ram[1286] = 0;
    exp_54_ram[1287] = 0;
    exp_54_ram[1288] = 0;
    exp_54_ram[1289] = 0;
    exp_54_ram[1290] = 0;
    exp_54_ram[1291] = 0;
    exp_54_ram[1292] = 0;
    exp_54_ram[1293] = 0;
    exp_54_ram[1294] = 0;
    exp_54_ram[1295] = 0;
    exp_54_ram[1296] = 0;
    exp_54_ram[1297] = 0;
    exp_54_ram[1298] = 0;
    exp_54_ram[1299] = 0;
    exp_54_ram[1300] = 0;
    exp_54_ram[1301] = 0;
    exp_54_ram[1302] = 0;
    exp_54_ram[1303] = 0;
    exp_54_ram[1304] = 0;
    exp_54_ram[1305] = 0;
    exp_54_ram[1306] = 0;
    exp_54_ram[1307] = 0;
    exp_54_ram[1308] = 0;
    exp_54_ram[1309] = 0;
    exp_54_ram[1310] = 0;
    exp_54_ram[1311] = 0;
    exp_54_ram[1312] = 0;
    exp_54_ram[1313] = 0;
    exp_54_ram[1314] = 0;
    exp_54_ram[1315] = 0;
    exp_54_ram[1316] = 0;
    exp_54_ram[1317] = 0;
    exp_54_ram[1318] = 0;
    exp_54_ram[1319] = 0;
    exp_54_ram[1320] = 0;
    exp_54_ram[1321] = 0;
    exp_54_ram[1322] = 0;
    exp_54_ram[1323] = 0;
    exp_54_ram[1324] = 0;
    exp_54_ram[1325] = 0;
    exp_54_ram[1326] = 0;
    exp_54_ram[1327] = 0;
    exp_54_ram[1328] = 0;
    exp_54_ram[1329] = 0;
    exp_54_ram[1330] = 0;
    exp_54_ram[1331] = 0;
    exp_54_ram[1332] = 0;
    exp_54_ram[1333] = 0;
    exp_54_ram[1334] = 0;
    exp_54_ram[1335] = 0;
    exp_54_ram[1336] = 0;
    exp_54_ram[1337] = 0;
    exp_54_ram[1338] = 0;
    exp_54_ram[1339] = 0;
    exp_54_ram[1340] = 0;
    exp_54_ram[1341] = 0;
    exp_54_ram[1342] = 0;
    exp_54_ram[1343] = 0;
    exp_54_ram[1344] = 0;
    exp_54_ram[1345] = 0;
    exp_54_ram[1346] = 0;
    exp_54_ram[1347] = 0;
    exp_54_ram[1348] = 0;
    exp_54_ram[1349] = 0;
    exp_54_ram[1350] = 0;
    exp_54_ram[1351] = 0;
    exp_54_ram[1352] = 0;
    exp_54_ram[1353] = 0;
    exp_54_ram[1354] = 0;
    exp_54_ram[1355] = 0;
    exp_54_ram[1356] = 0;
    exp_54_ram[1357] = 0;
    exp_54_ram[1358] = 0;
    exp_54_ram[1359] = 0;
    exp_54_ram[1360] = 0;
    exp_54_ram[1361] = 0;
    exp_54_ram[1362] = 0;
    exp_54_ram[1363] = 0;
    exp_54_ram[1364] = 0;
    exp_54_ram[1365] = 0;
    exp_54_ram[1366] = 0;
    exp_54_ram[1367] = 0;
    exp_54_ram[1368] = 0;
    exp_54_ram[1369] = 0;
    exp_54_ram[1370] = 0;
    exp_54_ram[1371] = 0;
    exp_54_ram[1372] = 0;
    exp_54_ram[1373] = 0;
    exp_54_ram[1374] = 0;
    exp_54_ram[1375] = 0;
    exp_54_ram[1376] = 0;
    exp_54_ram[1377] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_230;
  assign exp_230 = exp_511;

  reg [3:0] exp_511_reg;
  always@(*) begin
    case (exp_363)
      0:exp_511_reg <= exp_498;
      1:exp_511_reg <= exp_503;
      2:exp_511_reg <= exp_504;
      3:exp_511_reg <= exp_505;
      4:exp_511_reg <= exp_506;
      5:exp_511_reg <= exp_507;
      6:exp_511_reg <= exp_508;
      7:exp_511_reg <= exp_509;
      default:exp_511_reg <= exp_510;
    endcase
  end
  assign exp_511 = exp_511_reg;
  assign exp_510 = 0;
  assign exp_498 = exp_494 << exp_497;
  assign exp_494 = 1;
  assign exp_497 = exp_496 + exp_495;
  assign exp_496 = 0;
  assign exp_495 = exp_431[1:0];
  assign exp_503 = exp_499 << exp_502;
  assign exp_499 = 3;
  assign exp_502 = exp_501 + exp_500;
  assign exp_501 = 0;
  assign exp_500 = exp_431[1:1];
  assign exp_504 = 15;
  assign exp_505 = 0;
  assign exp_506 = 0;
  assign exp_507 = 0;
  assign exp_508 = 0;
  assign exp_509 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_225;
  assign exp_225 = exp_493;

  reg [31:0] exp_493_reg;
  always@(*) begin
    case (exp_363)
      0:exp_493_reg <= exp_480;
      1:exp_493_reg <= exp_484;
      2:exp_493_reg <= exp_486;
      3:exp_493_reg <= exp_487;
      4:exp_493_reg <= exp_488;
      5:exp_493_reg <= exp_489;
      6:exp_493_reg <= exp_490;
      7:exp_493_reg <= exp_491;
      default:exp_493_reg <= exp_492;
    endcase
  end
  assign exp_493 = exp_493_reg;
  assign exp_492 = 0;

  reg [31:0] exp_480_reg;
  always@(*) begin
    case (exp_434)
      0:exp_480_reg <= exp_466;
      1:exp_480_reg <= exp_474;
      2:exp_480_reg <= exp_476;
      3:exp_480_reg <= exp_478;
      default:exp_480_reg <= exp_479;
    endcase
  end
  assign exp_480 = exp_480_reg;
  assign exp_479 = 0;
  assign exp_466 = exp_465;
  assign exp_465 = exp_464 + exp_463;
  assign exp_464 = 0;
  assign exp_463 = exp_353[7:0];

      reg [31:0] exp_353_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_353_reg <= exp_296;
        end
      end
      assign exp_353 = exp_353_reg;
      assign exp_474 = exp_466 << exp_473;
  assign exp_473 = 8;
  assign exp_476 = exp_466 << exp_475;
  assign exp_475 = 16;
  assign exp_478 = exp_466 << exp_477;
  assign exp_477 = 24;

  reg [31:0] exp_484_reg;
  always@(*) begin
    case (exp_437)
      0:exp_484_reg <= exp_470;
      1:exp_484_reg <= exp_482;
      default:exp_484_reg <= exp_483;
    endcase
  end
  assign exp_484 = exp_484_reg;
  assign exp_437 = exp_436 + exp_435;
  assign exp_436 = 0;
  assign exp_435 = exp_431[1:1];
  assign exp_483 = 0;
  assign exp_470 = exp_469;
  assign exp_469 = exp_468 + exp_467;
  assign exp_468 = 0;
  assign exp_467 = exp_353[15:0];
  assign exp_482 = exp_470 << exp_481;
  assign exp_481 = 16;
  assign exp_486 = exp_485 + exp_472;
  assign exp_485 = 0;
  assign exp_472 = exp_471 + exp_353;
  assign exp_471 = 0;
  assign exp_487 = 0;
  assign exp_488 = 0;
  assign exp_489 = 0;
  assign exp_490 = 0;
  assign exp_491 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 0;
    exp_47_ram[32] = 1;
    exp_47_ram[33] = 0;
    exp_47_ram[34] = 0;
    exp_47_ram[35] = 108;
    exp_47_ram[36] = 87;
    exp_47_ram[37] = 100;
    exp_47_ram[38] = 0;
    exp_47_ram[39] = 1;
    exp_47_ram[40] = 129;
    exp_47_ram[41] = 1;
    exp_47_ram[42] = 164;
    exp_47_ram[43] = 180;
    exp_47_ram[44] = 132;
    exp_47_ram[45] = 244;
    exp_47_ram[46] = 196;
    exp_47_ram[47] = 196;
    exp_47_ram[48] = 231;
    exp_47_ram[49] = 196;
    exp_47_ram[50] = 7;
    exp_47_ram[51] = 193;
    exp_47_ram[52] = 1;
    exp_47_ram[53] = 0;
    exp_47_ram[54] = 1;
    exp_47_ram[55] = 129;
    exp_47_ram[56] = 1;
    exp_47_ram[57] = 5;
    exp_47_ram[58] = 180;
    exp_47_ram[59] = 196;
    exp_47_ram[60] = 212;
    exp_47_ram[61] = 244;
    exp_47_ram[62] = 0;
    exp_47_ram[63] = 193;
    exp_47_ram[64] = 1;
    exp_47_ram[65] = 0;
    exp_47_ram[66] = 1;
    exp_47_ram[67] = 17;
    exp_47_ram[68] = 129;
    exp_47_ram[69] = 1;
    exp_47_ram[70] = 5;
    exp_47_ram[71] = 180;
    exp_47_ram[72] = 196;
    exp_47_ram[73] = 212;
    exp_47_ram[74] = 244;
    exp_47_ram[75] = 244;
    exp_47_ram[76] = 7;
    exp_47_ram[77] = 244;
    exp_47_ram[78] = 7;
    exp_47_ram[79] = 64;
    exp_47_ram[80] = 0;
    exp_47_ram[81] = 193;
    exp_47_ram[82] = 129;
    exp_47_ram[83] = 1;
    exp_47_ram[84] = 0;
    exp_47_ram[85] = 1;
    exp_47_ram[86] = 129;
    exp_47_ram[87] = 1;
    exp_47_ram[88] = 164;
    exp_47_ram[89] = 180;
    exp_47_ram[90] = 196;
    exp_47_ram[91] = 244;
    exp_47_ram[92] = 0;
    exp_47_ram[93] = 196;
    exp_47_ram[94] = 23;
    exp_47_ram[95] = 244;
    exp_47_ram[96] = 196;
    exp_47_ram[97] = 7;
    exp_47_ram[98] = 7;
    exp_47_ram[99] = 132;
    exp_47_ram[100] = 247;
    exp_47_ram[101] = 228;
    exp_47_ram[102] = 7;
    exp_47_ram[103] = 196;
    exp_47_ram[104] = 196;
    exp_47_ram[105] = 247;
    exp_47_ram[106] = 7;
    exp_47_ram[107] = 193;
    exp_47_ram[108] = 1;
    exp_47_ram[109] = 0;
    exp_47_ram[110] = 1;
    exp_47_ram[111] = 129;
    exp_47_ram[112] = 1;
    exp_47_ram[113] = 5;
    exp_47_ram[114] = 244;
    exp_47_ram[115] = 244;
    exp_47_ram[116] = 240;
    exp_47_ram[117] = 231;
    exp_47_ram[118] = 244;
    exp_47_ram[119] = 144;
    exp_47_ram[120] = 231;
    exp_47_ram[121] = 16;
    exp_47_ram[122] = 128;
    exp_47_ram[123] = 0;
    exp_47_ram[124] = 23;
    exp_47_ram[125] = 247;
    exp_47_ram[126] = 7;
    exp_47_ram[127] = 193;
    exp_47_ram[128] = 1;
    exp_47_ram[129] = 0;
    exp_47_ram[130] = 1;
    exp_47_ram[131] = 17;
    exp_47_ram[132] = 129;
    exp_47_ram[133] = 1;
    exp_47_ram[134] = 164;
    exp_47_ram[135] = 4;
    exp_47_ram[136] = 0;
    exp_47_ram[137] = 196;
    exp_47_ram[138] = 7;
    exp_47_ram[139] = 39;
    exp_47_ram[140] = 231;
    exp_47_ram[141] = 23;
    exp_47_ram[142] = 7;
    exp_47_ram[143] = 196;
    exp_47_ram[144] = 7;
    exp_47_ram[145] = 23;
    exp_47_ram[146] = 196;
    exp_47_ram[147] = 215;
    exp_47_ram[148] = 7;
    exp_47_ram[149] = 246;
    exp_47_ram[150] = 7;
    exp_47_ram[151] = 244;
    exp_47_ram[152] = 196;
    exp_47_ram[153] = 7;
    exp_47_ram[154] = 7;
    exp_47_ram[155] = 7;
    exp_47_ram[156] = 159;
    exp_47_ram[157] = 5;
    exp_47_ram[158] = 7;
    exp_47_ram[159] = 196;
    exp_47_ram[160] = 7;
    exp_47_ram[161] = 193;
    exp_47_ram[162] = 129;
    exp_47_ram[163] = 1;
    exp_47_ram[164] = 0;
    exp_47_ram[165] = 1;
    exp_47_ram[166] = 17;
    exp_47_ram[167] = 129;
    exp_47_ram[168] = 1;
    exp_47_ram[169] = 164;
    exp_47_ram[170] = 180;
    exp_47_ram[171] = 196;
    exp_47_ram[172] = 212;
    exp_47_ram[173] = 228;
    exp_47_ram[174] = 244;
    exp_47_ram[175] = 4;
    exp_47_ram[176] = 20;
    exp_47_ram[177] = 68;
    exp_47_ram[178] = 244;
    exp_47_ram[179] = 4;
    exp_47_ram[180] = 39;
    exp_47_ram[181] = 7;
    exp_47_ram[182] = 4;
    exp_47_ram[183] = 23;
    exp_47_ram[184] = 7;
    exp_47_ram[185] = 132;
    exp_47_ram[186] = 244;
    exp_47_ram[187] = 64;
    exp_47_ram[188] = 68;
    exp_47_ram[189] = 23;
    exp_47_ram[190] = 228;
    exp_47_ram[191] = 196;
    exp_47_ram[192] = 4;
    exp_47_ram[193] = 7;
    exp_47_ram[194] = 132;
    exp_47_ram[195] = 0;
    exp_47_ram[196] = 7;
    exp_47_ram[197] = 196;
    exp_47_ram[198] = 23;
    exp_47_ram[199] = 244;
    exp_47_ram[200] = 196;
    exp_47_ram[201] = 68;
    exp_47_ram[202] = 247;
    exp_47_ram[203] = 0;
    exp_47_ram[204] = 132;
    exp_47_ram[205] = 247;
    exp_47_ram[206] = 244;
    exp_47_ram[207] = 196;
    exp_47_ram[208] = 132;
    exp_47_ram[209] = 247;
    exp_47_ram[210] = 7;
    exp_47_ram[211] = 68;
    exp_47_ram[212] = 23;
    exp_47_ram[213] = 228;
    exp_47_ram[214] = 196;
    exp_47_ram[215] = 4;
    exp_47_ram[216] = 7;
    exp_47_ram[217] = 132;
    exp_47_ram[218] = 7;
    exp_47_ram[219] = 132;
    exp_47_ram[220] = 7;
    exp_47_ram[221] = 4;
    exp_47_ram[222] = 39;
    exp_47_ram[223] = 7;
    exp_47_ram[224] = 128;
    exp_47_ram[225] = 68;
    exp_47_ram[226] = 23;
    exp_47_ram[227] = 228;
    exp_47_ram[228] = 196;
    exp_47_ram[229] = 4;
    exp_47_ram[230] = 7;
    exp_47_ram[231] = 132;
    exp_47_ram[232] = 0;
    exp_47_ram[233] = 7;
    exp_47_ram[234] = 68;
    exp_47_ram[235] = 132;
    exp_47_ram[236] = 247;
    exp_47_ram[237] = 68;
    exp_47_ram[238] = 231;
    exp_47_ram[239] = 68;
    exp_47_ram[240] = 7;
    exp_47_ram[241] = 193;
    exp_47_ram[242] = 129;
    exp_47_ram[243] = 1;
    exp_47_ram[244] = 0;
    exp_47_ram[245] = 1;
    exp_47_ram[246] = 17;
    exp_47_ram[247] = 129;
    exp_47_ram[248] = 1;
    exp_47_ram[249] = 164;
    exp_47_ram[250] = 180;
    exp_47_ram[251] = 196;
    exp_47_ram[252] = 212;
    exp_47_ram[253] = 228;
    exp_47_ram[254] = 244;
    exp_47_ram[255] = 8;
    exp_47_ram[256] = 20;
    exp_47_ram[257] = 244;
    exp_47_ram[258] = 132;
    exp_47_ram[259] = 39;
    exp_47_ram[260] = 7;
    exp_47_ram[261] = 68;
    exp_47_ram[262] = 7;
    exp_47_ram[263] = 132;
    exp_47_ram[264] = 23;
    exp_47_ram[265] = 7;
    exp_47_ram[266] = 116;
    exp_47_ram[267] = 7;
    exp_47_ram[268] = 132;
    exp_47_ram[269] = 199;
    exp_47_ram[270] = 7;
    exp_47_ram[271] = 68;
    exp_47_ram[272] = 247;
    exp_47_ram[273] = 244;
    exp_47_ram[274] = 0;
    exp_47_ram[275] = 132;
    exp_47_ram[276] = 23;
    exp_47_ram[277] = 228;
    exp_47_ram[278] = 196;
    exp_47_ram[279] = 247;
    exp_47_ram[280] = 0;
    exp_47_ram[281] = 231;
    exp_47_ram[282] = 132;
    exp_47_ram[283] = 4;
    exp_47_ram[284] = 247;
    exp_47_ram[285] = 132;
    exp_47_ram[286] = 240;
    exp_47_ram[287] = 231;
    exp_47_ram[288] = 0;
    exp_47_ram[289] = 132;
    exp_47_ram[290] = 23;
    exp_47_ram[291] = 228;
    exp_47_ram[292] = 196;
    exp_47_ram[293] = 247;
    exp_47_ram[294] = 0;
    exp_47_ram[295] = 231;
    exp_47_ram[296] = 132;
    exp_47_ram[297] = 23;
    exp_47_ram[298] = 7;
    exp_47_ram[299] = 132;
    exp_47_ram[300] = 68;
    exp_47_ram[301] = 247;
    exp_47_ram[302] = 132;
    exp_47_ram[303] = 240;
    exp_47_ram[304] = 231;
    exp_47_ram[305] = 132;
    exp_47_ram[306] = 7;
    exp_47_ram[307] = 7;
    exp_47_ram[308] = 132;
    exp_47_ram[309] = 7;
    exp_47_ram[310] = 7;
    exp_47_ram[311] = 132;
    exp_47_ram[312] = 7;
    exp_47_ram[313] = 132;
    exp_47_ram[314] = 4;
    exp_47_ram[315] = 247;
    exp_47_ram[316] = 132;
    exp_47_ram[317] = 68;
    exp_47_ram[318] = 247;
    exp_47_ram[319] = 132;
    exp_47_ram[320] = 247;
    exp_47_ram[321] = 244;
    exp_47_ram[322] = 132;
    exp_47_ram[323] = 7;
    exp_47_ram[324] = 4;
    exp_47_ram[325] = 0;
    exp_47_ram[326] = 247;
    exp_47_ram[327] = 132;
    exp_47_ram[328] = 247;
    exp_47_ram[329] = 244;
    exp_47_ram[330] = 4;
    exp_47_ram[331] = 0;
    exp_47_ram[332] = 247;
    exp_47_ram[333] = 132;
    exp_47_ram[334] = 7;
    exp_47_ram[335] = 7;
    exp_47_ram[336] = 132;
    exp_47_ram[337] = 240;
    exp_47_ram[338] = 231;
    exp_47_ram[339] = 132;
    exp_47_ram[340] = 23;
    exp_47_ram[341] = 228;
    exp_47_ram[342] = 196;
    exp_47_ram[343] = 247;
    exp_47_ram[344] = 128;
    exp_47_ram[345] = 231;
    exp_47_ram[346] = 192;
    exp_47_ram[347] = 4;
    exp_47_ram[348] = 0;
    exp_47_ram[349] = 247;
    exp_47_ram[350] = 132;
    exp_47_ram[351] = 7;
    exp_47_ram[352] = 7;
    exp_47_ram[353] = 132;
    exp_47_ram[354] = 240;
    exp_47_ram[355] = 231;
    exp_47_ram[356] = 132;
    exp_47_ram[357] = 23;
    exp_47_ram[358] = 228;
    exp_47_ram[359] = 196;
    exp_47_ram[360] = 247;
    exp_47_ram[361] = 128;
    exp_47_ram[362] = 231;
    exp_47_ram[363] = 128;
    exp_47_ram[364] = 4;
    exp_47_ram[365] = 32;
    exp_47_ram[366] = 247;
    exp_47_ram[367] = 132;
    exp_47_ram[368] = 240;
    exp_47_ram[369] = 231;
    exp_47_ram[370] = 132;
    exp_47_ram[371] = 23;
    exp_47_ram[372] = 228;
    exp_47_ram[373] = 196;
    exp_47_ram[374] = 247;
    exp_47_ram[375] = 32;
    exp_47_ram[376] = 231;
    exp_47_ram[377] = 132;
    exp_47_ram[378] = 240;
    exp_47_ram[379] = 231;
    exp_47_ram[380] = 132;
    exp_47_ram[381] = 23;
    exp_47_ram[382] = 228;
    exp_47_ram[383] = 196;
    exp_47_ram[384] = 247;
    exp_47_ram[385] = 0;
    exp_47_ram[386] = 231;
    exp_47_ram[387] = 132;
    exp_47_ram[388] = 240;
    exp_47_ram[389] = 231;
    exp_47_ram[390] = 116;
    exp_47_ram[391] = 7;
    exp_47_ram[392] = 132;
    exp_47_ram[393] = 23;
    exp_47_ram[394] = 228;
    exp_47_ram[395] = 196;
    exp_47_ram[396] = 247;
    exp_47_ram[397] = 208;
    exp_47_ram[398] = 231;
    exp_47_ram[399] = 128;
    exp_47_ram[400] = 132;
    exp_47_ram[401] = 71;
    exp_47_ram[402] = 7;
    exp_47_ram[403] = 132;
    exp_47_ram[404] = 23;
    exp_47_ram[405] = 228;
    exp_47_ram[406] = 196;
    exp_47_ram[407] = 247;
    exp_47_ram[408] = 176;
    exp_47_ram[409] = 231;
    exp_47_ram[410] = 192;
    exp_47_ram[411] = 132;
    exp_47_ram[412] = 135;
    exp_47_ram[413] = 7;
    exp_47_ram[414] = 132;
    exp_47_ram[415] = 23;
    exp_47_ram[416] = 228;
    exp_47_ram[417] = 196;
    exp_47_ram[418] = 247;
    exp_47_ram[419] = 0;
    exp_47_ram[420] = 231;
    exp_47_ram[421] = 132;
    exp_47_ram[422] = 68;
    exp_47_ram[423] = 132;
    exp_47_ram[424] = 196;
    exp_47_ram[425] = 4;
    exp_47_ram[426] = 68;
    exp_47_ram[427] = 132;
    exp_47_ram[428] = 196;
    exp_47_ram[429] = 31;
    exp_47_ram[430] = 5;
    exp_47_ram[431] = 7;
    exp_47_ram[432] = 193;
    exp_47_ram[433] = 129;
    exp_47_ram[434] = 1;
    exp_47_ram[435] = 0;
    exp_47_ram[436] = 1;
    exp_47_ram[437] = 17;
    exp_47_ram[438] = 129;
    exp_47_ram[439] = 1;
    exp_47_ram[440] = 164;
    exp_47_ram[441] = 180;
    exp_47_ram[442] = 196;
    exp_47_ram[443] = 212;
    exp_47_ram[444] = 228;
    exp_47_ram[445] = 4;
    exp_47_ram[446] = 20;
    exp_47_ram[447] = 244;
    exp_47_ram[448] = 4;
    exp_47_ram[449] = 196;
    exp_47_ram[450] = 7;
    exp_47_ram[451] = 68;
    exp_47_ram[452] = 247;
    exp_47_ram[453] = 244;
    exp_47_ram[454] = 68;
    exp_47_ram[455] = 7;
    exp_47_ram[456] = 7;
    exp_47_ram[457] = 196;
    exp_47_ram[458] = 7;
    exp_47_ram[459] = 196;
    exp_47_ram[460] = 68;
    exp_47_ram[461] = 247;
    exp_47_ram[462] = 244;
    exp_47_ram[463] = 180;
    exp_47_ram[464] = 144;
    exp_47_ram[465] = 231;
    exp_47_ram[466] = 180;
    exp_47_ram[467] = 7;
    exp_47_ram[468] = 247;
    exp_47_ram[469] = 0;
    exp_47_ram[470] = 68;
    exp_47_ram[471] = 7;
    exp_47_ram[472] = 7;
    exp_47_ram[473] = 16;
    exp_47_ram[474] = 128;
    exp_47_ram[475] = 16;
    exp_47_ram[476] = 180;
    exp_47_ram[477] = 231;
    exp_47_ram[478] = 247;
    exp_47_ram[479] = 103;
    exp_47_ram[480] = 247;
    exp_47_ram[481] = 196;
    exp_47_ram[482] = 23;
    exp_47_ram[483] = 212;
    exp_47_ram[484] = 4;
    exp_47_ram[485] = 230;
    exp_47_ram[486] = 247;
    exp_47_ram[487] = 196;
    exp_47_ram[488] = 68;
    exp_47_ram[489] = 247;
    exp_47_ram[490] = 244;
    exp_47_ram[491] = 196;
    exp_47_ram[492] = 7;
    exp_47_ram[493] = 196;
    exp_47_ram[494] = 240;
    exp_47_ram[495] = 231;
    exp_47_ram[496] = 180;
    exp_47_ram[497] = 132;
    exp_47_ram[498] = 68;
    exp_47_ram[499] = 241;
    exp_47_ram[500] = 4;
    exp_47_ram[501] = 241;
    exp_47_ram[502] = 4;
    exp_47_ram[503] = 241;
    exp_47_ram[504] = 68;
    exp_47_ram[505] = 6;
    exp_47_ram[506] = 196;
    exp_47_ram[507] = 4;
    exp_47_ram[508] = 68;
    exp_47_ram[509] = 132;
    exp_47_ram[510] = 196;
    exp_47_ram[511] = 159;
    exp_47_ram[512] = 5;
    exp_47_ram[513] = 7;
    exp_47_ram[514] = 193;
    exp_47_ram[515] = 129;
    exp_47_ram[516] = 1;
    exp_47_ram[517] = 0;
    exp_47_ram[518] = 1;
    exp_47_ram[519] = 17;
    exp_47_ram[520] = 129;
    exp_47_ram[521] = 1;
    exp_47_ram[522] = 164;
    exp_47_ram[523] = 180;
    exp_47_ram[524] = 196;
    exp_47_ram[525] = 212;
    exp_47_ram[526] = 228;
    exp_47_ram[527] = 4;
    exp_47_ram[528] = 132;
    exp_47_ram[529] = 7;
    exp_47_ram[530] = 128;
    exp_47_ram[531] = 244;
    exp_47_ram[532] = 208;
    exp_47_ram[533] = 4;
    exp_47_ram[534] = 7;
    exp_47_ram[535] = 80;
    exp_47_ram[536] = 247;
    exp_47_ram[537] = 4;
    exp_47_ram[538] = 7;
    exp_47_ram[539] = 196;
    exp_47_ram[540] = 23;
    exp_47_ram[541] = 228;
    exp_47_ram[542] = 196;
    exp_47_ram[543] = 68;
    exp_47_ram[544] = 7;
    exp_47_ram[545] = 132;
    exp_47_ram[546] = 7;
    exp_47_ram[547] = 4;
    exp_47_ram[548] = 23;
    exp_47_ram[549] = 244;
    exp_47_ram[550] = 80;
    exp_47_ram[551] = 4;
    exp_47_ram[552] = 23;
    exp_47_ram[553] = 244;
    exp_47_ram[554] = 4;
    exp_47_ram[555] = 4;
    exp_47_ram[556] = 7;
    exp_47_ram[557] = 7;
    exp_47_ram[558] = 0;
    exp_47_ram[559] = 247;
    exp_47_ram[560] = 39;
    exp_47_ram[561] = 0;
    exp_47_ram[562] = 71;
    exp_47_ram[563] = 247;
    exp_47_ram[564] = 7;
    exp_47_ram[565] = 7;
    exp_47_ram[566] = 196;
    exp_47_ram[567] = 23;
    exp_47_ram[568] = 244;
    exp_47_ram[569] = 4;
    exp_47_ram[570] = 23;
    exp_47_ram[571] = 244;
    exp_47_ram[572] = 16;
    exp_47_ram[573] = 244;
    exp_47_ram[574] = 192;
    exp_47_ram[575] = 196;
    exp_47_ram[576] = 39;
    exp_47_ram[577] = 244;
    exp_47_ram[578] = 4;
    exp_47_ram[579] = 23;
    exp_47_ram[580] = 244;
    exp_47_ram[581] = 16;
    exp_47_ram[582] = 244;
    exp_47_ram[583] = 128;
    exp_47_ram[584] = 196;
    exp_47_ram[585] = 71;
    exp_47_ram[586] = 244;
    exp_47_ram[587] = 4;
    exp_47_ram[588] = 23;
    exp_47_ram[589] = 244;
    exp_47_ram[590] = 16;
    exp_47_ram[591] = 244;
    exp_47_ram[592] = 64;
    exp_47_ram[593] = 196;
    exp_47_ram[594] = 135;
    exp_47_ram[595] = 244;
    exp_47_ram[596] = 4;
    exp_47_ram[597] = 23;
    exp_47_ram[598] = 244;
    exp_47_ram[599] = 16;
    exp_47_ram[600] = 244;
    exp_47_ram[601] = 0;
    exp_47_ram[602] = 196;
    exp_47_ram[603] = 7;
    exp_47_ram[604] = 244;
    exp_47_ram[605] = 4;
    exp_47_ram[606] = 23;
    exp_47_ram[607] = 244;
    exp_47_ram[608] = 16;
    exp_47_ram[609] = 244;
    exp_47_ram[610] = 192;
    exp_47_ram[611] = 4;
    exp_47_ram[612] = 0;
    exp_47_ram[613] = 4;
    exp_47_ram[614] = 7;
    exp_47_ram[615] = 4;
    exp_47_ram[616] = 4;
    exp_47_ram[617] = 7;
    exp_47_ram[618] = 7;
    exp_47_ram[619] = 223;
    exp_47_ram[620] = 5;
    exp_47_ram[621] = 7;
    exp_47_ram[622] = 4;
    exp_47_ram[623] = 7;
    exp_47_ram[624] = 159;
    exp_47_ram[625] = 164;
    exp_47_ram[626] = 0;
    exp_47_ram[627] = 4;
    exp_47_ram[628] = 7;
    exp_47_ram[629] = 160;
    exp_47_ram[630] = 247;
    exp_47_ram[631] = 196;
    exp_47_ram[632] = 71;
    exp_47_ram[633] = 228;
    exp_47_ram[634] = 7;
    exp_47_ram[635] = 244;
    exp_47_ram[636] = 132;
    exp_47_ram[637] = 7;
    exp_47_ram[638] = 196;
    exp_47_ram[639] = 39;
    exp_47_ram[640] = 244;
    exp_47_ram[641] = 132;
    exp_47_ram[642] = 240;
    exp_47_ram[643] = 244;
    exp_47_ram[644] = 192;
    exp_47_ram[645] = 132;
    exp_47_ram[646] = 244;
    exp_47_ram[647] = 4;
    exp_47_ram[648] = 23;
    exp_47_ram[649] = 244;
    exp_47_ram[650] = 4;
    exp_47_ram[651] = 4;
    exp_47_ram[652] = 7;
    exp_47_ram[653] = 224;
    exp_47_ram[654] = 247;
    exp_47_ram[655] = 196;
    exp_47_ram[656] = 7;
    exp_47_ram[657] = 244;
    exp_47_ram[658] = 4;
    exp_47_ram[659] = 23;
    exp_47_ram[660] = 244;
    exp_47_ram[661] = 4;
    exp_47_ram[662] = 7;
    exp_47_ram[663] = 7;
    exp_47_ram[664] = 143;
    exp_47_ram[665] = 5;
    exp_47_ram[666] = 7;
    exp_47_ram[667] = 4;
    exp_47_ram[668] = 7;
    exp_47_ram[669] = 79;
    exp_47_ram[670] = 164;
    exp_47_ram[671] = 64;
    exp_47_ram[672] = 4;
    exp_47_ram[673] = 7;
    exp_47_ram[674] = 160;
    exp_47_ram[675] = 247;
    exp_47_ram[676] = 196;
    exp_47_ram[677] = 71;
    exp_47_ram[678] = 228;
    exp_47_ram[679] = 7;
    exp_47_ram[680] = 244;
    exp_47_ram[681] = 68;
    exp_47_ram[682] = 7;
    exp_47_ram[683] = 0;
    exp_47_ram[684] = 244;
    exp_47_ram[685] = 4;
    exp_47_ram[686] = 23;
    exp_47_ram[687] = 244;
    exp_47_ram[688] = 4;
    exp_47_ram[689] = 7;
    exp_47_ram[690] = 135;
    exp_47_ram[691] = 32;
    exp_47_ram[692] = 247;
    exp_47_ram[693] = 39;
    exp_47_ram[694] = 0;
    exp_47_ram[695] = 135;
    exp_47_ram[696] = 247;
    exp_47_ram[697] = 7;
    exp_47_ram[698] = 7;
    exp_47_ram[699] = 196;
    exp_47_ram[700] = 7;
    exp_47_ram[701] = 244;
    exp_47_ram[702] = 4;
    exp_47_ram[703] = 23;
    exp_47_ram[704] = 244;
    exp_47_ram[705] = 4;
    exp_47_ram[706] = 7;
    exp_47_ram[707] = 192;
    exp_47_ram[708] = 247;
    exp_47_ram[709] = 196;
    exp_47_ram[710] = 7;
    exp_47_ram[711] = 244;
    exp_47_ram[712] = 4;
    exp_47_ram[713] = 23;
    exp_47_ram[714] = 244;
    exp_47_ram[715] = 64;
    exp_47_ram[716] = 196;
    exp_47_ram[717] = 7;
    exp_47_ram[718] = 244;
    exp_47_ram[719] = 4;
    exp_47_ram[720] = 23;
    exp_47_ram[721] = 244;
    exp_47_ram[722] = 4;
    exp_47_ram[723] = 7;
    exp_47_ram[724] = 128;
    exp_47_ram[725] = 247;
    exp_47_ram[726] = 196;
    exp_47_ram[727] = 7;
    exp_47_ram[728] = 244;
    exp_47_ram[729] = 4;
    exp_47_ram[730] = 23;
    exp_47_ram[731] = 244;
    exp_47_ram[732] = 128;
    exp_47_ram[733] = 196;
    exp_47_ram[734] = 7;
    exp_47_ram[735] = 244;
    exp_47_ram[736] = 4;
    exp_47_ram[737] = 23;
    exp_47_ram[738] = 244;
    exp_47_ram[739] = 0;
    exp_47_ram[740] = 196;
    exp_47_ram[741] = 7;
    exp_47_ram[742] = 244;
    exp_47_ram[743] = 4;
    exp_47_ram[744] = 23;
    exp_47_ram[745] = 244;
    exp_47_ram[746] = 64;
    exp_47_ram[747] = 196;
    exp_47_ram[748] = 7;
    exp_47_ram[749] = 244;
    exp_47_ram[750] = 4;
    exp_47_ram[751] = 23;
    exp_47_ram[752] = 244;
    exp_47_ram[753] = 128;
    exp_47_ram[754] = 0;
    exp_47_ram[755] = 0;
    exp_47_ram[756] = 0;
    exp_47_ram[757] = 128;
    exp_47_ram[758] = 0;
    exp_47_ram[759] = 4;
    exp_47_ram[760] = 7;
    exp_47_ram[761] = 183;
    exp_47_ram[762] = 48;
    exp_47_ram[763] = 247;
    exp_47_ram[764] = 39;
    exp_47_ram[765] = 0;
    exp_47_ram[766] = 71;
    exp_47_ram[767] = 247;
    exp_47_ram[768] = 7;
    exp_47_ram[769] = 7;
    exp_47_ram[770] = 4;
    exp_47_ram[771] = 7;
    exp_47_ram[772] = 128;
    exp_47_ram[773] = 247;
    exp_47_ram[774] = 4;
    exp_47_ram[775] = 7;
    exp_47_ram[776] = 128;
    exp_47_ram[777] = 247;
    exp_47_ram[778] = 0;
    exp_47_ram[779] = 244;
    exp_47_ram[780] = 0;
    exp_47_ram[781] = 4;
    exp_47_ram[782] = 7;
    exp_47_ram[783] = 240;
    exp_47_ram[784] = 247;
    exp_47_ram[785] = 128;
    exp_47_ram[786] = 244;
    exp_47_ram[787] = 64;
    exp_47_ram[788] = 4;
    exp_47_ram[789] = 7;
    exp_47_ram[790] = 32;
    exp_47_ram[791] = 247;
    exp_47_ram[792] = 32;
    exp_47_ram[793] = 244;
    exp_47_ram[794] = 128;
    exp_47_ram[795] = 160;
    exp_47_ram[796] = 244;
    exp_47_ram[797] = 196;
    exp_47_ram[798] = 247;
    exp_47_ram[799] = 244;
    exp_47_ram[800] = 4;
    exp_47_ram[801] = 7;
    exp_47_ram[802] = 128;
    exp_47_ram[803] = 247;
    exp_47_ram[804] = 196;
    exp_47_ram[805] = 7;
    exp_47_ram[806] = 244;
    exp_47_ram[807] = 4;
    exp_47_ram[808] = 7;
    exp_47_ram[809] = 144;
    exp_47_ram[810] = 247;
    exp_47_ram[811] = 4;
    exp_47_ram[812] = 7;
    exp_47_ram[813] = 64;
    exp_47_ram[814] = 247;
    exp_47_ram[815] = 196;
    exp_47_ram[816] = 55;
    exp_47_ram[817] = 244;
    exp_47_ram[818] = 196;
    exp_47_ram[819] = 7;
    exp_47_ram[820] = 7;
    exp_47_ram[821] = 196;
    exp_47_ram[822] = 231;
    exp_47_ram[823] = 244;
    exp_47_ram[824] = 4;
    exp_47_ram[825] = 7;
    exp_47_ram[826] = 144;
    exp_47_ram[827] = 247;
    exp_47_ram[828] = 4;
    exp_47_ram[829] = 7;
    exp_47_ram[830] = 64;
    exp_47_ram[831] = 247;
    exp_47_ram[832] = 196;
    exp_47_ram[833] = 7;
    exp_47_ram[834] = 7;
    exp_47_ram[835] = 196;
    exp_47_ram[836] = 7;
    exp_47_ram[837] = 7;
    exp_47_ram[838] = 196;
    exp_47_ram[839] = 71;
    exp_47_ram[840] = 228;
    exp_47_ram[841] = 7;
    exp_47_ram[842] = 244;
    exp_47_ram[843] = 132;
    exp_47_ram[844] = 247;
    exp_47_ram[845] = 132;
    exp_47_ram[846] = 247;
    exp_47_ram[847] = 231;
    exp_47_ram[848] = 7;
    exp_47_ram[849] = 132;
    exp_47_ram[850] = 247;
    exp_47_ram[851] = 247;
    exp_47_ram[852] = 196;
    exp_47_ram[853] = 241;
    exp_47_ram[854] = 132;
    exp_47_ram[855] = 241;
    exp_47_ram[856] = 68;
    exp_47_ram[857] = 132;
    exp_47_ram[858] = 7;
    exp_47_ram[859] = 6;
    exp_47_ram[860] = 68;
    exp_47_ram[861] = 196;
    exp_47_ram[862] = 132;
    exp_47_ram[863] = 196;
    exp_47_ram[864] = 31;
    exp_47_ram[865] = 164;
    exp_47_ram[866] = 192;
    exp_47_ram[867] = 196;
    exp_47_ram[868] = 7;
    exp_47_ram[869] = 7;
    exp_47_ram[870] = 196;
    exp_47_ram[871] = 71;
    exp_47_ram[872] = 228;
    exp_47_ram[873] = 7;
    exp_47_ram[874] = 247;
    exp_47_ram[875] = 192;
    exp_47_ram[876] = 196;
    exp_47_ram[877] = 7;
    exp_47_ram[878] = 7;
    exp_47_ram[879] = 196;
    exp_47_ram[880] = 71;
    exp_47_ram[881] = 228;
    exp_47_ram[882] = 7;
    exp_47_ram[883] = 7;
    exp_47_ram[884] = 7;
    exp_47_ram[885] = 64;
    exp_47_ram[886] = 196;
    exp_47_ram[887] = 71;
    exp_47_ram[888] = 228;
    exp_47_ram[889] = 7;
    exp_47_ram[890] = 244;
    exp_47_ram[891] = 196;
    exp_47_ram[892] = 247;
    exp_47_ram[893] = 196;
    exp_47_ram[894] = 247;
    exp_47_ram[895] = 231;
    exp_47_ram[896] = 7;
    exp_47_ram[897] = 196;
    exp_47_ram[898] = 247;
    exp_47_ram[899] = 247;
    exp_47_ram[900] = 196;
    exp_47_ram[901] = 241;
    exp_47_ram[902] = 132;
    exp_47_ram[903] = 241;
    exp_47_ram[904] = 68;
    exp_47_ram[905] = 132;
    exp_47_ram[906] = 7;
    exp_47_ram[907] = 6;
    exp_47_ram[908] = 68;
    exp_47_ram[909] = 196;
    exp_47_ram[910] = 132;
    exp_47_ram[911] = 196;
    exp_47_ram[912] = 31;
    exp_47_ram[913] = 164;
    exp_47_ram[914] = 192;
    exp_47_ram[915] = 196;
    exp_47_ram[916] = 7;
    exp_47_ram[917] = 7;
    exp_47_ram[918] = 196;
    exp_47_ram[919] = 7;
    exp_47_ram[920] = 7;
    exp_47_ram[921] = 196;
    exp_47_ram[922] = 71;
    exp_47_ram[923] = 228;
    exp_47_ram[924] = 7;
    exp_47_ram[925] = 196;
    exp_47_ram[926] = 241;
    exp_47_ram[927] = 132;
    exp_47_ram[928] = 241;
    exp_47_ram[929] = 68;
    exp_47_ram[930] = 132;
    exp_47_ram[931] = 0;
    exp_47_ram[932] = 68;
    exp_47_ram[933] = 196;
    exp_47_ram[934] = 132;
    exp_47_ram[935] = 196;
    exp_47_ram[936] = 31;
    exp_47_ram[937] = 164;
    exp_47_ram[938] = 192;
    exp_47_ram[939] = 196;
    exp_47_ram[940] = 7;
    exp_47_ram[941] = 7;
    exp_47_ram[942] = 196;
    exp_47_ram[943] = 71;
    exp_47_ram[944] = 228;
    exp_47_ram[945] = 7;
    exp_47_ram[946] = 247;
    exp_47_ram[947] = 192;
    exp_47_ram[948] = 196;
    exp_47_ram[949] = 7;
    exp_47_ram[950] = 7;
    exp_47_ram[951] = 196;
    exp_47_ram[952] = 71;
    exp_47_ram[953] = 228;
    exp_47_ram[954] = 7;
    exp_47_ram[955] = 7;
    exp_47_ram[956] = 7;
    exp_47_ram[957] = 64;
    exp_47_ram[958] = 196;
    exp_47_ram[959] = 71;
    exp_47_ram[960] = 228;
    exp_47_ram[961] = 7;
    exp_47_ram[962] = 244;
    exp_47_ram[963] = 196;
    exp_47_ram[964] = 241;
    exp_47_ram[965] = 132;
    exp_47_ram[966] = 241;
    exp_47_ram[967] = 68;
    exp_47_ram[968] = 132;
    exp_47_ram[969] = 0;
    exp_47_ram[970] = 4;
    exp_47_ram[971] = 68;
    exp_47_ram[972] = 196;
    exp_47_ram[973] = 132;
    exp_47_ram[974] = 196;
    exp_47_ram[975] = 79;
    exp_47_ram[976] = 164;
    exp_47_ram[977] = 4;
    exp_47_ram[978] = 23;
    exp_47_ram[979] = 244;
    exp_47_ram[980] = 192;
    exp_47_ram[981] = 16;
    exp_47_ram[982] = 244;
    exp_47_ram[983] = 196;
    exp_47_ram[984] = 39;
    exp_47_ram[985] = 7;
    exp_47_ram[986] = 128;
    exp_47_ram[987] = 196;
    exp_47_ram[988] = 23;
    exp_47_ram[989] = 228;
    exp_47_ram[990] = 196;
    exp_47_ram[991] = 68;
    exp_47_ram[992] = 7;
    exp_47_ram[993] = 132;
    exp_47_ram[994] = 0;
    exp_47_ram[995] = 7;
    exp_47_ram[996] = 68;
    exp_47_ram[997] = 23;
    exp_47_ram[998] = 228;
    exp_47_ram[999] = 132;
    exp_47_ram[1000] = 231;
    exp_47_ram[1001] = 196;
    exp_47_ram[1002] = 71;
    exp_47_ram[1003] = 228;
    exp_47_ram[1004] = 7;
    exp_47_ram[1005] = 247;
    exp_47_ram[1006] = 196;
    exp_47_ram[1007] = 23;
    exp_47_ram[1008] = 228;
    exp_47_ram[1009] = 196;
    exp_47_ram[1010] = 68;
    exp_47_ram[1011] = 7;
    exp_47_ram[1012] = 132;
    exp_47_ram[1013] = 7;
    exp_47_ram[1014] = 196;
    exp_47_ram[1015] = 39;
    exp_47_ram[1016] = 7;
    exp_47_ram[1017] = 128;
    exp_47_ram[1018] = 196;
    exp_47_ram[1019] = 23;
    exp_47_ram[1020] = 228;
    exp_47_ram[1021] = 196;
    exp_47_ram[1022] = 68;
    exp_47_ram[1023] = 7;
    exp_47_ram[1024] = 132;
    exp_47_ram[1025] = 0;
    exp_47_ram[1026] = 7;
    exp_47_ram[1027] = 68;
    exp_47_ram[1028] = 23;
    exp_47_ram[1029] = 228;
    exp_47_ram[1030] = 132;
    exp_47_ram[1031] = 231;
    exp_47_ram[1032] = 4;
    exp_47_ram[1033] = 23;
    exp_47_ram[1034] = 244;
    exp_47_ram[1035] = 0;
    exp_47_ram[1036] = 196;
    exp_47_ram[1037] = 71;
    exp_47_ram[1038] = 228;
    exp_47_ram[1039] = 7;
    exp_47_ram[1040] = 244;
    exp_47_ram[1041] = 68;
    exp_47_ram[1042] = 7;
    exp_47_ram[1043] = 68;
    exp_47_ram[1044] = 128;
    exp_47_ram[1045] = 240;
    exp_47_ram[1046] = 7;
    exp_47_ram[1047] = 4;
    exp_47_ram[1048] = 79;
    exp_47_ram[1049] = 164;
    exp_47_ram[1050] = 196;
    exp_47_ram[1051] = 7;
    exp_47_ram[1052] = 7;
    exp_47_ram[1053] = 196;
    exp_47_ram[1054] = 68;
    exp_47_ram[1055] = 247;
    exp_47_ram[1056] = 7;
    exp_47_ram[1057] = 244;
    exp_47_ram[1058] = 196;
    exp_47_ram[1059] = 39;
    exp_47_ram[1060] = 7;
    exp_47_ram[1061] = 128;
    exp_47_ram[1062] = 196;
    exp_47_ram[1063] = 23;
    exp_47_ram[1064] = 228;
    exp_47_ram[1065] = 196;
    exp_47_ram[1066] = 68;
    exp_47_ram[1067] = 7;
    exp_47_ram[1068] = 132;
    exp_47_ram[1069] = 0;
    exp_47_ram[1070] = 7;
    exp_47_ram[1071] = 196;
    exp_47_ram[1072] = 23;
    exp_47_ram[1073] = 228;
    exp_47_ram[1074] = 132;
    exp_47_ram[1075] = 231;
    exp_47_ram[1076] = 64;
    exp_47_ram[1077] = 4;
    exp_47_ram[1078] = 23;
    exp_47_ram[1079] = 228;
    exp_47_ram[1080] = 7;
    exp_47_ram[1081] = 196;
    exp_47_ram[1082] = 23;
    exp_47_ram[1083] = 228;
    exp_47_ram[1084] = 196;
    exp_47_ram[1085] = 68;
    exp_47_ram[1086] = 7;
    exp_47_ram[1087] = 132;
    exp_47_ram[1088] = 7;
    exp_47_ram[1089] = 4;
    exp_47_ram[1090] = 7;
    exp_47_ram[1091] = 7;
    exp_47_ram[1092] = 196;
    exp_47_ram[1093] = 7;
    exp_47_ram[1094] = 7;
    exp_47_ram[1095] = 68;
    exp_47_ram[1096] = 247;
    exp_47_ram[1097] = 228;
    exp_47_ram[1098] = 7;
    exp_47_ram[1099] = 196;
    exp_47_ram[1100] = 39;
    exp_47_ram[1101] = 7;
    exp_47_ram[1102] = 128;
    exp_47_ram[1103] = 196;
    exp_47_ram[1104] = 23;
    exp_47_ram[1105] = 228;
    exp_47_ram[1106] = 196;
    exp_47_ram[1107] = 68;
    exp_47_ram[1108] = 7;
    exp_47_ram[1109] = 132;
    exp_47_ram[1110] = 0;
    exp_47_ram[1111] = 7;
    exp_47_ram[1112] = 196;
    exp_47_ram[1113] = 23;
    exp_47_ram[1114] = 228;
    exp_47_ram[1115] = 132;
    exp_47_ram[1116] = 231;
    exp_47_ram[1117] = 4;
    exp_47_ram[1118] = 23;
    exp_47_ram[1119] = 244;
    exp_47_ram[1120] = 192;
    exp_47_ram[1121] = 128;
    exp_47_ram[1122] = 244;
    exp_47_ram[1123] = 196;
    exp_47_ram[1124] = 23;
    exp_47_ram[1125] = 244;
    exp_47_ram[1126] = 196;
    exp_47_ram[1127] = 71;
    exp_47_ram[1128] = 228;
    exp_47_ram[1129] = 7;
    exp_47_ram[1130] = 7;
    exp_47_ram[1131] = 196;
    exp_47_ram[1132] = 241;
    exp_47_ram[1133] = 132;
    exp_47_ram[1134] = 241;
    exp_47_ram[1135] = 68;
    exp_47_ram[1136] = 0;
    exp_47_ram[1137] = 0;
    exp_47_ram[1138] = 68;
    exp_47_ram[1139] = 196;
    exp_47_ram[1140] = 132;
    exp_47_ram[1141] = 196;
    exp_47_ram[1142] = 143;
    exp_47_ram[1143] = 164;
    exp_47_ram[1144] = 4;
    exp_47_ram[1145] = 23;
    exp_47_ram[1146] = 244;
    exp_47_ram[1147] = 0;
    exp_47_ram[1148] = 196;
    exp_47_ram[1149] = 23;
    exp_47_ram[1150] = 228;
    exp_47_ram[1151] = 196;
    exp_47_ram[1152] = 68;
    exp_47_ram[1153] = 7;
    exp_47_ram[1154] = 132;
    exp_47_ram[1155] = 80;
    exp_47_ram[1156] = 7;
    exp_47_ram[1157] = 4;
    exp_47_ram[1158] = 23;
    exp_47_ram[1159] = 244;
    exp_47_ram[1160] = 192;
    exp_47_ram[1161] = 4;
    exp_47_ram[1162] = 7;
    exp_47_ram[1163] = 196;
    exp_47_ram[1164] = 23;
    exp_47_ram[1165] = 228;
    exp_47_ram[1166] = 196;
    exp_47_ram[1167] = 68;
    exp_47_ram[1168] = 7;
    exp_47_ram[1169] = 132;
    exp_47_ram[1170] = 7;
    exp_47_ram[1171] = 4;
    exp_47_ram[1172] = 23;
    exp_47_ram[1173] = 244;
    exp_47_ram[1174] = 0;
    exp_47_ram[1175] = 4;
    exp_47_ram[1176] = 7;
    exp_47_ram[1177] = 7;
    exp_47_ram[1178] = 196;
    exp_47_ram[1179] = 68;
    exp_47_ram[1180] = 247;
    exp_47_ram[1181] = 68;
    exp_47_ram[1182] = 247;
    exp_47_ram[1183] = 128;
    exp_47_ram[1184] = 196;
    exp_47_ram[1185] = 196;
    exp_47_ram[1186] = 68;
    exp_47_ram[1187] = 7;
    exp_47_ram[1188] = 132;
    exp_47_ram[1189] = 0;
    exp_47_ram[1190] = 7;
    exp_47_ram[1191] = 196;
    exp_47_ram[1192] = 7;
    exp_47_ram[1193] = 193;
    exp_47_ram[1194] = 129;
    exp_47_ram[1195] = 1;
    exp_47_ram[1196] = 0;
    exp_47_ram[1197] = 1;
    exp_47_ram[1198] = 17;
    exp_47_ram[1199] = 129;
    exp_47_ram[1200] = 1;
    exp_47_ram[1201] = 164;
    exp_47_ram[1202] = 180;
    exp_47_ram[1203] = 196;
    exp_47_ram[1204] = 212;
    exp_47_ram[1205] = 228;
    exp_47_ram[1206] = 244;
    exp_47_ram[1207] = 4;
    exp_47_ram[1208] = 20;
    exp_47_ram[1209] = 4;
    exp_47_ram[1210] = 244;
    exp_47_ram[1211] = 132;
    exp_47_ram[1212] = 71;
    exp_47_ram[1213] = 244;
    exp_47_ram[1214] = 132;
    exp_47_ram[1215] = 68;
    exp_47_ram[1216] = 196;
    exp_47_ram[1217] = 240;
    exp_47_ram[1218] = 7;
    exp_47_ram[1219] = 128;
    exp_47_ram[1220] = 143;
    exp_47_ram[1221] = 164;
    exp_47_ram[1222] = 196;
    exp_47_ram[1223] = 7;
    exp_47_ram[1224] = 193;
    exp_47_ram[1225] = 129;
    exp_47_ram[1226] = 1;
    exp_47_ram[1227] = 0;
    exp_47_ram[1228] = 1;
    exp_47_ram[1229] = 17;
    exp_47_ram[1230] = 129;
    exp_47_ram[1231] = 1;
    exp_47_ram[1232] = 5;
    exp_47_ram[1233] = 244;
    exp_47_ram[1234] = 244;
    exp_47_ram[1235] = 0;
    exp_47_ram[1236] = 7;
    exp_47_ram[1237] = 7;
    exp_47_ram[1238] = 7;
    exp_47_ram[1239] = 31;
    exp_47_ram[1240] = 0;
    exp_47_ram[1241] = 193;
    exp_47_ram[1242] = 129;
    exp_47_ram[1243] = 1;
    exp_47_ram[1244] = 0;
    exp_47_ram[1245] = 1;
    exp_47_ram[1246] = 17;
    exp_47_ram[1247] = 129;
    exp_47_ram[1248] = 1;
    exp_47_ram[1249] = 192;
    exp_47_ram[1250] = 223;
    exp_47_ram[1251] = 0;
    exp_47_ram[1252] = 193;
    exp_47_ram[1253] = 129;
    exp_47_ram[1254] = 1;
    exp_47_ram[1255] = 0;
    exp_47_ram[1256] = 0;
    exp_47_ram[1257] = 0;
    exp_47_ram[1258] = 0;
    exp_47_ram[1259] = 0;
    exp_47_ram[1260] = 0;
    exp_47_ram[1261] = 0;
    exp_47_ram[1262] = 0;
    exp_47_ram[1263] = 0;
    exp_47_ram[1264] = 0;
    exp_47_ram[1265] = 0;
    exp_47_ram[1266] = 0;
    exp_47_ram[1267] = 0;
    exp_47_ram[1268] = 0;
    exp_47_ram[1269] = 0;
    exp_47_ram[1270] = 0;
    exp_47_ram[1271] = 0;
    exp_47_ram[1272] = 0;
    exp_47_ram[1273] = 0;
    exp_47_ram[1274] = 0;
    exp_47_ram[1275] = 0;
    exp_47_ram[1276] = 0;
    exp_47_ram[1277] = 0;
    exp_47_ram[1278] = 0;
    exp_47_ram[1279] = 0;
    exp_47_ram[1280] = 0;
    exp_47_ram[1281] = 0;
    exp_47_ram[1282] = 0;
    exp_47_ram[1283] = 0;
    exp_47_ram[1284] = 0;
    exp_47_ram[1285] = 0;
    exp_47_ram[1286] = 0;
    exp_47_ram[1287] = 0;
    exp_47_ram[1288] = 0;
    exp_47_ram[1289] = 0;
    exp_47_ram[1290] = 0;
    exp_47_ram[1291] = 0;
    exp_47_ram[1292] = 0;
    exp_47_ram[1293] = 0;
    exp_47_ram[1294] = 0;
    exp_47_ram[1295] = 0;
    exp_47_ram[1296] = 0;
    exp_47_ram[1297] = 0;
    exp_47_ram[1298] = 0;
    exp_47_ram[1299] = 0;
    exp_47_ram[1300] = 0;
    exp_47_ram[1301] = 0;
    exp_47_ram[1302] = 0;
    exp_47_ram[1303] = 0;
    exp_47_ram[1304] = 0;
    exp_47_ram[1305] = 0;
    exp_47_ram[1306] = 0;
    exp_47_ram[1307] = 0;
    exp_47_ram[1308] = 0;
    exp_47_ram[1309] = 0;
    exp_47_ram[1310] = 0;
    exp_47_ram[1311] = 0;
    exp_47_ram[1312] = 0;
    exp_47_ram[1313] = 0;
    exp_47_ram[1314] = 0;
    exp_47_ram[1315] = 0;
    exp_47_ram[1316] = 0;
    exp_47_ram[1317] = 0;
    exp_47_ram[1318] = 0;
    exp_47_ram[1319] = 0;
    exp_47_ram[1320] = 0;
    exp_47_ram[1321] = 0;
    exp_47_ram[1322] = 0;
    exp_47_ram[1323] = 0;
    exp_47_ram[1324] = 0;
    exp_47_ram[1325] = 0;
    exp_47_ram[1326] = 0;
    exp_47_ram[1327] = 0;
    exp_47_ram[1328] = 0;
    exp_47_ram[1329] = 0;
    exp_47_ram[1330] = 0;
    exp_47_ram[1331] = 0;
    exp_47_ram[1332] = 0;
    exp_47_ram[1333] = 0;
    exp_47_ram[1334] = 0;
    exp_47_ram[1335] = 0;
    exp_47_ram[1336] = 0;
    exp_47_ram[1337] = 0;
    exp_47_ram[1338] = 0;
    exp_47_ram[1339] = 0;
    exp_47_ram[1340] = 0;
    exp_47_ram[1341] = 0;
    exp_47_ram[1342] = 0;
    exp_47_ram[1343] = 0;
    exp_47_ram[1344] = 0;
    exp_47_ram[1345] = 0;
    exp_47_ram[1346] = 0;
    exp_47_ram[1347] = 0;
    exp_47_ram[1348] = 0;
    exp_47_ram[1349] = 0;
    exp_47_ram[1350] = 0;
    exp_47_ram[1351] = 0;
    exp_47_ram[1352] = 0;
    exp_47_ram[1353] = 0;
    exp_47_ram[1354] = 0;
    exp_47_ram[1355] = 0;
    exp_47_ram[1356] = 0;
    exp_47_ram[1357] = 0;
    exp_47_ram[1358] = 0;
    exp_47_ram[1359] = 0;
    exp_47_ram[1360] = 0;
    exp_47_ram[1361] = 0;
    exp_47_ram[1362] = 0;
    exp_47_ram[1363] = 0;
    exp_47_ram[1364] = 0;
    exp_47_ram[1365] = 0;
    exp_47_ram[1366] = 0;
    exp_47_ram[1367] = 0;
    exp_47_ram[1368] = 0;
    exp_47_ram[1369] = 0;
    exp_47_ram[1370] = 0;
    exp_47_ram[1371] = 0;
    exp_47_ram[1372] = 0;
    exp_47_ram[1373] = 0;
    exp_47_ram[1374] = 0;
    exp_47_ram[1375] = 0;
    exp_47_ram[1376] = 0;
    exp_47_ram[1377] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 33;
    exp_40_ram[32] = 1;
    exp_40_ram[33] = 16;
    exp_40_ram[34] = 0;
    exp_40_ram[35] = 101;
    exp_40_ram[36] = 32;
    exp_40_ram[37] = 108;
    exp_40_ram[38] = 0;
    exp_40_ram[39] = 1;
    exp_40_ram[40] = 38;
    exp_40_ram[41] = 4;
    exp_40_ram[42] = 46;
    exp_40_ram[43] = 44;
    exp_40_ram[44] = 39;
    exp_40_ram[45] = 38;
    exp_40_ram[46] = 39;
    exp_40_ram[47] = 39;
    exp_40_ram[48] = 160;
    exp_40_ram[49] = 39;
    exp_40_ram[50] = 133;
    exp_40_ram[51] = 36;
    exp_40_ram[52] = 1;
    exp_40_ram[53] = 128;
    exp_40_ram[54] = 1;
    exp_40_ram[55] = 46;
    exp_40_ram[56] = 4;
    exp_40_ram[57] = 7;
    exp_40_ram[58] = 36;
    exp_40_ram[59] = 34;
    exp_40_ram[60] = 32;
    exp_40_ram[61] = 7;
    exp_40_ram[62] = 0;
    exp_40_ram[63] = 36;
    exp_40_ram[64] = 1;
    exp_40_ram[65] = 128;
    exp_40_ram[66] = 1;
    exp_40_ram[67] = 46;
    exp_40_ram[68] = 44;
    exp_40_ram[69] = 4;
    exp_40_ram[70] = 7;
    exp_40_ram[71] = 36;
    exp_40_ram[72] = 34;
    exp_40_ram[73] = 32;
    exp_40_ram[74] = 7;
    exp_40_ram[75] = 71;
    exp_40_ram[76] = 136;
    exp_40_ram[77] = 71;
    exp_40_ram[78] = 133;
    exp_40_ram[79] = 16;
    exp_40_ram[80] = 0;
    exp_40_ram[81] = 32;
    exp_40_ram[82] = 36;
    exp_40_ram[83] = 1;
    exp_40_ram[84] = 128;
    exp_40_ram[85] = 1;
    exp_40_ram[86] = 38;
    exp_40_ram[87] = 4;
    exp_40_ram[88] = 46;
    exp_40_ram[89] = 44;
    exp_40_ram[90] = 39;
    exp_40_ram[91] = 38;
    exp_40_ram[92] = 0;
    exp_40_ram[93] = 39;
    exp_40_ram[94] = 135;
    exp_40_ram[95] = 38;
    exp_40_ram[96] = 39;
    exp_40_ram[97] = 199;
    exp_40_ram[98] = 138;
    exp_40_ram[99] = 39;
    exp_40_ram[100] = 135;
    exp_40_ram[101] = 44;
    exp_40_ram[102] = 158;
    exp_40_ram[103] = 39;
    exp_40_ram[104] = 39;
    exp_40_ram[105] = 7;
    exp_40_ram[106] = 133;
    exp_40_ram[107] = 36;
    exp_40_ram[108] = 1;
    exp_40_ram[109] = 128;
    exp_40_ram[110] = 1;
    exp_40_ram[111] = 46;
    exp_40_ram[112] = 4;
    exp_40_ram[113] = 7;
    exp_40_ram[114] = 7;
    exp_40_ram[115] = 71;
    exp_40_ram[116] = 7;
    exp_40_ram[117] = 252;
    exp_40_ram[118] = 71;
    exp_40_ram[119] = 7;
    exp_40_ram[120] = 230;
    exp_40_ram[121] = 7;
    exp_40_ram[122] = 0;
    exp_40_ram[123] = 7;
    exp_40_ram[124] = 247;
    exp_40_ram[125] = 247;
    exp_40_ram[126] = 133;
    exp_40_ram[127] = 36;
    exp_40_ram[128] = 1;
    exp_40_ram[129] = 128;
    exp_40_ram[130] = 1;
    exp_40_ram[131] = 38;
    exp_40_ram[132] = 36;
    exp_40_ram[133] = 4;
    exp_40_ram[134] = 46;
    exp_40_ram[135] = 38;
    exp_40_ram[136] = 0;
    exp_40_ram[137] = 39;
    exp_40_ram[138] = 7;
    exp_40_ram[139] = 151;
    exp_40_ram[140] = 135;
    exp_40_ram[141] = 151;
    exp_40_ram[142] = 134;
    exp_40_ram[143] = 39;
    exp_40_ram[144] = 167;
    exp_40_ram[145] = 134;
    exp_40_ram[146] = 39;
    exp_40_ram[147] = 32;
    exp_40_ram[148] = 199;
    exp_40_ram[149] = 7;
    exp_40_ram[150] = 135;
    exp_40_ram[151] = 38;
    exp_40_ram[152] = 39;
    exp_40_ram[153] = 167;
    exp_40_ram[154] = 199;
    exp_40_ram[155] = 133;
    exp_40_ram[156] = 240;
    exp_40_ram[157] = 7;
    exp_40_ram[158] = 150;
    exp_40_ram[159] = 39;
    exp_40_ram[160] = 133;
    exp_40_ram[161] = 32;
    exp_40_ram[162] = 36;
    exp_40_ram[163] = 1;
    exp_40_ram[164] = 128;
    exp_40_ram[165] = 1;
    exp_40_ram[166] = 46;
    exp_40_ram[167] = 44;
    exp_40_ram[168] = 4;
    exp_40_ram[169] = 46;
    exp_40_ram[170] = 44;
    exp_40_ram[171] = 42;
    exp_40_ram[172] = 40;
    exp_40_ram[173] = 38;
    exp_40_ram[174] = 36;
    exp_40_ram[175] = 34;
    exp_40_ram[176] = 32;
    exp_40_ram[177] = 39;
    exp_40_ram[178] = 36;
    exp_40_ram[179] = 39;
    exp_40_ram[180] = 247;
    exp_40_ram[181] = 156;
    exp_40_ram[182] = 39;
    exp_40_ram[183] = 247;
    exp_40_ram[184] = 150;
    exp_40_ram[185] = 39;
    exp_40_ram[186] = 38;
    exp_40_ram[187] = 0;
    exp_40_ram[188] = 39;
    exp_40_ram[189] = 135;
    exp_40_ram[190] = 42;
    exp_40_ram[191] = 39;
    exp_40_ram[192] = 38;
    exp_40_ram[193] = 134;
    exp_40_ram[194] = 37;
    exp_40_ram[195] = 5;
    exp_40_ram[196] = 0;
    exp_40_ram[197] = 39;
    exp_40_ram[198] = 135;
    exp_40_ram[199] = 38;
    exp_40_ram[200] = 39;
    exp_40_ram[201] = 39;
    exp_40_ram[202] = 100;
    exp_40_ram[203] = 0;
    exp_40_ram[204] = 39;
    exp_40_ram[205] = 135;
    exp_40_ram[206] = 36;
    exp_40_ram[207] = 39;
    exp_40_ram[208] = 39;
    exp_40_ram[209] = 7;
    exp_40_ram[210] = 197;
    exp_40_ram[211] = 39;
    exp_40_ram[212] = 135;
    exp_40_ram[213] = 42;
    exp_40_ram[214] = 39;
    exp_40_ram[215] = 38;
    exp_40_ram[216] = 134;
    exp_40_ram[217] = 37;
    exp_40_ram[218] = 0;
    exp_40_ram[219] = 39;
    exp_40_ram[220] = 144;
    exp_40_ram[221] = 39;
    exp_40_ram[222] = 247;
    exp_40_ram[223] = 128;
    exp_40_ram[224] = 0;
    exp_40_ram[225] = 39;
    exp_40_ram[226] = 135;
    exp_40_ram[227] = 42;
    exp_40_ram[228] = 39;
    exp_40_ram[229] = 38;
    exp_40_ram[230] = 134;
    exp_40_ram[231] = 37;
    exp_40_ram[232] = 5;
    exp_40_ram[233] = 0;
    exp_40_ram[234] = 39;
    exp_40_ram[235] = 39;
    exp_40_ram[236] = 7;
    exp_40_ram[237] = 39;
    exp_40_ram[238] = 230;
    exp_40_ram[239] = 39;
    exp_40_ram[240] = 133;
    exp_40_ram[241] = 32;
    exp_40_ram[242] = 36;
    exp_40_ram[243] = 1;
    exp_40_ram[244] = 128;
    exp_40_ram[245] = 1;
    exp_40_ram[246] = 38;
    exp_40_ram[247] = 36;
    exp_40_ram[248] = 4;
    exp_40_ram[249] = 38;
    exp_40_ram[250] = 36;
    exp_40_ram[251] = 34;
    exp_40_ram[252] = 32;
    exp_40_ram[253] = 46;
    exp_40_ram[254] = 44;
    exp_40_ram[255] = 7;
    exp_40_ram[256] = 40;
    exp_40_ram[257] = 11;
    exp_40_ram[258] = 39;
    exp_40_ram[259] = 247;
    exp_40_ram[260] = 154;
    exp_40_ram[261] = 39;
    exp_40_ram[262] = 136;
    exp_40_ram[263] = 39;
    exp_40_ram[264] = 247;
    exp_40_ram[265] = 130;
    exp_40_ram[266] = 71;
    exp_40_ram[267] = 152;
    exp_40_ram[268] = 39;
    exp_40_ram[269] = 247;
    exp_40_ram[270] = 136;
    exp_40_ram[271] = 39;
    exp_40_ram[272] = 135;
    exp_40_ram[273] = 34;
    exp_40_ram[274] = 0;
    exp_40_ram[275] = 39;
    exp_40_ram[276] = 135;
    exp_40_ram[277] = 44;
    exp_40_ram[278] = 39;
    exp_40_ram[279] = 7;
    exp_40_ram[280] = 7;
    exp_40_ram[281] = 128;
    exp_40_ram[282] = 39;
    exp_40_ram[283] = 39;
    exp_40_ram[284] = 120;
    exp_40_ram[285] = 39;
    exp_40_ram[286] = 7;
    exp_40_ram[287] = 248;
    exp_40_ram[288] = 0;
    exp_40_ram[289] = 39;
    exp_40_ram[290] = 135;
    exp_40_ram[291] = 44;
    exp_40_ram[292] = 39;
    exp_40_ram[293] = 7;
    exp_40_ram[294] = 7;
    exp_40_ram[295] = 128;
    exp_40_ram[296] = 39;
    exp_40_ram[297] = 247;
    exp_40_ram[298] = 142;
    exp_40_ram[299] = 39;
    exp_40_ram[300] = 39;
    exp_40_ram[301] = 120;
    exp_40_ram[302] = 39;
    exp_40_ram[303] = 7;
    exp_40_ram[304] = 242;
    exp_40_ram[305] = 39;
    exp_40_ram[306] = 247;
    exp_40_ram[307] = 128;
    exp_40_ram[308] = 39;
    exp_40_ram[309] = 247;
    exp_40_ram[310] = 152;
    exp_40_ram[311] = 39;
    exp_40_ram[312] = 132;
    exp_40_ram[313] = 39;
    exp_40_ram[314] = 39;
    exp_40_ram[315] = 8;
    exp_40_ram[316] = 39;
    exp_40_ram[317] = 39;
    exp_40_ram[318] = 24;
    exp_40_ram[319] = 39;
    exp_40_ram[320] = 135;
    exp_40_ram[321] = 44;
    exp_40_ram[322] = 39;
    exp_40_ram[323] = 142;
    exp_40_ram[324] = 39;
    exp_40_ram[325] = 7;
    exp_40_ram[326] = 24;
    exp_40_ram[327] = 39;
    exp_40_ram[328] = 135;
    exp_40_ram[329] = 44;
    exp_40_ram[330] = 39;
    exp_40_ram[331] = 7;
    exp_40_ram[332] = 30;
    exp_40_ram[333] = 39;
    exp_40_ram[334] = 247;
    exp_40_ram[335] = 152;
    exp_40_ram[336] = 39;
    exp_40_ram[337] = 7;
    exp_40_ram[338] = 226;
    exp_40_ram[339] = 39;
    exp_40_ram[340] = 135;
    exp_40_ram[341] = 44;
    exp_40_ram[342] = 39;
    exp_40_ram[343] = 7;
    exp_40_ram[344] = 7;
    exp_40_ram[345] = 128;
    exp_40_ram[346] = 0;
    exp_40_ram[347] = 39;
    exp_40_ram[348] = 7;
    exp_40_ram[349] = 30;
    exp_40_ram[350] = 39;
    exp_40_ram[351] = 247;
    exp_40_ram[352] = 136;
    exp_40_ram[353] = 39;
    exp_40_ram[354] = 7;
    exp_40_ram[355] = 226;
    exp_40_ram[356] = 39;
    exp_40_ram[357] = 135;
    exp_40_ram[358] = 44;
    exp_40_ram[359] = 39;
    exp_40_ram[360] = 7;
    exp_40_ram[361] = 7;
    exp_40_ram[362] = 128;
    exp_40_ram[363] = 0;
    exp_40_ram[364] = 39;
    exp_40_ram[365] = 7;
    exp_40_ram[366] = 22;
    exp_40_ram[367] = 39;
    exp_40_ram[368] = 7;
    exp_40_ram[369] = 224;
    exp_40_ram[370] = 39;
    exp_40_ram[371] = 135;
    exp_40_ram[372] = 44;
    exp_40_ram[373] = 39;
    exp_40_ram[374] = 7;
    exp_40_ram[375] = 7;
    exp_40_ram[376] = 128;
    exp_40_ram[377] = 39;
    exp_40_ram[378] = 7;
    exp_40_ram[379] = 224;
    exp_40_ram[380] = 39;
    exp_40_ram[381] = 135;
    exp_40_ram[382] = 44;
    exp_40_ram[383] = 39;
    exp_40_ram[384] = 7;
    exp_40_ram[385] = 7;
    exp_40_ram[386] = 128;
    exp_40_ram[387] = 39;
    exp_40_ram[388] = 7;
    exp_40_ram[389] = 224;
    exp_40_ram[390] = 71;
    exp_40_ram[391] = 130;
    exp_40_ram[392] = 39;
    exp_40_ram[393] = 135;
    exp_40_ram[394] = 44;
    exp_40_ram[395] = 39;
    exp_40_ram[396] = 7;
    exp_40_ram[397] = 7;
    exp_40_ram[398] = 128;
    exp_40_ram[399] = 0;
    exp_40_ram[400] = 39;
    exp_40_ram[401] = 247;
    exp_40_ram[402] = 130;
    exp_40_ram[403] = 39;
    exp_40_ram[404] = 135;
    exp_40_ram[405] = 44;
    exp_40_ram[406] = 39;
    exp_40_ram[407] = 7;
    exp_40_ram[408] = 7;
    exp_40_ram[409] = 128;
    exp_40_ram[410] = 0;
    exp_40_ram[411] = 39;
    exp_40_ram[412] = 247;
    exp_40_ram[413] = 128;
    exp_40_ram[414] = 39;
    exp_40_ram[415] = 135;
    exp_40_ram[416] = 44;
    exp_40_ram[417] = 39;
    exp_40_ram[418] = 7;
    exp_40_ram[419] = 7;
    exp_40_ram[420] = 128;
    exp_40_ram[421] = 40;
    exp_40_ram[422] = 40;
    exp_40_ram[423] = 39;
    exp_40_ram[424] = 39;
    exp_40_ram[425] = 38;
    exp_40_ram[426] = 38;
    exp_40_ram[427] = 37;
    exp_40_ram[428] = 37;
    exp_40_ram[429] = 240;
    exp_40_ram[430] = 7;
    exp_40_ram[431] = 133;
    exp_40_ram[432] = 32;
    exp_40_ram[433] = 36;
    exp_40_ram[434] = 1;
    exp_40_ram[435] = 128;
    exp_40_ram[436] = 1;
    exp_40_ram[437] = 38;
    exp_40_ram[438] = 36;
    exp_40_ram[439] = 4;
    exp_40_ram[440] = 46;
    exp_40_ram[441] = 44;
    exp_40_ram[442] = 42;
    exp_40_ram[443] = 40;
    exp_40_ram[444] = 38;
    exp_40_ram[445] = 34;
    exp_40_ram[446] = 32;
    exp_40_ram[447] = 5;
    exp_40_ram[448] = 38;
    exp_40_ram[449] = 39;
    exp_40_ram[450] = 152;
    exp_40_ram[451] = 39;
    exp_40_ram[452] = 247;
    exp_40_ram[453] = 34;
    exp_40_ram[454] = 39;
    exp_40_ram[455] = 247;
    exp_40_ram[456] = 134;
    exp_40_ram[457] = 39;
    exp_40_ram[458] = 140;
    exp_40_ram[459] = 39;
    exp_40_ram[460] = 39;
    exp_40_ram[461] = 119;
    exp_40_ram[462] = 5;
    exp_40_ram[463] = 71;
    exp_40_ram[464] = 7;
    exp_40_ram[465] = 234;
    exp_40_ram[466] = 71;
    exp_40_ram[467] = 135;
    exp_40_ram[468] = 247;
    exp_40_ram[469] = 0;
    exp_40_ram[470] = 39;
    exp_40_ram[471] = 247;
    exp_40_ram[472] = 134;
    exp_40_ram[473] = 7;
    exp_40_ram[474] = 0;
    exp_40_ram[475] = 7;
    exp_40_ram[476] = 71;
    exp_40_ram[477] = 135;
    exp_40_ram[478] = 247;
    exp_40_ram[479] = 135;
    exp_40_ram[480] = 247;
    exp_40_ram[481] = 39;
    exp_40_ram[482] = 6;
    exp_40_ram[483] = 38;
    exp_40_ram[484] = 6;
    exp_40_ram[485] = 135;
    exp_40_ram[486] = 12;
    exp_40_ram[487] = 39;
    exp_40_ram[488] = 39;
    exp_40_ram[489] = 87;
    exp_40_ram[490] = 38;
    exp_40_ram[491] = 39;
    exp_40_ram[492] = 136;
    exp_40_ram[493] = 39;
    exp_40_ram[494] = 7;
    exp_40_ram[495] = 248;
    exp_40_ram[496] = 70;
    exp_40_ram[497] = 7;
    exp_40_ram[498] = 39;
    exp_40_ram[499] = 36;
    exp_40_ram[500] = 39;
    exp_40_ram[501] = 34;
    exp_40_ram[502] = 39;
    exp_40_ram[503] = 32;
    exp_40_ram[504] = 40;
    exp_40_ram[505] = 136;
    exp_40_ram[506] = 39;
    exp_40_ram[507] = 38;
    exp_40_ram[508] = 38;
    exp_40_ram[509] = 37;
    exp_40_ram[510] = 37;
    exp_40_ram[511] = 240;
    exp_40_ram[512] = 7;
    exp_40_ram[513] = 133;
    exp_40_ram[514] = 32;
    exp_40_ram[515] = 36;
    exp_40_ram[516] = 1;
    exp_40_ram[517] = 128;
    exp_40_ram[518] = 1;
    exp_40_ram[519] = 46;
    exp_40_ram[520] = 44;
    exp_40_ram[521] = 4;
    exp_40_ram[522] = 38;
    exp_40_ram[523] = 36;
    exp_40_ram[524] = 34;
    exp_40_ram[525] = 32;
    exp_40_ram[526] = 46;
    exp_40_ram[527] = 46;
    exp_40_ram[528] = 39;
    exp_40_ram[529] = 156;
    exp_40_ram[530] = 7;
    exp_40_ram[531] = 38;
    exp_40_ram[532] = 0;
    exp_40_ram[533] = 39;
    exp_40_ram[534] = 199;
    exp_40_ram[535] = 7;
    exp_40_ram[536] = 14;
    exp_40_ram[537] = 39;
    exp_40_ram[538] = 197;
    exp_40_ram[539] = 39;
    exp_40_ram[540] = 135;
    exp_40_ram[541] = 46;
    exp_40_ram[542] = 39;
    exp_40_ram[543] = 38;
    exp_40_ram[544] = 134;
    exp_40_ram[545] = 37;
    exp_40_ram[546] = 0;
    exp_40_ram[547] = 39;
    exp_40_ram[548] = 135;
    exp_40_ram[549] = 32;
    exp_40_ram[550] = 0;
    exp_40_ram[551] = 39;
    exp_40_ram[552] = 135;
    exp_40_ram[553] = 32;
    exp_40_ram[554] = 38;
    exp_40_ram[555] = 39;
    exp_40_ram[556] = 199;
    exp_40_ram[557] = 135;
    exp_40_ram[558] = 7;
    exp_40_ram[559] = 104;
    exp_40_ram[560] = 151;
    exp_40_ram[561] = 23;
    exp_40_ram[562] = 135;
    exp_40_ram[563] = 7;
    exp_40_ram[564] = 167;
    exp_40_ram[565] = 128;
    exp_40_ram[566] = 39;
    exp_40_ram[567] = 231;
    exp_40_ram[568] = 38;
    exp_40_ram[569] = 39;
    exp_40_ram[570] = 135;
    exp_40_ram[571] = 32;
    exp_40_ram[572] = 7;
    exp_40_ram[573] = 32;
    exp_40_ram[574] = 0;
    exp_40_ram[575] = 39;
    exp_40_ram[576] = 231;
    exp_40_ram[577] = 38;
    exp_40_ram[578] = 39;
    exp_40_ram[579] = 135;
    exp_40_ram[580] = 32;
    exp_40_ram[581] = 7;
    exp_40_ram[582] = 32;
    exp_40_ram[583] = 0;
    exp_40_ram[584] = 39;
    exp_40_ram[585] = 231;
    exp_40_ram[586] = 38;
    exp_40_ram[587] = 39;
    exp_40_ram[588] = 135;
    exp_40_ram[589] = 32;
    exp_40_ram[590] = 7;
    exp_40_ram[591] = 32;
    exp_40_ram[592] = 0;
    exp_40_ram[593] = 39;
    exp_40_ram[594] = 231;
    exp_40_ram[595] = 38;
    exp_40_ram[596] = 39;
    exp_40_ram[597] = 135;
    exp_40_ram[598] = 32;
    exp_40_ram[599] = 7;
    exp_40_ram[600] = 32;
    exp_40_ram[601] = 0;
    exp_40_ram[602] = 39;
    exp_40_ram[603] = 231;
    exp_40_ram[604] = 38;
    exp_40_ram[605] = 39;
    exp_40_ram[606] = 135;
    exp_40_ram[607] = 32;
    exp_40_ram[608] = 7;
    exp_40_ram[609] = 32;
    exp_40_ram[610] = 0;
    exp_40_ram[611] = 32;
    exp_40_ram[612] = 0;
    exp_40_ram[613] = 39;
    exp_40_ram[614] = 154;
    exp_40_ram[615] = 36;
    exp_40_ram[616] = 39;
    exp_40_ram[617] = 199;
    exp_40_ram[618] = 133;
    exp_40_ram[619] = 240;
    exp_40_ram[620] = 7;
    exp_40_ram[621] = 140;
    exp_40_ram[622] = 7;
    exp_40_ram[623] = 133;
    exp_40_ram[624] = 240;
    exp_40_ram[625] = 36;
    exp_40_ram[626] = 0;
    exp_40_ram[627] = 39;
    exp_40_ram[628] = 199;
    exp_40_ram[629] = 7;
    exp_40_ram[630] = 24;
    exp_40_ram[631] = 39;
    exp_40_ram[632] = 135;
    exp_40_ram[633] = 46;
    exp_40_ram[634] = 167;
    exp_40_ram[635] = 36;
    exp_40_ram[636] = 39;
    exp_40_ram[637] = 208;
    exp_40_ram[638] = 39;
    exp_40_ram[639] = 231;
    exp_40_ram[640] = 38;
    exp_40_ram[641] = 39;
    exp_40_ram[642] = 7;
    exp_40_ram[643] = 36;
    exp_40_ram[644] = 0;
    exp_40_ram[645] = 39;
    exp_40_ram[646] = 36;
    exp_40_ram[647] = 39;
    exp_40_ram[648] = 135;
    exp_40_ram[649] = 32;
    exp_40_ram[650] = 34;
    exp_40_ram[651] = 39;
    exp_40_ram[652] = 199;
    exp_40_ram[653] = 7;
    exp_40_ram[654] = 20;
    exp_40_ram[655] = 39;
    exp_40_ram[656] = 231;
    exp_40_ram[657] = 38;
    exp_40_ram[658] = 39;
    exp_40_ram[659] = 135;
    exp_40_ram[660] = 32;
    exp_40_ram[661] = 39;
    exp_40_ram[662] = 199;
    exp_40_ram[663] = 133;
    exp_40_ram[664] = 240;
    exp_40_ram[665] = 7;
    exp_40_ram[666] = 140;
    exp_40_ram[667] = 7;
    exp_40_ram[668] = 133;
    exp_40_ram[669] = 240;
    exp_40_ram[670] = 34;
    exp_40_ram[671] = 0;
    exp_40_ram[672] = 39;
    exp_40_ram[673] = 199;
    exp_40_ram[674] = 7;
    exp_40_ram[675] = 26;
    exp_40_ram[676] = 39;
    exp_40_ram[677] = 135;
    exp_40_ram[678] = 46;
    exp_40_ram[679] = 167;
    exp_40_ram[680] = 34;
    exp_40_ram[681] = 39;
    exp_40_ram[682] = 212;
    exp_40_ram[683] = 7;
    exp_40_ram[684] = 34;
    exp_40_ram[685] = 39;
    exp_40_ram[686] = 135;
    exp_40_ram[687] = 32;
    exp_40_ram[688] = 39;
    exp_40_ram[689] = 199;
    exp_40_ram[690] = 135;
    exp_40_ram[691] = 7;
    exp_40_ram[692] = 108;
    exp_40_ram[693] = 151;
    exp_40_ram[694] = 23;
    exp_40_ram[695] = 135;
    exp_40_ram[696] = 7;
    exp_40_ram[697] = 167;
    exp_40_ram[698] = 128;
    exp_40_ram[699] = 39;
    exp_40_ram[700] = 231;
    exp_40_ram[701] = 38;
    exp_40_ram[702] = 39;
    exp_40_ram[703] = 135;
    exp_40_ram[704] = 32;
    exp_40_ram[705] = 39;
    exp_40_ram[706] = 199;
    exp_40_ram[707] = 7;
    exp_40_ram[708] = 16;
    exp_40_ram[709] = 39;
    exp_40_ram[710] = 231;
    exp_40_ram[711] = 38;
    exp_40_ram[712] = 39;
    exp_40_ram[713] = 135;
    exp_40_ram[714] = 32;
    exp_40_ram[715] = 0;
    exp_40_ram[716] = 39;
    exp_40_ram[717] = 231;
    exp_40_ram[718] = 38;
    exp_40_ram[719] = 39;
    exp_40_ram[720] = 135;
    exp_40_ram[721] = 32;
    exp_40_ram[722] = 39;
    exp_40_ram[723] = 199;
    exp_40_ram[724] = 7;
    exp_40_ram[725] = 18;
    exp_40_ram[726] = 39;
    exp_40_ram[727] = 231;
    exp_40_ram[728] = 38;
    exp_40_ram[729] = 39;
    exp_40_ram[730] = 135;
    exp_40_ram[731] = 32;
    exp_40_ram[732] = 0;
    exp_40_ram[733] = 39;
    exp_40_ram[734] = 231;
    exp_40_ram[735] = 38;
    exp_40_ram[736] = 39;
    exp_40_ram[737] = 135;
    exp_40_ram[738] = 32;
    exp_40_ram[739] = 0;
    exp_40_ram[740] = 39;
    exp_40_ram[741] = 231;
    exp_40_ram[742] = 38;
    exp_40_ram[743] = 39;
    exp_40_ram[744] = 135;
    exp_40_ram[745] = 32;
    exp_40_ram[746] = 0;
    exp_40_ram[747] = 39;
    exp_40_ram[748] = 231;
    exp_40_ram[749] = 38;
    exp_40_ram[750] = 39;
    exp_40_ram[751] = 135;
    exp_40_ram[752] = 32;
    exp_40_ram[753] = 0;
    exp_40_ram[754] = 0;
    exp_40_ram[755] = 0;
    exp_40_ram[756] = 0;
    exp_40_ram[757] = 0;
    exp_40_ram[758] = 0;
    exp_40_ram[759] = 39;
    exp_40_ram[760] = 199;
    exp_40_ram[761] = 135;
    exp_40_ram[762] = 7;
    exp_40_ram[763] = 108;
    exp_40_ram[764] = 151;
    exp_40_ram[765] = 23;
    exp_40_ram[766] = 135;
    exp_40_ram[767] = 7;
    exp_40_ram[768] = 167;
    exp_40_ram[769] = 128;
    exp_40_ram[770] = 39;
    exp_40_ram[771] = 199;
    exp_40_ram[772] = 7;
    exp_40_ram[773] = 10;
    exp_40_ram[774] = 39;
    exp_40_ram[775] = 199;
    exp_40_ram[776] = 7;
    exp_40_ram[777] = 24;
    exp_40_ram[778] = 7;
    exp_40_ram[779] = 44;
    exp_40_ram[780] = 0;
    exp_40_ram[781] = 39;
    exp_40_ram[782] = 199;
    exp_40_ram[783] = 7;
    exp_40_ram[784] = 24;
    exp_40_ram[785] = 7;
    exp_40_ram[786] = 44;
    exp_40_ram[787] = 0;
    exp_40_ram[788] = 39;
    exp_40_ram[789] = 199;
    exp_40_ram[790] = 7;
    exp_40_ram[791] = 24;
    exp_40_ram[792] = 7;
    exp_40_ram[793] = 44;
    exp_40_ram[794] = 0;
    exp_40_ram[795] = 7;
    exp_40_ram[796] = 44;
    exp_40_ram[797] = 39;
    exp_40_ram[798] = 247;
    exp_40_ram[799] = 38;
    exp_40_ram[800] = 39;
    exp_40_ram[801] = 199;
    exp_40_ram[802] = 7;
    exp_40_ram[803] = 24;
    exp_40_ram[804] = 39;
    exp_40_ram[805] = 231;
    exp_40_ram[806] = 38;
    exp_40_ram[807] = 39;
    exp_40_ram[808] = 199;
    exp_40_ram[809] = 7;
    exp_40_ram[810] = 0;
    exp_40_ram[811] = 39;
    exp_40_ram[812] = 199;
    exp_40_ram[813] = 7;
    exp_40_ram[814] = 8;
    exp_40_ram[815] = 39;
    exp_40_ram[816] = 247;
    exp_40_ram[817] = 38;
    exp_40_ram[818] = 39;
    exp_40_ram[819] = 247;
    exp_40_ram[820] = 136;
    exp_40_ram[821] = 39;
    exp_40_ram[822] = 247;
    exp_40_ram[823] = 38;
    exp_40_ram[824] = 39;
    exp_40_ram[825] = 199;
    exp_40_ram[826] = 7;
    exp_40_ram[827] = 10;
    exp_40_ram[828] = 39;
    exp_40_ram[829] = 199;
    exp_40_ram[830] = 7;
    exp_40_ram[831] = 24;
    exp_40_ram[832] = 39;
    exp_40_ram[833] = 247;
    exp_40_ram[834] = 158;
    exp_40_ram[835] = 39;
    exp_40_ram[836] = 247;
    exp_40_ram[837] = 140;
    exp_40_ram[838] = 39;
    exp_40_ram[839] = 135;
    exp_40_ram[840] = 46;
    exp_40_ram[841] = 167;
    exp_40_ram[842] = 44;
    exp_40_ram[843] = 39;
    exp_40_ram[844] = 215;
    exp_40_ram[845] = 39;
    exp_40_ram[846] = 71;
    exp_40_ram[847] = 135;
    exp_40_ram[848] = 134;
    exp_40_ram[849] = 39;
    exp_40_ram[850] = 215;
    exp_40_ram[851] = 247;
    exp_40_ram[852] = 39;
    exp_40_ram[853] = 34;
    exp_40_ram[854] = 39;
    exp_40_ram[855] = 32;
    exp_40_ram[856] = 40;
    exp_40_ram[857] = 40;
    exp_40_ram[858] = 7;
    exp_40_ram[859] = 135;
    exp_40_ram[860] = 38;
    exp_40_ram[861] = 38;
    exp_40_ram[862] = 37;
    exp_40_ram[863] = 37;
    exp_40_ram[864] = 240;
    exp_40_ram[865] = 46;
    exp_40_ram[866] = 0;
    exp_40_ram[867] = 39;
    exp_40_ram[868] = 247;
    exp_40_ram[869] = 142;
    exp_40_ram[870] = 39;
    exp_40_ram[871] = 135;
    exp_40_ram[872] = 46;
    exp_40_ram[873] = 167;
    exp_40_ram[874] = 247;
    exp_40_ram[875] = 0;
    exp_40_ram[876] = 39;
    exp_40_ram[877] = 247;
    exp_40_ram[878] = 128;
    exp_40_ram[879] = 39;
    exp_40_ram[880] = 135;
    exp_40_ram[881] = 46;
    exp_40_ram[882] = 167;
    exp_40_ram[883] = 151;
    exp_40_ram[884] = 215;
    exp_40_ram[885] = 0;
    exp_40_ram[886] = 39;
    exp_40_ram[887] = 135;
    exp_40_ram[888] = 46;
    exp_40_ram[889] = 167;
    exp_40_ram[890] = 46;
    exp_40_ram[891] = 39;
    exp_40_ram[892] = 215;
    exp_40_ram[893] = 39;
    exp_40_ram[894] = 71;
    exp_40_ram[895] = 135;
    exp_40_ram[896] = 134;
    exp_40_ram[897] = 39;
    exp_40_ram[898] = 215;
    exp_40_ram[899] = 247;
    exp_40_ram[900] = 39;
    exp_40_ram[901] = 34;
    exp_40_ram[902] = 39;
    exp_40_ram[903] = 32;
    exp_40_ram[904] = 40;
    exp_40_ram[905] = 40;
    exp_40_ram[906] = 7;
    exp_40_ram[907] = 135;
    exp_40_ram[908] = 38;
    exp_40_ram[909] = 38;
    exp_40_ram[910] = 37;
    exp_40_ram[911] = 37;
    exp_40_ram[912] = 240;
    exp_40_ram[913] = 46;
    exp_40_ram[914] = 0;
    exp_40_ram[915] = 39;
    exp_40_ram[916] = 247;
    exp_40_ram[917] = 152;
    exp_40_ram[918] = 39;
    exp_40_ram[919] = 247;
    exp_40_ram[920] = 134;
    exp_40_ram[921] = 39;
    exp_40_ram[922] = 135;
    exp_40_ram[923] = 46;
    exp_40_ram[924] = 167;
    exp_40_ram[925] = 39;
    exp_40_ram[926] = 34;
    exp_40_ram[927] = 39;
    exp_40_ram[928] = 32;
    exp_40_ram[929] = 40;
    exp_40_ram[930] = 40;
    exp_40_ram[931] = 7;
    exp_40_ram[932] = 38;
    exp_40_ram[933] = 38;
    exp_40_ram[934] = 37;
    exp_40_ram[935] = 37;
    exp_40_ram[936] = 240;
    exp_40_ram[937] = 46;
    exp_40_ram[938] = 0;
    exp_40_ram[939] = 39;
    exp_40_ram[940] = 247;
    exp_40_ram[941] = 142;
    exp_40_ram[942] = 39;
    exp_40_ram[943] = 135;
    exp_40_ram[944] = 46;
    exp_40_ram[945] = 167;
    exp_40_ram[946] = 247;
    exp_40_ram[947] = 0;
    exp_40_ram[948] = 39;
    exp_40_ram[949] = 247;
    exp_40_ram[950] = 128;
    exp_40_ram[951] = 39;
    exp_40_ram[952] = 135;
    exp_40_ram[953] = 46;
    exp_40_ram[954] = 167;
    exp_40_ram[955] = 151;
    exp_40_ram[956] = 215;
    exp_40_ram[957] = 0;
    exp_40_ram[958] = 39;
    exp_40_ram[959] = 135;
    exp_40_ram[960] = 46;
    exp_40_ram[961] = 167;
    exp_40_ram[962] = 32;
    exp_40_ram[963] = 39;
    exp_40_ram[964] = 34;
    exp_40_ram[965] = 39;
    exp_40_ram[966] = 32;
    exp_40_ram[967] = 40;
    exp_40_ram[968] = 40;
    exp_40_ram[969] = 7;
    exp_40_ram[970] = 39;
    exp_40_ram[971] = 38;
    exp_40_ram[972] = 38;
    exp_40_ram[973] = 37;
    exp_40_ram[974] = 37;
    exp_40_ram[975] = 240;
    exp_40_ram[976] = 46;
    exp_40_ram[977] = 39;
    exp_40_ram[978] = 135;
    exp_40_ram[979] = 32;
    exp_40_ram[980] = 0;
    exp_40_ram[981] = 7;
    exp_40_ram[982] = 42;
    exp_40_ram[983] = 39;
    exp_40_ram[984] = 247;
    exp_40_ram[985] = 144;
    exp_40_ram[986] = 0;
    exp_40_ram[987] = 39;
    exp_40_ram[988] = 135;
    exp_40_ram[989] = 46;
    exp_40_ram[990] = 39;
    exp_40_ram[991] = 38;
    exp_40_ram[992] = 134;
    exp_40_ram[993] = 37;
    exp_40_ram[994] = 5;
    exp_40_ram[995] = 0;
    exp_40_ram[996] = 39;
    exp_40_ram[997] = 135;
    exp_40_ram[998] = 42;
    exp_40_ram[999] = 39;
    exp_40_ram[1000] = 230;
    exp_40_ram[1001] = 39;
    exp_40_ram[1002] = 135;
    exp_40_ram[1003] = 46;
    exp_40_ram[1004] = 167;
    exp_40_ram[1005] = 245;
    exp_40_ram[1006] = 39;
    exp_40_ram[1007] = 135;
    exp_40_ram[1008] = 46;
    exp_40_ram[1009] = 39;
    exp_40_ram[1010] = 38;
    exp_40_ram[1011] = 134;
    exp_40_ram[1012] = 37;
    exp_40_ram[1013] = 0;
    exp_40_ram[1014] = 39;
    exp_40_ram[1015] = 247;
    exp_40_ram[1016] = 128;
    exp_40_ram[1017] = 0;
    exp_40_ram[1018] = 39;
    exp_40_ram[1019] = 135;
    exp_40_ram[1020] = 46;
    exp_40_ram[1021] = 39;
    exp_40_ram[1022] = 38;
    exp_40_ram[1023] = 134;
    exp_40_ram[1024] = 37;
    exp_40_ram[1025] = 5;
    exp_40_ram[1026] = 0;
    exp_40_ram[1027] = 39;
    exp_40_ram[1028] = 135;
    exp_40_ram[1029] = 42;
    exp_40_ram[1030] = 39;
    exp_40_ram[1031] = 230;
    exp_40_ram[1032] = 39;
    exp_40_ram[1033] = 135;
    exp_40_ram[1034] = 32;
    exp_40_ram[1035] = 0;
    exp_40_ram[1036] = 39;
    exp_40_ram[1037] = 135;
    exp_40_ram[1038] = 46;
    exp_40_ram[1039] = 167;
    exp_40_ram[1040] = 40;
    exp_40_ram[1041] = 39;
    exp_40_ram[1042] = 134;
    exp_40_ram[1043] = 39;
    exp_40_ram[1044] = 0;
    exp_40_ram[1045] = 7;
    exp_40_ram[1046] = 133;
    exp_40_ram[1047] = 37;
    exp_40_ram[1048] = 240;
    exp_40_ram[1049] = 38;
    exp_40_ram[1050] = 39;
    exp_40_ram[1051] = 247;
    exp_40_ram[1052] = 140;
    exp_40_ram[1053] = 39;
    exp_40_ram[1054] = 39;
    exp_40_ram[1055] = 116;
    exp_40_ram[1056] = 7;
    exp_40_ram[1057] = 38;
    exp_40_ram[1058] = 39;
    exp_40_ram[1059] = 247;
    exp_40_ram[1060] = 154;
    exp_40_ram[1061] = 0;
    exp_40_ram[1062] = 39;
    exp_40_ram[1063] = 135;
    exp_40_ram[1064] = 46;
    exp_40_ram[1065] = 39;
    exp_40_ram[1066] = 38;
    exp_40_ram[1067] = 134;
    exp_40_ram[1068] = 37;
    exp_40_ram[1069] = 5;
    exp_40_ram[1070] = 0;
    exp_40_ram[1071] = 39;
    exp_40_ram[1072] = 135;
    exp_40_ram[1073] = 38;
    exp_40_ram[1074] = 39;
    exp_40_ram[1075] = 230;
    exp_40_ram[1076] = 0;
    exp_40_ram[1077] = 39;
    exp_40_ram[1078] = 135;
    exp_40_ram[1079] = 40;
    exp_40_ram[1080] = 197;
    exp_40_ram[1081] = 39;
    exp_40_ram[1082] = 135;
    exp_40_ram[1083] = 46;
    exp_40_ram[1084] = 39;
    exp_40_ram[1085] = 38;
    exp_40_ram[1086] = 134;
    exp_40_ram[1087] = 37;
    exp_40_ram[1088] = 0;
    exp_40_ram[1089] = 39;
    exp_40_ram[1090] = 199;
    exp_40_ram[1091] = 128;
    exp_40_ram[1092] = 39;
    exp_40_ram[1093] = 247;
    exp_40_ram[1094] = 142;
    exp_40_ram[1095] = 39;
    exp_40_ram[1096] = 135;
    exp_40_ram[1097] = 34;
    exp_40_ram[1098] = 150;
    exp_40_ram[1099] = 39;
    exp_40_ram[1100] = 247;
    exp_40_ram[1101] = 128;
    exp_40_ram[1102] = 0;
    exp_40_ram[1103] = 39;
    exp_40_ram[1104] = 135;
    exp_40_ram[1105] = 46;
    exp_40_ram[1106] = 39;
    exp_40_ram[1107] = 38;
    exp_40_ram[1108] = 134;
    exp_40_ram[1109] = 37;
    exp_40_ram[1110] = 5;
    exp_40_ram[1111] = 0;
    exp_40_ram[1112] = 39;
    exp_40_ram[1113] = 135;
    exp_40_ram[1114] = 38;
    exp_40_ram[1115] = 39;
    exp_40_ram[1116] = 230;
    exp_40_ram[1117] = 39;
    exp_40_ram[1118] = 135;
    exp_40_ram[1119] = 32;
    exp_40_ram[1120] = 0;
    exp_40_ram[1121] = 7;
    exp_40_ram[1122] = 36;
    exp_40_ram[1123] = 39;
    exp_40_ram[1124] = 231;
    exp_40_ram[1125] = 38;
    exp_40_ram[1126] = 39;
    exp_40_ram[1127] = 135;
    exp_40_ram[1128] = 46;
    exp_40_ram[1129] = 167;
    exp_40_ram[1130] = 135;
    exp_40_ram[1131] = 39;
    exp_40_ram[1132] = 34;
    exp_40_ram[1133] = 39;
    exp_40_ram[1134] = 32;
    exp_40_ram[1135] = 40;
    exp_40_ram[1136] = 8;
    exp_40_ram[1137] = 7;
    exp_40_ram[1138] = 38;
    exp_40_ram[1139] = 38;
    exp_40_ram[1140] = 37;
    exp_40_ram[1141] = 37;
    exp_40_ram[1142] = 240;
    exp_40_ram[1143] = 46;
    exp_40_ram[1144] = 39;
    exp_40_ram[1145] = 135;
    exp_40_ram[1146] = 32;
    exp_40_ram[1147] = 0;
    exp_40_ram[1148] = 39;
    exp_40_ram[1149] = 135;
    exp_40_ram[1150] = 46;
    exp_40_ram[1151] = 39;
    exp_40_ram[1152] = 38;
    exp_40_ram[1153] = 134;
    exp_40_ram[1154] = 37;
    exp_40_ram[1155] = 5;
    exp_40_ram[1156] = 0;
    exp_40_ram[1157] = 39;
    exp_40_ram[1158] = 135;
    exp_40_ram[1159] = 32;
    exp_40_ram[1160] = 0;
    exp_40_ram[1161] = 39;
    exp_40_ram[1162] = 197;
    exp_40_ram[1163] = 39;
    exp_40_ram[1164] = 135;
    exp_40_ram[1165] = 46;
    exp_40_ram[1166] = 39;
    exp_40_ram[1167] = 38;
    exp_40_ram[1168] = 134;
    exp_40_ram[1169] = 37;
    exp_40_ram[1170] = 0;
    exp_40_ram[1171] = 39;
    exp_40_ram[1172] = 135;
    exp_40_ram[1173] = 32;
    exp_40_ram[1174] = 0;
    exp_40_ram[1175] = 39;
    exp_40_ram[1176] = 199;
    exp_40_ram[1177] = 152;
    exp_40_ram[1178] = 39;
    exp_40_ram[1179] = 39;
    exp_40_ram[1180] = 104;
    exp_40_ram[1181] = 39;
    exp_40_ram[1182] = 135;
    exp_40_ram[1183] = 0;
    exp_40_ram[1184] = 39;
    exp_40_ram[1185] = 39;
    exp_40_ram[1186] = 38;
    exp_40_ram[1187] = 134;
    exp_40_ram[1188] = 37;
    exp_40_ram[1189] = 5;
    exp_40_ram[1190] = 0;
    exp_40_ram[1191] = 39;
    exp_40_ram[1192] = 133;
    exp_40_ram[1193] = 32;
    exp_40_ram[1194] = 36;
    exp_40_ram[1195] = 1;
    exp_40_ram[1196] = 128;
    exp_40_ram[1197] = 1;
    exp_40_ram[1198] = 38;
    exp_40_ram[1199] = 36;
    exp_40_ram[1200] = 4;
    exp_40_ram[1201] = 46;
    exp_40_ram[1202] = 34;
    exp_40_ram[1203] = 36;
    exp_40_ram[1204] = 38;
    exp_40_ram[1205] = 40;
    exp_40_ram[1206] = 42;
    exp_40_ram[1207] = 44;
    exp_40_ram[1208] = 46;
    exp_40_ram[1209] = 7;
    exp_40_ram[1210] = 44;
    exp_40_ram[1211] = 39;
    exp_40_ram[1212] = 135;
    exp_40_ram[1213] = 36;
    exp_40_ram[1214] = 39;
    exp_40_ram[1215] = 7;
    exp_40_ram[1216] = 38;
    exp_40_ram[1217] = 6;
    exp_40_ram[1218] = 133;
    exp_40_ram[1219] = 5;
    exp_40_ram[1220] = 240;
    exp_40_ram[1221] = 38;
    exp_40_ram[1222] = 39;
    exp_40_ram[1223] = 133;
    exp_40_ram[1224] = 32;
    exp_40_ram[1225] = 36;
    exp_40_ram[1226] = 1;
    exp_40_ram[1227] = 128;
    exp_40_ram[1228] = 1;
    exp_40_ram[1229] = 46;
    exp_40_ram[1230] = 44;
    exp_40_ram[1231] = 4;
    exp_40_ram[1232] = 7;
    exp_40_ram[1233] = 7;
    exp_40_ram[1234] = 71;
    exp_40_ram[1235] = 23;
    exp_40_ram[1236] = 167;
    exp_40_ram[1237] = 133;
    exp_40_ram[1238] = 5;
    exp_40_ram[1239] = 224;
    exp_40_ram[1240] = 0;
    exp_40_ram[1241] = 32;
    exp_40_ram[1242] = 36;
    exp_40_ram[1243] = 1;
    exp_40_ram[1244] = 128;
    exp_40_ram[1245] = 1;
    exp_40_ram[1246] = 38;
    exp_40_ram[1247] = 36;
    exp_40_ram[1248] = 4;
    exp_40_ram[1249] = 5;
    exp_40_ram[1250] = 240;
    exp_40_ram[1251] = 0;
    exp_40_ram[1252] = 32;
    exp_40_ram[1253] = 36;
    exp_40_ram[1254] = 1;
    exp_40_ram[1255] = 128;
    exp_40_ram[1256] = 0;
    exp_40_ram[1257] = 9;
    exp_40_ram[1258] = 9;
    exp_40_ram[1259] = 9;
    exp_40_ram[1260] = 9;
    exp_40_ram[1261] = 9;
    exp_40_ram[1262] = 9;
    exp_40_ram[1263] = 9;
    exp_40_ram[1264] = 9;
    exp_40_ram[1265] = 9;
    exp_40_ram[1266] = 9;
    exp_40_ram[1267] = 9;
    exp_40_ram[1268] = 9;
    exp_40_ram[1269] = 9;
    exp_40_ram[1270] = 8;
    exp_40_ram[1271] = 9;
    exp_40_ram[1272] = 9;
    exp_40_ram[1273] = 8;
    exp_40_ram[1274] = 11;
    exp_40_ram[1275] = 11;
    exp_40_ram[1276] = 11;
    exp_40_ram[1277] = 11;
    exp_40_ram[1278] = 10;
    exp_40_ram[1279] = 11;
    exp_40_ram[1280] = 11;
    exp_40_ram[1281] = 11;
    exp_40_ram[1282] = 11;
    exp_40_ram[1283] = 11;
    exp_40_ram[1284] = 11;
    exp_40_ram[1285] = 11;
    exp_40_ram[1286] = 11;
    exp_40_ram[1287] = 11;
    exp_40_ram[1288] = 11;
    exp_40_ram[1289] = 11;
    exp_40_ram[1290] = 11;
    exp_40_ram[1291] = 11;
    exp_40_ram[1292] = 11;
    exp_40_ram[1293] = 17;
    exp_40_ram[1294] = 18;
    exp_40_ram[1295] = 18;
    exp_40_ram[1296] = 18;
    exp_40_ram[1297] = 18;
    exp_40_ram[1298] = 18;
    exp_40_ram[1299] = 18;
    exp_40_ram[1300] = 18;
    exp_40_ram[1301] = 18;
    exp_40_ram[1302] = 18;
    exp_40_ram[1303] = 18;
    exp_40_ram[1304] = 18;
    exp_40_ram[1305] = 18;
    exp_40_ram[1306] = 18;
    exp_40_ram[1307] = 18;
    exp_40_ram[1308] = 18;
    exp_40_ram[1309] = 18;
    exp_40_ram[1310] = 18;
    exp_40_ram[1311] = 18;
    exp_40_ram[1312] = 18;
    exp_40_ram[1313] = 18;
    exp_40_ram[1314] = 18;
    exp_40_ram[1315] = 18;
    exp_40_ram[1316] = 18;
    exp_40_ram[1317] = 18;
    exp_40_ram[1318] = 18;
    exp_40_ram[1319] = 18;
    exp_40_ram[1320] = 18;
    exp_40_ram[1321] = 18;
    exp_40_ram[1322] = 18;
    exp_40_ram[1323] = 18;
    exp_40_ram[1324] = 18;
    exp_40_ram[1325] = 18;
    exp_40_ram[1326] = 18;
    exp_40_ram[1327] = 18;
    exp_40_ram[1328] = 18;
    exp_40_ram[1329] = 18;
    exp_40_ram[1330] = 18;
    exp_40_ram[1331] = 18;
    exp_40_ram[1332] = 18;
    exp_40_ram[1333] = 18;
    exp_40_ram[1334] = 18;
    exp_40_ram[1335] = 18;
    exp_40_ram[1336] = 18;
    exp_40_ram[1337] = 18;
    exp_40_ram[1338] = 18;
    exp_40_ram[1339] = 18;
    exp_40_ram[1340] = 18;
    exp_40_ram[1341] = 18;
    exp_40_ram[1342] = 18;
    exp_40_ram[1343] = 18;
    exp_40_ram[1344] = 12;
    exp_40_ram[1345] = 18;
    exp_40_ram[1346] = 18;
    exp_40_ram[1347] = 18;
    exp_40_ram[1348] = 18;
    exp_40_ram[1349] = 18;
    exp_40_ram[1350] = 18;
    exp_40_ram[1351] = 18;
    exp_40_ram[1352] = 18;
    exp_40_ram[1353] = 18;
    exp_40_ram[1354] = 12;
    exp_40_ram[1355] = 15;
    exp_40_ram[1356] = 12;
    exp_40_ram[1357] = 18;
    exp_40_ram[1358] = 18;
    exp_40_ram[1359] = 18;
    exp_40_ram[1360] = 18;
    exp_40_ram[1361] = 12;
    exp_40_ram[1362] = 18;
    exp_40_ram[1363] = 18;
    exp_40_ram[1364] = 18;
    exp_40_ram[1365] = 18;
    exp_40_ram[1366] = 18;
    exp_40_ram[1367] = 12;
    exp_40_ram[1368] = 17;
    exp_40_ram[1369] = 18;
    exp_40_ram[1370] = 18;
    exp_40_ram[1371] = 16;
    exp_40_ram[1372] = 18;
    exp_40_ram[1373] = 12;
    exp_40_ram[1374] = 18;
    exp_40_ram[1375] = 18;
    exp_40_ram[1376] = 12;
    exp_40_ram[1377] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [2047:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 55;
    exp_33_ram[32] = 19;
    exp_33_ram[33] = 239;
    exp_33_ram[34] = 111;
    exp_33_ram[35] = 72;
    exp_33_ram[36] = 111;
    exp_33_ram[37] = 114;
    exp_33_ram[38] = 10;
    exp_33_ram[39] = 19;
    exp_33_ram[40] = 35;
    exp_33_ram[41] = 19;
    exp_33_ram[42] = 35;
    exp_33_ram[43] = 35;
    exp_33_ram[44] = 131;
    exp_33_ram[45] = 35;
    exp_33_ram[46] = 3;
    exp_33_ram[47] = 131;
    exp_33_ram[48] = 35;
    exp_33_ram[49] = 131;
    exp_33_ram[50] = 19;
    exp_33_ram[51] = 3;
    exp_33_ram[52] = 19;
    exp_33_ram[53] = 103;
    exp_33_ram[54] = 19;
    exp_33_ram[55] = 35;
    exp_33_ram[56] = 19;
    exp_33_ram[57] = 147;
    exp_33_ram[58] = 35;
    exp_33_ram[59] = 35;
    exp_33_ram[60] = 35;
    exp_33_ram[61] = 163;
    exp_33_ram[62] = 19;
    exp_33_ram[63] = 3;
    exp_33_ram[64] = 19;
    exp_33_ram[65] = 103;
    exp_33_ram[66] = 19;
    exp_33_ram[67] = 35;
    exp_33_ram[68] = 35;
    exp_33_ram[69] = 19;
    exp_33_ram[70] = 147;
    exp_33_ram[71] = 35;
    exp_33_ram[72] = 35;
    exp_33_ram[73] = 35;
    exp_33_ram[74] = 163;
    exp_33_ram[75] = 131;
    exp_33_ram[76] = 99;
    exp_33_ram[77] = 131;
    exp_33_ram[78] = 19;
    exp_33_ram[79] = 239;
    exp_33_ram[80] = 19;
    exp_33_ram[81] = 131;
    exp_33_ram[82] = 3;
    exp_33_ram[83] = 19;
    exp_33_ram[84] = 103;
    exp_33_ram[85] = 19;
    exp_33_ram[86] = 35;
    exp_33_ram[87] = 19;
    exp_33_ram[88] = 35;
    exp_33_ram[89] = 35;
    exp_33_ram[90] = 131;
    exp_33_ram[91] = 35;
    exp_33_ram[92] = 111;
    exp_33_ram[93] = 131;
    exp_33_ram[94] = 147;
    exp_33_ram[95] = 35;
    exp_33_ram[96] = 131;
    exp_33_ram[97] = 131;
    exp_33_ram[98] = 99;
    exp_33_ram[99] = 131;
    exp_33_ram[100] = 19;
    exp_33_ram[101] = 35;
    exp_33_ram[102] = 227;
    exp_33_ram[103] = 3;
    exp_33_ram[104] = 131;
    exp_33_ram[105] = 179;
    exp_33_ram[106] = 19;
    exp_33_ram[107] = 3;
    exp_33_ram[108] = 19;
    exp_33_ram[109] = 103;
    exp_33_ram[110] = 19;
    exp_33_ram[111] = 35;
    exp_33_ram[112] = 19;
    exp_33_ram[113] = 147;
    exp_33_ram[114] = 163;
    exp_33_ram[115] = 3;
    exp_33_ram[116] = 147;
    exp_33_ram[117] = 99;
    exp_33_ram[118] = 3;
    exp_33_ram[119] = 147;
    exp_33_ram[120] = 99;
    exp_33_ram[121] = 147;
    exp_33_ram[122] = 111;
    exp_33_ram[123] = 147;
    exp_33_ram[124] = 147;
    exp_33_ram[125] = 147;
    exp_33_ram[126] = 19;
    exp_33_ram[127] = 3;
    exp_33_ram[128] = 19;
    exp_33_ram[129] = 103;
    exp_33_ram[130] = 19;
    exp_33_ram[131] = 35;
    exp_33_ram[132] = 35;
    exp_33_ram[133] = 19;
    exp_33_ram[134] = 35;
    exp_33_ram[135] = 35;
    exp_33_ram[136] = 111;
    exp_33_ram[137] = 3;
    exp_33_ram[138] = 147;
    exp_33_ram[139] = 147;
    exp_33_ram[140] = 179;
    exp_33_ram[141] = 147;
    exp_33_ram[142] = 19;
    exp_33_ram[143] = 131;
    exp_33_ram[144] = 131;
    exp_33_ram[145] = 147;
    exp_33_ram[146] = 3;
    exp_33_ram[147] = 35;
    exp_33_ram[148] = 131;
    exp_33_ram[149] = 179;
    exp_33_ram[150] = 147;
    exp_33_ram[151] = 35;
    exp_33_ram[152] = 131;
    exp_33_ram[153] = 131;
    exp_33_ram[154] = 131;
    exp_33_ram[155] = 19;
    exp_33_ram[156] = 239;
    exp_33_ram[157] = 147;
    exp_33_ram[158] = 227;
    exp_33_ram[159] = 131;
    exp_33_ram[160] = 19;
    exp_33_ram[161] = 131;
    exp_33_ram[162] = 3;
    exp_33_ram[163] = 19;
    exp_33_ram[164] = 103;
    exp_33_ram[165] = 19;
    exp_33_ram[166] = 35;
    exp_33_ram[167] = 35;
    exp_33_ram[168] = 19;
    exp_33_ram[169] = 35;
    exp_33_ram[170] = 35;
    exp_33_ram[171] = 35;
    exp_33_ram[172] = 35;
    exp_33_ram[173] = 35;
    exp_33_ram[174] = 35;
    exp_33_ram[175] = 35;
    exp_33_ram[176] = 35;
    exp_33_ram[177] = 131;
    exp_33_ram[178] = 35;
    exp_33_ram[179] = 131;
    exp_33_ram[180] = 147;
    exp_33_ram[181] = 99;
    exp_33_ram[182] = 131;
    exp_33_ram[183] = 147;
    exp_33_ram[184] = 99;
    exp_33_ram[185] = 131;
    exp_33_ram[186] = 35;
    exp_33_ram[187] = 111;
    exp_33_ram[188] = 131;
    exp_33_ram[189] = 19;
    exp_33_ram[190] = 35;
    exp_33_ram[191] = 3;
    exp_33_ram[192] = 131;
    exp_33_ram[193] = 19;
    exp_33_ram[194] = 131;
    exp_33_ram[195] = 19;
    exp_33_ram[196] = 231;
    exp_33_ram[197] = 131;
    exp_33_ram[198] = 147;
    exp_33_ram[199] = 35;
    exp_33_ram[200] = 3;
    exp_33_ram[201] = 131;
    exp_33_ram[202] = 227;
    exp_33_ram[203] = 111;
    exp_33_ram[204] = 131;
    exp_33_ram[205] = 147;
    exp_33_ram[206] = 35;
    exp_33_ram[207] = 3;
    exp_33_ram[208] = 131;
    exp_33_ram[209] = 179;
    exp_33_ram[210] = 3;
    exp_33_ram[211] = 131;
    exp_33_ram[212] = 19;
    exp_33_ram[213] = 35;
    exp_33_ram[214] = 3;
    exp_33_ram[215] = 131;
    exp_33_ram[216] = 19;
    exp_33_ram[217] = 131;
    exp_33_ram[218] = 231;
    exp_33_ram[219] = 131;
    exp_33_ram[220] = 227;
    exp_33_ram[221] = 131;
    exp_33_ram[222] = 147;
    exp_33_ram[223] = 99;
    exp_33_ram[224] = 111;
    exp_33_ram[225] = 131;
    exp_33_ram[226] = 19;
    exp_33_ram[227] = 35;
    exp_33_ram[228] = 3;
    exp_33_ram[229] = 131;
    exp_33_ram[230] = 19;
    exp_33_ram[231] = 131;
    exp_33_ram[232] = 19;
    exp_33_ram[233] = 231;
    exp_33_ram[234] = 3;
    exp_33_ram[235] = 131;
    exp_33_ram[236] = 179;
    exp_33_ram[237] = 3;
    exp_33_ram[238] = 227;
    exp_33_ram[239] = 131;
    exp_33_ram[240] = 19;
    exp_33_ram[241] = 131;
    exp_33_ram[242] = 3;
    exp_33_ram[243] = 19;
    exp_33_ram[244] = 103;
    exp_33_ram[245] = 19;
    exp_33_ram[246] = 35;
    exp_33_ram[247] = 35;
    exp_33_ram[248] = 19;
    exp_33_ram[249] = 35;
    exp_33_ram[250] = 35;
    exp_33_ram[251] = 35;
    exp_33_ram[252] = 35;
    exp_33_ram[253] = 35;
    exp_33_ram[254] = 35;
    exp_33_ram[255] = 147;
    exp_33_ram[256] = 35;
    exp_33_ram[257] = 163;
    exp_33_ram[258] = 131;
    exp_33_ram[259] = 147;
    exp_33_ram[260] = 99;
    exp_33_ram[261] = 131;
    exp_33_ram[262] = 99;
    exp_33_ram[263] = 131;
    exp_33_ram[264] = 147;
    exp_33_ram[265] = 99;
    exp_33_ram[266] = 131;
    exp_33_ram[267] = 99;
    exp_33_ram[268] = 131;
    exp_33_ram[269] = 147;
    exp_33_ram[270] = 99;
    exp_33_ram[271] = 131;
    exp_33_ram[272] = 147;
    exp_33_ram[273] = 35;
    exp_33_ram[274] = 111;
    exp_33_ram[275] = 131;
    exp_33_ram[276] = 19;
    exp_33_ram[277] = 35;
    exp_33_ram[278] = 3;
    exp_33_ram[279] = 179;
    exp_33_ram[280] = 19;
    exp_33_ram[281] = 35;
    exp_33_ram[282] = 3;
    exp_33_ram[283] = 131;
    exp_33_ram[284] = 99;
    exp_33_ram[285] = 3;
    exp_33_ram[286] = 147;
    exp_33_ram[287] = 227;
    exp_33_ram[288] = 111;
    exp_33_ram[289] = 131;
    exp_33_ram[290] = 19;
    exp_33_ram[291] = 35;
    exp_33_ram[292] = 3;
    exp_33_ram[293] = 179;
    exp_33_ram[294] = 19;
    exp_33_ram[295] = 35;
    exp_33_ram[296] = 131;
    exp_33_ram[297] = 147;
    exp_33_ram[298] = 99;
    exp_33_ram[299] = 3;
    exp_33_ram[300] = 131;
    exp_33_ram[301] = 99;
    exp_33_ram[302] = 3;
    exp_33_ram[303] = 147;
    exp_33_ram[304] = 227;
    exp_33_ram[305] = 131;
    exp_33_ram[306] = 147;
    exp_33_ram[307] = 99;
    exp_33_ram[308] = 131;
    exp_33_ram[309] = 147;
    exp_33_ram[310] = 99;
    exp_33_ram[311] = 131;
    exp_33_ram[312] = 99;
    exp_33_ram[313] = 3;
    exp_33_ram[314] = 131;
    exp_33_ram[315] = 99;
    exp_33_ram[316] = 3;
    exp_33_ram[317] = 131;
    exp_33_ram[318] = 99;
    exp_33_ram[319] = 131;
    exp_33_ram[320] = 147;
    exp_33_ram[321] = 35;
    exp_33_ram[322] = 131;
    exp_33_ram[323] = 99;
    exp_33_ram[324] = 3;
    exp_33_ram[325] = 147;
    exp_33_ram[326] = 99;
    exp_33_ram[327] = 131;
    exp_33_ram[328] = 147;
    exp_33_ram[329] = 35;
    exp_33_ram[330] = 3;
    exp_33_ram[331] = 147;
    exp_33_ram[332] = 99;
    exp_33_ram[333] = 131;
    exp_33_ram[334] = 147;
    exp_33_ram[335] = 99;
    exp_33_ram[336] = 3;
    exp_33_ram[337] = 147;
    exp_33_ram[338] = 99;
    exp_33_ram[339] = 131;
    exp_33_ram[340] = 19;
    exp_33_ram[341] = 35;
    exp_33_ram[342] = 3;
    exp_33_ram[343] = 179;
    exp_33_ram[344] = 19;
    exp_33_ram[345] = 35;
    exp_33_ram[346] = 111;
    exp_33_ram[347] = 3;
    exp_33_ram[348] = 147;
    exp_33_ram[349] = 99;
    exp_33_ram[350] = 131;
    exp_33_ram[351] = 147;
    exp_33_ram[352] = 99;
    exp_33_ram[353] = 3;
    exp_33_ram[354] = 147;
    exp_33_ram[355] = 99;
    exp_33_ram[356] = 131;
    exp_33_ram[357] = 19;
    exp_33_ram[358] = 35;
    exp_33_ram[359] = 3;
    exp_33_ram[360] = 179;
    exp_33_ram[361] = 19;
    exp_33_ram[362] = 35;
    exp_33_ram[363] = 111;
    exp_33_ram[364] = 3;
    exp_33_ram[365] = 147;
    exp_33_ram[366] = 99;
    exp_33_ram[367] = 3;
    exp_33_ram[368] = 147;
    exp_33_ram[369] = 99;
    exp_33_ram[370] = 131;
    exp_33_ram[371] = 19;
    exp_33_ram[372] = 35;
    exp_33_ram[373] = 3;
    exp_33_ram[374] = 179;
    exp_33_ram[375] = 19;
    exp_33_ram[376] = 35;
    exp_33_ram[377] = 3;
    exp_33_ram[378] = 147;
    exp_33_ram[379] = 99;
    exp_33_ram[380] = 131;
    exp_33_ram[381] = 19;
    exp_33_ram[382] = 35;
    exp_33_ram[383] = 3;
    exp_33_ram[384] = 179;
    exp_33_ram[385] = 19;
    exp_33_ram[386] = 35;
    exp_33_ram[387] = 3;
    exp_33_ram[388] = 147;
    exp_33_ram[389] = 99;
    exp_33_ram[390] = 131;
    exp_33_ram[391] = 99;
    exp_33_ram[392] = 131;
    exp_33_ram[393] = 19;
    exp_33_ram[394] = 35;
    exp_33_ram[395] = 3;
    exp_33_ram[396] = 179;
    exp_33_ram[397] = 19;
    exp_33_ram[398] = 35;
    exp_33_ram[399] = 111;
    exp_33_ram[400] = 131;
    exp_33_ram[401] = 147;
    exp_33_ram[402] = 99;
    exp_33_ram[403] = 131;
    exp_33_ram[404] = 19;
    exp_33_ram[405] = 35;
    exp_33_ram[406] = 3;
    exp_33_ram[407] = 179;
    exp_33_ram[408] = 19;
    exp_33_ram[409] = 35;
    exp_33_ram[410] = 111;
    exp_33_ram[411] = 131;
    exp_33_ram[412] = 147;
    exp_33_ram[413] = 99;
    exp_33_ram[414] = 131;
    exp_33_ram[415] = 19;
    exp_33_ram[416] = 35;
    exp_33_ram[417] = 3;
    exp_33_ram[418] = 179;
    exp_33_ram[419] = 19;
    exp_33_ram[420] = 35;
    exp_33_ram[421] = 131;
    exp_33_ram[422] = 3;
    exp_33_ram[423] = 131;
    exp_33_ram[424] = 3;
    exp_33_ram[425] = 131;
    exp_33_ram[426] = 3;
    exp_33_ram[427] = 131;
    exp_33_ram[428] = 3;
    exp_33_ram[429] = 239;
    exp_33_ram[430] = 147;
    exp_33_ram[431] = 19;
    exp_33_ram[432] = 131;
    exp_33_ram[433] = 3;
    exp_33_ram[434] = 19;
    exp_33_ram[435] = 103;
    exp_33_ram[436] = 19;
    exp_33_ram[437] = 35;
    exp_33_ram[438] = 35;
    exp_33_ram[439] = 19;
    exp_33_ram[440] = 35;
    exp_33_ram[441] = 35;
    exp_33_ram[442] = 35;
    exp_33_ram[443] = 35;
    exp_33_ram[444] = 35;
    exp_33_ram[445] = 35;
    exp_33_ram[446] = 35;
    exp_33_ram[447] = 163;
    exp_33_ram[448] = 35;
    exp_33_ram[449] = 131;
    exp_33_ram[450] = 99;
    exp_33_ram[451] = 131;
    exp_33_ram[452] = 147;
    exp_33_ram[453] = 35;
    exp_33_ram[454] = 131;
    exp_33_ram[455] = 147;
    exp_33_ram[456] = 99;
    exp_33_ram[457] = 131;
    exp_33_ram[458] = 99;
    exp_33_ram[459] = 3;
    exp_33_ram[460] = 131;
    exp_33_ram[461] = 179;
    exp_33_ram[462] = 163;
    exp_33_ram[463] = 3;
    exp_33_ram[464] = 147;
    exp_33_ram[465] = 99;
    exp_33_ram[466] = 131;
    exp_33_ram[467] = 147;
    exp_33_ram[468] = 147;
    exp_33_ram[469] = 111;
    exp_33_ram[470] = 131;
    exp_33_ram[471] = 147;
    exp_33_ram[472] = 99;
    exp_33_ram[473] = 147;
    exp_33_ram[474] = 111;
    exp_33_ram[475] = 147;
    exp_33_ram[476] = 3;
    exp_33_ram[477] = 179;
    exp_33_ram[478] = 147;
    exp_33_ram[479] = 147;
    exp_33_ram[480] = 147;
    exp_33_ram[481] = 3;
    exp_33_ram[482] = 147;
    exp_33_ram[483] = 35;
    exp_33_ram[484] = 147;
    exp_33_ram[485] = 51;
    exp_33_ram[486] = 35;
    exp_33_ram[487] = 3;
    exp_33_ram[488] = 131;
    exp_33_ram[489] = 179;
    exp_33_ram[490] = 35;
    exp_33_ram[491] = 131;
    exp_33_ram[492] = 99;
    exp_33_ram[493] = 3;
    exp_33_ram[494] = 147;
    exp_33_ram[495] = 227;
    exp_33_ram[496] = 131;
    exp_33_ram[497] = 19;
    exp_33_ram[498] = 131;
    exp_33_ram[499] = 35;
    exp_33_ram[500] = 131;
    exp_33_ram[501] = 35;
    exp_33_ram[502] = 131;
    exp_33_ram[503] = 35;
    exp_33_ram[504] = 131;
    exp_33_ram[505] = 19;
    exp_33_ram[506] = 131;
    exp_33_ram[507] = 131;
    exp_33_ram[508] = 3;
    exp_33_ram[509] = 131;
    exp_33_ram[510] = 3;
    exp_33_ram[511] = 239;
    exp_33_ram[512] = 147;
    exp_33_ram[513] = 19;
    exp_33_ram[514] = 131;
    exp_33_ram[515] = 3;
    exp_33_ram[516] = 19;
    exp_33_ram[517] = 103;
    exp_33_ram[518] = 19;
    exp_33_ram[519] = 35;
    exp_33_ram[520] = 35;
    exp_33_ram[521] = 19;
    exp_33_ram[522] = 35;
    exp_33_ram[523] = 35;
    exp_33_ram[524] = 35;
    exp_33_ram[525] = 35;
    exp_33_ram[526] = 35;
    exp_33_ram[527] = 35;
    exp_33_ram[528] = 131;
    exp_33_ram[529] = 227;
    exp_33_ram[530] = 147;
    exp_33_ram[531] = 35;
    exp_33_ram[532] = 111;
    exp_33_ram[533] = 131;
    exp_33_ram[534] = 3;
    exp_33_ram[535] = 147;
    exp_33_ram[536] = 99;
    exp_33_ram[537] = 131;
    exp_33_ram[538] = 3;
    exp_33_ram[539] = 131;
    exp_33_ram[540] = 19;
    exp_33_ram[541] = 35;
    exp_33_ram[542] = 3;
    exp_33_ram[543] = 131;
    exp_33_ram[544] = 19;
    exp_33_ram[545] = 131;
    exp_33_ram[546] = 231;
    exp_33_ram[547] = 131;
    exp_33_ram[548] = 147;
    exp_33_ram[549] = 35;
    exp_33_ram[550] = 111;
    exp_33_ram[551] = 131;
    exp_33_ram[552] = 147;
    exp_33_ram[553] = 35;
    exp_33_ram[554] = 35;
    exp_33_ram[555] = 131;
    exp_33_ram[556] = 131;
    exp_33_ram[557] = 147;
    exp_33_ram[558] = 19;
    exp_33_ram[559] = 99;
    exp_33_ram[560] = 19;
    exp_33_ram[561] = 183;
    exp_33_ram[562] = 147;
    exp_33_ram[563] = 179;
    exp_33_ram[564] = 131;
    exp_33_ram[565] = 103;
    exp_33_ram[566] = 131;
    exp_33_ram[567] = 147;
    exp_33_ram[568] = 35;
    exp_33_ram[569] = 131;
    exp_33_ram[570] = 147;
    exp_33_ram[571] = 35;
    exp_33_ram[572] = 147;
    exp_33_ram[573] = 35;
    exp_33_ram[574] = 111;
    exp_33_ram[575] = 131;
    exp_33_ram[576] = 147;
    exp_33_ram[577] = 35;
    exp_33_ram[578] = 131;
    exp_33_ram[579] = 147;
    exp_33_ram[580] = 35;
    exp_33_ram[581] = 147;
    exp_33_ram[582] = 35;
    exp_33_ram[583] = 111;
    exp_33_ram[584] = 131;
    exp_33_ram[585] = 147;
    exp_33_ram[586] = 35;
    exp_33_ram[587] = 131;
    exp_33_ram[588] = 147;
    exp_33_ram[589] = 35;
    exp_33_ram[590] = 147;
    exp_33_ram[591] = 35;
    exp_33_ram[592] = 111;
    exp_33_ram[593] = 131;
    exp_33_ram[594] = 147;
    exp_33_ram[595] = 35;
    exp_33_ram[596] = 131;
    exp_33_ram[597] = 147;
    exp_33_ram[598] = 35;
    exp_33_ram[599] = 147;
    exp_33_ram[600] = 35;
    exp_33_ram[601] = 111;
    exp_33_ram[602] = 131;
    exp_33_ram[603] = 147;
    exp_33_ram[604] = 35;
    exp_33_ram[605] = 131;
    exp_33_ram[606] = 147;
    exp_33_ram[607] = 35;
    exp_33_ram[608] = 147;
    exp_33_ram[609] = 35;
    exp_33_ram[610] = 111;
    exp_33_ram[611] = 35;
    exp_33_ram[612] = 19;
    exp_33_ram[613] = 131;
    exp_33_ram[614] = 227;
    exp_33_ram[615] = 35;
    exp_33_ram[616] = 131;
    exp_33_ram[617] = 131;
    exp_33_ram[618] = 19;
    exp_33_ram[619] = 239;
    exp_33_ram[620] = 147;
    exp_33_ram[621] = 99;
    exp_33_ram[622] = 147;
    exp_33_ram[623] = 19;
    exp_33_ram[624] = 239;
    exp_33_ram[625] = 35;
    exp_33_ram[626] = 111;
    exp_33_ram[627] = 131;
    exp_33_ram[628] = 3;
    exp_33_ram[629] = 147;
    exp_33_ram[630] = 99;
    exp_33_ram[631] = 131;
    exp_33_ram[632] = 19;
    exp_33_ram[633] = 35;
    exp_33_ram[634] = 131;
    exp_33_ram[635] = 35;
    exp_33_ram[636] = 131;
    exp_33_ram[637] = 99;
    exp_33_ram[638] = 131;
    exp_33_ram[639] = 147;
    exp_33_ram[640] = 35;
    exp_33_ram[641] = 131;
    exp_33_ram[642] = 179;
    exp_33_ram[643] = 35;
    exp_33_ram[644] = 111;
    exp_33_ram[645] = 131;
    exp_33_ram[646] = 35;
    exp_33_ram[647] = 131;
    exp_33_ram[648] = 147;
    exp_33_ram[649] = 35;
    exp_33_ram[650] = 35;
    exp_33_ram[651] = 131;
    exp_33_ram[652] = 3;
    exp_33_ram[653] = 147;
    exp_33_ram[654] = 99;
    exp_33_ram[655] = 131;
    exp_33_ram[656] = 147;
    exp_33_ram[657] = 35;
    exp_33_ram[658] = 131;
    exp_33_ram[659] = 147;
    exp_33_ram[660] = 35;
    exp_33_ram[661] = 131;
    exp_33_ram[662] = 131;
    exp_33_ram[663] = 19;
    exp_33_ram[664] = 239;
    exp_33_ram[665] = 147;
    exp_33_ram[666] = 99;
    exp_33_ram[667] = 147;
    exp_33_ram[668] = 19;
    exp_33_ram[669] = 239;
    exp_33_ram[670] = 35;
    exp_33_ram[671] = 111;
    exp_33_ram[672] = 131;
    exp_33_ram[673] = 3;
    exp_33_ram[674] = 147;
    exp_33_ram[675] = 99;
    exp_33_ram[676] = 131;
    exp_33_ram[677] = 19;
    exp_33_ram[678] = 35;
    exp_33_ram[679] = 131;
    exp_33_ram[680] = 35;
    exp_33_ram[681] = 131;
    exp_33_ram[682] = 99;
    exp_33_ram[683] = 147;
    exp_33_ram[684] = 35;
    exp_33_ram[685] = 131;
    exp_33_ram[686] = 147;
    exp_33_ram[687] = 35;
    exp_33_ram[688] = 131;
    exp_33_ram[689] = 131;
    exp_33_ram[690] = 147;
    exp_33_ram[691] = 19;
    exp_33_ram[692] = 99;
    exp_33_ram[693] = 19;
    exp_33_ram[694] = 183;
    exp_33_ram[695] = 147;
    exp_33_ram[696] = 179;
    exp_33_ram[697] = 131;
    exp_33_ram[698] = 103;
    exp_33_ram[699] = 131;
    exp_33_ram[700] = 147;
    exp_33_ram[701] = 35;
    exp_33_ram[702] = 131;
    exp_33_ram[703] = 147;
    exp_33_ram[704] = 35;
    exp_33_ram[705] = 131;
    exp_33_ram[706] = 3;
    exp_33_ram[707] = 147;
    exp_33_ram[708] = 99;
    exp_33_ram[709] = 131;
    exp_33_ram[710] = 147;
    exp_33_ram[711] = 35;
    exp_33_ram[712] = 131;
    exp_33_ram[713] = 147;
    exp_33_ram[714] = 35;
    exp_33_ram[715] = 111;
    exp_33_ram[716] = 131;
    exp_33_ram[717] = 147;
    exp_33_ram[718] = 35;
    exp_33_ram[719] = 131;
    exp_33_ram[720] = 147;
    exp_33_ram[721] = 35;
    exp_33_ram[722] = 131;
    exp_33_ram[723] = 3;
    exp_33_ram[724] = 147;
    exp_33_ram[725] = 99;
    exp_33_ram[726] = 131;
    exp_33_ram[727] = 147;
    exp_33_ram[728] = 35;
    exp_33_ram[729] = 131;
    exp_33_ram[730] = 147;
    exp_33_ram[731] = 35;
    exp_33_ram[732] = 111;
    exp_33_ram[733] = 131;
    exp_33_ram[734] = 147;
    exp_33_ram[735] = 35;
    exp_33_ram[736] = 131;
    exp_33_ram[737] = 147;
    exp_33_ram[738] = 35;
    exp_33_ram[739] = 111;
    exp_33_ram[740] = 131;
    exp_33_ram[741] = 147;
    exp_33_ram[742] = 35;
    exp_33_ram[743] = 131;
    exp_33_ram[744] = 147;
    exp_33_ram[745] = 35;
    exp_33_ram[746] = 111;
    exp_33_ram[747] = 131;
    exp_33_ram[748] = 147;
    exp_33_ram[749] = 35;
    exp_33_ram[750] = 131;
    exp_33_ram[751] = 147;
    exp_33_ram[752] = 35;
    exp_33_ram[753] = 111;
    exp_33_ram[754] = 19;
    exp_33_ram[755] = 111;
    exp_33_ram[756] = 19;
    exp_33_ram[757] = 111;
    exp_33_ram[758] = 19;
    exp_33_ram[759] = 131;
    exp_33_ram[760] = 131;
    exp_33_ram[761] = 147;
    exp_33_ram[762] = 19;
    exp_33_ram[763] = 99;
    exp_33_ram[764] = 19;
    exp_33_ram[765] = 183;
    exp_33_ram[766] = 147;
    exp_33_ram[767] = 179;
    exp_33_ram[768] = 131;
    exp_33_ram[769] = 103;
    exp_33_ram[770] = 131;
    exp_33_ram[771] = 3;
    exp_33_ram[772] = 147;
    exp_33_ram[773] = 99;
    exp_33_ram[774] = 131;
    exp_33_ram[775] = 3;
    exp_33_ram[776] = 147;
    exp_33_ram[777] = 99;
    exp_33_ram[778] = 147;
    exp_33_ram[779] = 35;
    exp_33_ram[780] = 111;
    exp_33_ram[781] = 131;
    exp_33_ram[782] = 3;
    exp_33_ram[783] = 147;
    exp_33_ram[784] = 99;
    exp_33_ram[785] = 147;
    exp_33_ram[786] = 35;
    exp_33_ram[787] = 111;
    exp_33_ram[788] = 131;
    exp_33_ram[789] = 3;
    exp_33_ram[790] = 147;
    exp_33_ram[791] = 99;
    exp_33_ram[792] = 147;
    exp_33_ram[793] = 35;
    exp_33_ram[794] = 111;
    exp_33_ram[795] = 147;
    exp_33_ram[796] = 35;
    exp_33_ram[797] = 131;
    exp_33_ram[798] = 147;
    exp_33_ram[799] = 35;
    exp_33_ram[800] = 131;
    exp_33_ram[801] = 3;
    exp_33_ram[802] = 147;
    exp_33_ram[803] = 99;
    exp_33_ram[804] = 131;
    exp_33_ram[805] = 147;
    exp_33_ram[806] = 35;
    exp_33_ram[807] = 131;
    exp_33_ram[808] = 3;
    exp_33_ram[809] = 147;
    exp_33_ram[810] = 99;
    exp_33_ram[811] = 131;
    exp_33_ram[812] = 3;
    exp_33_ram[813] = 147;
    exp_33_ram[814] = 99;
    exp_33_ram[815] = 131;
    exp_33_ram[816] = 147;
    exp_33_ram[817] = 35;
    exp_33_ram[818] = 131;
    exp_33_ram[819] = 147;
    exp_33_ram[820] = 99;
    exp_33_ram[821] = 131;
    exp_33_ram[822] = 147;
    exp_33_ram[823] = 35;
    exp_33_ram[824] = 131;
    exp_33_ram[825] = 3;
    exp_33_ram[826] = 147;
    exp_33_ram[827] = 99;
    exp_33_ram[828] = 131;
    exp_33_ram[829] = 3;
    exp_33_ram[830] = 147;
    exp_33_ram[831] = 99;
    exp_33_ram[832] = 131;
    exp_33_ram[833] = 147;
    exp_33_ram[834] = 99;
    exp_33_ram[835] = 131;
    exp_33_ram[836] = 147;
    exp_33_ram[837] = 99;
    exp_33_ram[838] = 131;
    exp_33_ram[839] = 19;
    exp_33_ram[840] = 35;
    exp_33_ram[841] = 131;
    exp_33_ram[842] = 35;
    exp_33_ram[843] = 131;
    exp_33_ram[844] = 19;
    exp_33_ram[845] = 131;
    exp_33_ram[846] = 179;
    exp_33_ram[847] = 179;
    exp_33_ram[848] = 147;
    exp_33_ram[849] = 131;
    exp_33_ram[850] = 147;
    exp_33_ram[851] = 19;
    exp_33_ram[852] = 131;
    exp_33_ram[853] = 35;
    exp_33_ram[854] = 131;
    exp_33_ram[855] = 35;
    exp_33_ram[856] = 131;
    exp_33_ram[857] = 3;
    exp_33_ram[858] = 147;
    exp_33_ram[859] = 19;
    exp_33_ram[860] = 131;
    exp_33_ram[861] = 3;
    exp_33_ram[862] = 131;
    exp_33_ram[863] = 3;
    exp_33_ram[864] = 239;
    exp_33_ram[865] = 35;
    exp_33_ram[866] = 111;
    exp_33_ram[867] = 131;
    exp_33_ram[868] = 147;
    exp_33_ram[869] = 99;
    exp_33_ram[870] = 131;
    exp_33_ram[871] = 19;
    exp_33_ram[872] = 35;
    exp_33_ram[873] = 131;
    exp_33_ram[874] = 147;
    exp_33_ram[875] = 111;
    exp_33_ram[876] = 131;
    exp_33_ram[877] = 147;
    exp_33_ram[878] = 99;
    exp_33_ram[879] = 131;
    exp_33_ram[880] = 19;
    exp_33_ram[881] = 35;
    exp_33_ram[882] = 131;
    exp_33_ram[883] = 147;
    exp_33_ram[884] = 147;
    exp_33_ram[885] = 111;
    exp_33_ram[886] = 131;
    exp_33_ram[887] = 19;
    exp_33_ram[888] = 35;
    exp_33_ram[889] = 131;
    exp_33_ram[890] = 35;
    exp_33_ram[891] = 131;
    exp_33_ram[892] = 19;
    exp_33_ram[893] = 131;
    exp_33_ram[894] = 179;
    exp_33_ram[895] = 179;
    exp_33_ram[896] = 147;
    exp_33_ram[897] = 131;
    exp_33_ram[898] = 147;
    exp_33_ram[899] = 19;
    exp_33_ram[900] = 131;
    exp_33_ram[901] = 35;
    exp_33_ram[902] = 131;
    exp_33_ram[903] = 35;
    exp_33_ram[904] = 131;
    exp_33_ram[905] = 3;
    exp_33_ram[906] = 147;
    exp_33_ram[907] = 19;
    exp_33_ram[908] = 131;
    exp_33_ram[909] = 3;
    exp_33_ram[910] = 131;
    exp_33_ram[911] = 3;
    exp_33_ram[912] = 239;
    exp_33_ram[913] = 35;
    exp_33_ram[914] = 111;
    exp_33_ram[915] = 131;
    exp_33_ram[916] = 147;
    exp_33_ram[917] = 99;
    exp_33_ram[918] = 131;
    exp_33_ram[919] = 147;
    exp_33_ram[920] = 99;
    exp_33_ram[921] = 131;
    exp_33_ram[922] = 19;
    exp_33_ram[923] = 35;
    exp_33_ram[924] = 3;
    exp_33_ram[925] = 131;
    exp_33_ram[926] = 35;
    exp_33_ram[927] = 131;
    exp_33_ram[928] = 35;
    exp_33_ram[929] = 131;
    exp_33_ram[930] = 3;
    exp_33_ram[931] = 147;
    exp_33_ram[932] = 131;
    exp_33_ram[933] = 3;
    exp_33_ram[934] = 131;
    exp_33_ram[935] = 3;
    exp_33_ram[936] = 239;
    exp_33_ram[937] = 35;
    exp_33_ram[938] = 111;
    exp_33_ram[939] = 131;
    exp_33_ram[940] = 147;
    exp_33_ram[941] = 99;
    exp_33_ram[942] = 131;
    exp_33_ram[943] = 19;
    exp_33_ram[944] = 35;
    exp_33_ram[945] = 131;
    exp_33_ram[946] = 147;
    exp_33_ram[947] = 111;
    exp_33_ram[948] = 131;
    exp_33_ram[949] = 147;
    exp_33_ram[950] = 99;
    exp_33_ram[951] = 131;
    exp_33_ram[952] = 19;
    exp_33_ram[953] = 35;
    exp_33_ram[954] = 131;
    exp_33_ram[955] = 147;
    exp_33_ram[956] = 147;
    exp_33_ram[957] = 111;
    exp_33_ram[958] = 131;
    exp_33_ram[959] = 19;
    exp_33_ram[960] = 35;
    exp_33_ram[961] = 131;
    exp_33_ram[962] = 35;
    exp_33_ram[963] = 131;
    exp_33_ram[964] = 35;
    exp_33_ram[965] = 131;
    exp_33_ram[966] = 35;
    exp_33_ram[967] = 131;
    exp_33_ram[968] = 3;
    exp_33_ram[969] = 147;
    exp_33_ram[970] = 3;
    exp_33_ram[971] = 131;
    exp_33_ram[972] = 3;
    exp_33_ram[973] = 131;
    exp_33_ram[974] = 3;
    exp_33_ram[975] = 239;
    exp_33_ram[976] = 35;
    exp_33_ram[977] = 131;
    exp_33_ram[978] = 147;
    exp_33_ram[979] = 35;
    exp_33_ram[980] = 111;
    exp_33_ram[981] = 147;
    exp_33_ram[982] = 35;
    exp_33_ram[983] = 131;
    exp_33_ram[984] = 147;
    exp_33_ram[985] = 99;
    exp_33_ram[986] = 111;
    exp_33_ram[987] = 131;
    exp_33_ram[988] = 19;
    exp_33_ram[989] = 35;
    exp_33_ram[990] = 3;
    exp_33_ram[991] = 131;
    exp_33_ram[992] = 19;
    exp_33_ram[993] = 131;
    exp_33_ram[994] = 19;
    exp_33_ram[995] = 231;
    exp_33_ram[996] = 131;
    exp_33_ram[997] = 19;
    exp_33_ram[998] = 35;
    exp_33_ram[999] = 3;
    exp_33_ram[1000] = 227;
    exp_33_ram[1001] = 131;
    exp_33_ram[1002] = 19;
    exp_33_ram[1003] = 35;
    exp_33_ram[1004] = 131;
    exp_33_ram[1005] = 19;
    exp_33_ram[1006] = 131;
    exp_33_ram[1007] = 19;
    exp_33_ram[1008] = 35;
    exp_33_ram[1009] = 3;
    exp_33_ram[1010] = 131;
    exp_33_ram[1011] = 19;
    exp_33_ram[1012] = 131;
    exp_33_ram[1013] = 231;
    exp_33_ram[1014] = 131;
    exp_33_ram[1015] = 147;
    exp_33_ram[1016] = 99;
    exp_33_ram[1017] = 111;
    exp_33_ram[1018] = 131;
    exp_33_ram[1019] = 19;
    exp_33_ram[1020] = 35;
    exp_33_ram[1021] = 3;
    exp_33_ram[1022] = 131;
    exp_33_ram[1023] = 19;
    exp_33_ram[1024] = 131;
    exp_33_ram[1025] = 19;
    exp_33_ram[1026] = 231;
    exp_33_ram[1027] = 131;
    exp_33_ram[1028] = 19;
    exp_33_ram[1029] = 35;
    exp_33_ram[1030] = 3;
    exp_33_ram[1031] = 227;
    exp_33_ram[1032] = 131;
    exp_33_ram[1033] = 147;
    exp_33_ram[1034] = 35;
    exp_33_ram[1035] = 111;
    exp_33_ram[1036] = 131;
    exp_33_ram[1037] = 19;
    exp_33_ram[1038] = 35;
    exp_33_ram[1039] = 131;
    exp_33_ram[1040] = 35;
    exp_33_ram[1041] = 131;
    exp_33_ram[1042] = 99;
    exp_33_ram[1043] = 131;
    exp_33_ram[1044] = 111;
    exp_33_ram[1045] = 147;
    exp_33_ram[1046] = 147;
    exp_33_ram[1047] = 3;
    exp_33_ram[1048] = 239;
    exp_33_ram[1049] = 35;
    exp_33_ram[1050] = 131;
    exp_33_ram[1051] = 147;
    exp_33_ram[1052] = 99;
    exp_33_ram[1053] = 3;
    exp_33_ram[1054] = 131;
    exp_33_ram[1055] = 99;
    exp_33_ram[1056] = 147;
    exp_33_ram[1057] = 35;
    exp_33_ram[1058] = 131;
    exp_33_ram[1059] = 147;
    exp_33_ram[1060] = 99;
    exp_33_ram[1061] = 111;
    exp_33_ram[1062] = 131;
    exp_33_ram[1063] = 19;
    exp_33_ram[1064] = 35;
    exp_33_ram[1065] = 3;
    exp_33_ram[1066] = 131;
    exp_33_ram[1067] = 19;
    exp_33_ram[1068] = 131;
    exp_33_ram[1069] = 19;
    exp_33_ram[1070] = 231;
    exp_33_ram[1071] = 131;
    exp_33_ram[1072] = 19;
    exp_33_ram[1073] = 35;
    exp_33_ram[1074] = 3;
    exp_33_ram[1075] = 227;
    exp_33_ram[1076] = 111;
    exp_33_ram[1077] = 131;
    exp_33_ram[1078] = 19;
    exp_33_ram[1079] = 35;
    exp_33_ram[1080] = 3;
    exp_33_ram[1081] = 131;
    exp_33_ram[1082] = 19;
    exp_33_ram[1083] = 35;
    exp_33_ram[1084] = 3;
    exp_33_ram[1085] = 131;
    exp_33_ram[1086] = 19;
    exp_33_ram[1087] = 131;
    exp_33_ram[1088] = 231;
    exp_33_ram[1089] = 131;
    exp_33_ram[1090] = 131;
    exp_33_ram[1091] = 99;
    exp_33_ram[1092] = 131;
    exp_33_ram[1093] = 147;
    exp_33_ram[1094] = 227;
    exp_33_ram[1095] = 131;
    exp_33_ram[1096] = 19;
    exp_33_ram[1097] = 35;
    exp_33_ram[1098] = 227;
    exp_33_ram[1099] = 131;
    exp_33_ram[1100] = 147;
    exp_33_ram[1101] = 99;
    exp_33_ram[1102] = 111;
    exp_33_ram[1103] = 131;
    exp_33_ram[1104] = 19;
    exp_33_ram[1105] = 35;
    exp_33_ram[1106] = 3;
    exp_33_ram[1107] = 131;
    exp_33_ram[1108] = 19;
    exp_33_ram[1109] = 131;
    exp_33_ram[1110] = 19;
    exp_33_ram[1111] = 231;
    exp_33_ram[1112] = 131;
    exp_33_ram[1113] = 19;
    exp_33_ram[1114] = 35;
    exp_33_ram[1115] = 3;
    exp_33_ram[1116] = 227;
    exp_33_ram[1117] = 131;
    exp_33_ram[1118] = 147;
    exp_33_ram[1119] = 35;
    exp_33_ram[1120] = 111;
    exp_33_ram[1121] = 147;
    exp_33_ram[1122] = 35;
    exp_33_ram[1123] = 131;
    exp_33_ram[1124] = 147;
    exp_33_ram[1125] = 35;
    exp_33_ram[1126] = 131;
    exp_33_ram[1127] = 19;
    exp_33_ram[1128] = 35;
    exp_33_ram[1129] = 131;
    exp_33_ram[1130] = 19;
    exp_33_ram[1131] = 131;
    exp_33_ram[1132] = 35;
    exp_33_ram[1133] = 131;
    exp_33_ram[1134] = 35;
    exp_33_ram[1135] = 131;
    exp_33_ram[1136] = 19;
    exp_33_ram[1137] = 147;
    exp_33_ram[1138] = 131;
    exp_33_ram[1139] = 3;
    exp_33_ram[1140] = 131;
    exp_33_ram[1141] = 3;
    exp_33_ram[1142] = 239;
    exp_33_ram[1143] = 35;
    exp_33_ram[1144] = 131;
    exp_33_ram[1145] = 147;
    exp_33_ram[1146] = 35;
    exp_33_ram[1147] = 111;
    exp_33_ram[1148] = 131;
    exp_33_ram[1149] = 19;
    exp_33_ram[1150] = 35;
    exp_33_ram[1151] = 3;
    exp_33_ram[1152] = 131;
    exp_33_ram[1153] = 19;
    exp_33_ram[1154] = 131;
    exp_33_ram[1155] = 19;
    exp_33_ram[1156] = 231;
    exp_33_ram[1157] = 131;
    exp_33_ram[1158] = 147;
    exp_33_ram[1159] = 35;
    exp_33_ram[1160] = 111;
    exp_33_ram[1161] = 131;
    exp_33_ram[1162] = 3;
    exp_33_ram[1163] = 131;
    exp_33_ram[1164] = 19;
    exp_33_ram[1165] = 35;
    exp_33_ram[1166] = 3;
    exp_33_ram[1167] = 131;
    exp_33_ram[1168] = 19;
    exp_33_ram[1169] = 131;
    exp_33_ram[1170] = 231;
    exp_33_ram[1171] = 131;
    exp_33_ram[1172] = 147;
    exp_33_ram[1173] = 35;
    exp_33_ram[1174] = 19;
    exp_33_ram[1175] = 131;
    exp_33_ram[1176] = 131;
    exp_33_ram[1177] = 99;
    exp_33_ram[1178] = 3;
    exp_33_ram[1179] = 131;
    exp_33_ram[1180] = 99;
    exp_33_ram[1181] = 131;
    exp_33_ram[1182] = 147;
    exp_33_ram[1183] = 111;
    exp_33_ram[1184] = 131;
    exp_33_ram[1185] = 3;
    exp_33_ram[1186] = 131;
    exp_33_ram[1187] = 19;
    exp_33_ram[1188] = 131;
    exp_33_ram[1189] = 19;
    exp_33_ram[1190] = 231;
    exp_33_ram[1191] = 131;
    exp_33_ram[1192] = 19;
    exp_33_ram[1193] = 131;
    exp_33_ram[1194] = 3;
    exp_33_ram[1195] = 19;
    exp_33_ram[1196] = 103;
    exp_33_ram[1197] = 19;
    exp_33_ram[1198] = 35;
    exp_33_ram[1199] = 35;
    exp_33_ram[1200] = 19;
    exp_33_ram[1201] = 35;
    exp_33_ram[1202] = 35;
    exp_33_ram[1203] = 35;
    exp_33_ram[1204] = 35;
    exp_33_ram[1205] = 35;
    exp_33_ram[1206] = 35;
    exp_33_ram[1207] = 35;
    exp_33_ram[1208] = 35;
    exp_33_ram[1209] = 147;
    exp_33_ram[1210] = 35;
    exp_33_ram[1211] = 131;
    exp_33_ram[1212] = 147;
    exp_33_ram[1213] = 35;
    exp_33_ram[1214] = 3;
    exp_33_ram[1215] = 147;
    exp_33_ram[1216] = 131;
    exp_33_ram[1217] = 19;
    exp_33_ram[1218] = 147;
    exp_33_ram[1219] = 19;
    exp_33_ram[1220] = 239;
    exp_33_ram[1221] = 35;
    exp_33_ram[1222] = 131;
    exp_33_ram[1223] = 19;
    exp_33_ram[1224] = 131;
    exp_33_ram[1225] = 3;
    exp_33_ram[1226] = 19;
    exp_33_ram[1227] = 103;
    exp_33_ram[1228] = 19;
    exp_33_ram[1229] = 35;
    exp_33_ram[1230] = 35;
    exp_33_ram[1231] = 19;
    exp_33_ram[1232] = 147;
    exp_33_ram[1233] = 163;
    exp_33_ram[1234] = 3;
    exp_33_ram[1235] = 183;
    exp_33_ram[1236] = 131;
    exp_33_ram[1237] = 147;
    exp_33_ram[1238] = 19;
    exp_33_ram[1239] = 239;
    exp_33_ram[1240] = 19;
    exp_33_ram[1241] = 131;
    exp_33_ram[1242] = 3;
    exp_33_ram[1243] = 19;
    exp_33_ram[1244] = 103;
    exp_33_ram[1245] = 19;
    exp_33_ram[1246] = 35;
    exp_33_ram[1247] = 35;
    exp_33_ram[1248] = 19;
    exp_33_ram[1249] = 19;
    exp_33_ram[1250] = 239;
    exp_33_ram[1251] = 19;
    exp_33_ram[1252] = 131;
    exp_33_ram[1253] = 3;
    exp_33_ram[1254] = 19;
    exp_33_ram[1255] = 103;
    exp_33_ram[1256] = 8;
    exp_33_ram[1257] = 68;
    exp_33_ram[1258] = 140;
    exp_33_ram[1259] = 140;
    exp_33_ram[1260] = 104;
    exp_33_ram[1261] = 140;
    exp_33_ram[1262] = 140;
    exp_33_ram[1263] = 140;
    exp_33_ram[1264] = 140;
    exp_33_ram[1265] = 140;
    exp_33_ram[1266] = 140;
    exp_33_ram[1267] = 140;
    exp_33_ram[1268] = 32;
    exp_33_ram[1269] = 140;
    exp_33_ram[1270] = 252;
    exp_33_ram[1271] = 140;
    exp_33_ram[1272] = 140;
    exp_33_ram[1273] = 216;
    exp_33_ram[1274] = 48;
    exp_33_ram[1275] = 200;
    exp_33_ram[1276] = 144;
    exp_33_ram[1277] = 200;
    exp_33_ram[1278] = 236;
    exp_33_ram[1279] = 200;
    exp_33_ram[1280] = 200;
    exp_33_ram[1281] = 200;
    exp_33_ram[1282] = 200;
    exp_33_ram[1283] = 200;
    exp_33_ram[1284] = 200;
    exp_33_ram[1285] = 200;
    exp_33_ram[1286] = 116;
    exp_33_ram[1287] = 200;
    exp_33_ram[1288] = 200;
    exp_33_ram[1289] = 200;
    exp_33_ram[1290] = 200;
    exp_33_ram[1291] = 200;
    exp_33_ram[1292] = 172;
    exp_33_ram[1293] = 240;
    exp_33_ram[1294] = 36;
    exp_33_ram[1295] = 36;
    exp_33_ram[1296] = 36;
    exp_33_ram[1297] = 36;
    exp_33_ram[1298] = 36;
    exp_33_ram[1299] = 36;
    exp_33_ram[1300] = 36;
    exp_33_ram[1301] = 36;
    exp_33_ram[1302] = 36;
    exp_33_ram[1303] = 36;
    exp_33_ram[1304] = 36;
    exp_33_ram[1305] = 36;
    exp_33_ram[1306] = 36;
    exp_33_ram[1307] = 36;
    exp_33_ram[1308] = 36;
    exp_33_ram[1309] = 36;
    exp_33_ram[1310] = 36;
    exp_33_ram[1311] = 36;
    exp_33_ram[1312] = 36;
    exp_33_ram[1313] = 36;
    exp_33_ram[1314] = 36;
    exp_33_ram[1315] = 36;
    exp_33_ram[1316] = 36;
    exp_33_ram[1317] = 36;
    exp_33_ram[1318] = 36;
    exp_33_ram[1319] = 36;
    exp_33_ram[1320] = 36;
    exp_33_ram[1321] = 36;
    exp_33_ram[1322] = 36;
    exp_33_ram[1323] = 36;
    exp_33_ram[1324] = 36;
    exp_33_ram[1325] = 36;
    exp_33_ram[1326] = 36;
    exp_33_ram[1327] = 36;
    exp_33_ram[1328] = 36;
    exp_33_ram[1329] = 36;
    exp_33_ram[1330] = 36;
    exp_33_ram[1331] = 36;
    exp_33_ram[1332] = 36;
    exp_33_ram[1333] = 36;
    exp_33_ram[1334] = 36;
    exp_33_ram[1335] = 36;
    exp_33_ram[1336] = 36;
    exp_33_ram[1337] = 36;
    exp_33_ram[1338] = 36;
    exp_33_ram[1339] = 36;
    exp_33_ram[1340] = 36;
    exp_33_ram[1341] = 36;
    exp_33_ram[1342] = 36;
    exp_33_ram[1343] = 36;
    exp_33_ram[1344] = 8;
    exp_33_ram[1345] = 36;
    exp_33_ram[1346] = 36;
    exp_33_ram[1347] = 36;
    exp_33_ram[1348] = 36;
    exp_33_ram[1349] = 36;
    exp_33_ram[1350] = 36;
    exp_33_ram[1351] = 36;
    exp_33_ram[1352] = 36;
    exp_33_ram[1353] = 36;
    exp_33_ram[1354] = 8;
    exp_33_ram[1355] = 84;
    exp_33_ram[1356] = 8;
    exp_33_ram[1357] = 36;
    exp_33_ram[1358] = 36;
    exp_33_ram[1359] = 36;
    exp_33_ram[1360] = 36;
    exp_33_ram[1361] = 8;
    exp_33_ram[1362] = 36;
    exp_33_ram[1363] = 36;
    exp_33_ram[1364] = 36;
    exp_33_ram[1365] = 36;
    exp_33_ram[1366] = 36;
    exp_33_ram[1367] = 8;
    exp_33_ram[1368] = 132;
    exp_33_ram[1369] = 36;
    exp_33_ram[1370] = 36;
    exp_33_ram[1371] = 48;
    exp_33_ram[1372] = 36;
    exp_33_ram[1373] = 8;
    exp_33_ram[1374] = 36;
    exp_33_ram[1375] = 36;
    exp_33_ram[1376] = 8;
    exp_33_ram[1377] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_179;

  reg [31:0] exp_179_reg;
  always@(*) begin
    case (exp_177)
      0:exp_179_reg <= exp_157;
      1:exp_179_reg <= exp_167;
      default:exp_179_reg <= exp_178;
    endcase
  end
  assign exp_179 = exp_179_reg;
  assign exp_177 = exp_139[2:2];
  assign exp_139 = exp_1;
  assign exp_178 = 0;

      reg [31:0] exp_157_reg = 0;
      always@(posedge clk) begin
        if (exp_156) begin
          exp_157_reg <= exp_164;
        end
      end
      assign exp_157 = exp_157_reg;
    
  reg [31:0] exp_164_reg;
  always@(*) begin
    case (exp_159)
      0:exp_164_reg <= exp_161;
      1:exp_164_reg <= exp_162;
      default:exp_164_reg <= exp_163;
    endcase
  end
  assign exp_164 = exp_164_reg;
  assign exp_159 = exp_157 == exp_158;
  assign exp_158 = 4294967295;
  assign exp_163 = 0;
  assign exp_161 = exp_157 + exp_160;
  assign exp_160 = 1;
  assign exp_162 = 0;
  assign exp_156 = 1;

      reg [31:0] exp_167_reg = 0;
      always@(posedge clk) begin
        if (exp_166) begin
          exp_167_reg <= exp_174;
        end
      end
      assign exp_167 = exp_167_reg;
    
  reg [31:0] exp_174_reg;
  always@(*) begin
    case (exp_169)
      0:exp_174_reg <= exp_171;
      1:exp_174_reg <= exp_172;
      default:exp_174_reg <= exp_173;
    endcase
  end
  assign exp_174 = exp_174_reg;
  assign exp_169 = exp_167 == exp_168;
  assign exp_168 = 4294967295;
  assign exp_173 = 0;
  assign exp_171 = exp_167 + exp_170;
  assign exp_170 = 1;
  assign exp_172 = 0;
  assign exp_166 = exp_159 & exp_165;
  assign exp_165 = 1;
  assign exp_182 = exp_201;
  assign exp_201 = 0;
  assign exp_204 = exp_219;
  assign exp_219 = stdin_in;
  assign exp_439 = exp_226[15:8];
  assign exp_440 = exp_226[23:16];
  assign exp_441 = exp_226[31:24];
  assign exp_453 = $signed(exp_452);
  assign exp_452 = exp_451 + exp_447;
  assign exp_451 = 0;

  reg [15:0] exp_447_reg;
  always@(*) begin
    case (exp_437)
      0:exp_447_reg <= exp_444;
      1:exp_447_reg <= exp_445;
      default:exp_447_reg <= exp_446;
    endcase
  end
  assign exp_447 = exp_447_reg;
  assign exp_446 = 0;
  assign exp_444 = exp_226[15:0];
  assign exp_445 = exp_226[31:16];
  assign exp_454 = 0;
  assign exp_455 = exp_443;
  assign exp_456 = exp_447;
  assign exp_457 = 0;
  assign exp_458 = 0;

  reg [31:0] exp_817_reg;
  always@(*) begin
    case (exp_607)
      0:exp_817_reg <= exp_813;
      1:exp_817_reg <= exp_815;
      default:exp_817_reg <= exp_816;
    endcase
  end
  assign exp_817 = exp_817_reg;
  assign exp_816 = 0;

  reg [31:0] exp_813_reg;
  always@(*) begin
    case (exp_584)
      0:exp_813_reg <= exp_808;
      1:exp_813_reg <= exp_809;
      default:exp_813_reg <= exp_812;
    endcase
  end
  assign exp_813 = exp_813_reg;
  assign exp_584 = exp_583 & exp_581;
  assign exp_583 = exp_576 == exp_582;
  assign exp_582 = 0;
  assign exp_812 = 0;
  assign exp_808 = exp_807[63:32];

  reg [63:0] exp_807_reg;
  always@(*) begin
    case (exp_804)
      0:exp_807_reg <= exp_803;
      1:exp_807_reg <= exp_805;
      default:exp_807_reg <= exp_806;
    endcase
  end
  assign exp_807 = exp_807_reg;

      reg [0:0] exp_804_reg = 0;
      always@(posedge clk) begin
        if (exp_789) begin
          exp_804_reg <= exp_787;
        end
      end
      assign exp_804 = exp_804_reg;
    
      reg [0:0] exp_787_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_787_reg <= exp_764;
        end
      end
      assign exp_787 = exp_787_reg;
    
      reg [0:0] exp_764_reg = 0;
      always@(posedge clk) begin
        if (exp_746) begin
          exp_764_reg <= exp_761;
        end
      end
      assign exp_764 = exp_764_reg;
      assign exp_761 = exp_759 ^ exp_760;
  assign exp_759 = exp_741 & exp_724;
  assign exp_741 = exp_740 + exp_739;
  assign exp_740 = 0;
  assign exp_739 = exp_737[31:31];

      reg [31:0] exp_737_reg = 0;
      always@(posedge clk) begin
        if (exp_736) begin
          exp_737_reg <= exp_354;
        end
      end
      assign exp_737 = exp_737_reg;
      assign exp_736 = exp_726 == exp_735;
  assign exp_735 = 0;
  assign exp_724 = exp_723 | exp_590;
  assign exp_723 = exp_584 | exp_587;
  assign exp_587 = exp_586 & exp_581;
  assign exp_586 = exp_576 == exp_585;
  assign exp_585 = 1;
  assign exp_590 = exp_589 & exp_581;
  assign exp_589 = exp_576 == exp_588;
  assign exp_588 = 2;
  assign exp_760 = exp_744 & exp_725;
  assign exp_744 = exp_743 + exp_742;
  assign exp_743 = 0;
  assign exp_742 = exp_738[31:31];

      reg [31:0] exp_738_reg = 0;
      always@(posedge clk) begin
        if (exp_736) begin
          exp_738_reg <= exp_355;
        end
      end
      assign exp_738 = exp_738_reg;
      assign exp_725 = exp_584 | exp_587;
  assign exp_746 = exp_726 == exp_745;
  assign exp_745 = 1;
  assign exp_766 = exp_726 == exp_765;
  assign exp_765 = 2;
  assign exp_789 = exp_726 == exp_788;
  assign exp_788 = 3;
  assign exp_806 = 0;

      reg [63:0] exp_803_reg = 0;
      always@(posedge clk) begin
        if (exp_789) begin
          exp_803_reg <= exp_802;
        end
      end
      assign exp_803 = exp_803_reg;
      assign exp_802 = exp_798 + exp_801;
  assign exp_798 = exp_794 + exp_797;
  assign exp_794 = exp_790 + exp_793;
  assign exp_790 = exp_783;

      reg [31:0] exp_783_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_783_reg <= exp_770;
        end
      end
      assign exp_783 = exp_783_reg;
      assign exp_770 = exp_768 * exp_769;
  assign exp_768 = exp_767;
  assign exp_767 = exp_762[15:0];

      reg [31:0] exp_762_reg = 0;
      always@(posedge clk) begin
        if (exp_746) begin
          exp_762_reg <= exp_752;
        end
      end
      assign exp_762 = exp_762_reg;
      assign exp_752 = exp_751 + exp_750;
  assign exp_751 = 0;

  reg [31:0] exp_750_reg;
  always@(*) begin
    case (exp_747)
      0:exp_750_reg <= exp_737;
      1:exp_750_reg <= exp_748;
      default:exp_750_reg <= exp_749;
    endcase
  end
  assign exp_750 = exp_750_reg;
  assign exp_747 = exp_741 & exp_724;
  assign exp_749 = 0;
  assign exp_748 = -exp_737;
  assign exp_769 = exp_763[15:0];

      reg [31:0] exp_763_reg = 0;
      always@(posedge clk) begin
        if (exp_746) begin
          exp_763_reg <= exp_758;
        end
      end
      assign exp_763 = exp_763_reg;
      assign exp_758 = exp_757 + exp_756;
  assign exp_757 = 0;

  reg [31:0] exp_756_reg;
  always@(*) begin
    case (exp_753)
      0:exp_756_reg <= exp_738;
      1:exp_756_reg <= exp_754;
      default:exp_756_reg <= exp_755;
    endcase
  end
  assign exp_756 = exp_756_reg;
  assign exp_753 = exp_744 & exp_725;
  assign exp_755 = 0;
  assign exp_754 = -exp_738;
  assign exp_793 = exp_791 << exp_792;
  assign exp_791 = exp_784;

      reg [31:0] exp_784_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_784_reg <= exp_774;
        end
      end
      assign exp_784 = exp_784_reg;
      assign exp_774 = exp_772 * exp_773;
  assign exp_772 = exp_771;
  assign exp_771 = exp_762[15:0];
  assign exp_773 = exp_763[31:16];
  assign exp_792 = 16;
  assign exp_797 = exp_795 << exp_796;
  assign exp_795 = exp_785;

      reg [31:0] exp_785_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_785_reg <= exp_778;
        end
      end
      assign exp_785 = exp_785_reg;
      assign exp_778 = exp_776 * exp_777;
  assign exp_776 = exp_775;
  assign exp_775 = exp_762[31:16];
  assign exp_777 = exp_763[15:0];
  assign exp_796 = 16;
  assign exp_801 = exp_799 << exp_800;
  assign exp_799 = exp_786;

      reg [31:0] exp_786_reg = 0;
      always@(posedge clk) begin
        if (exp_766) begin
          exp_786_reg <= exp_782;
        end
      end
      assign exp_786 = exp_786_reg;
      assign exp_782 = exp_780 * exp_781;
  assign exp_780 = exp_779;
  assign exp_779 = exp_762[31:16];
  assign exp_781 = exp_763[31:16];
  assign exp_800 = 32;
  assign exp_805 = -exp_803;
  assign exp_809 = exp_807[31:0];

  reg [31:0] exp_815_reg;
  always@(*) begin
    case (exp_608)
      0:exp_815_reg <= exp_718;
      1:exp_815_reg <= exp_719;
      default:exp_815_reg <= exp_814;
    endcase
  end
  assign exp_815 = exp_815_reg;
  assign exp_608 = exp_576[1:1];
  assign exp_814 = 0;

      reg [31:0] exp_718_reg = 0;
      always@(posedge clk) begin
        if (exp_627) begin
          exp_718_reg <= exp_712;
        end
      end
      assign exp_718 = exp_718_reg;
    
  reg [31:0] exp_712_reg;
  always@(*) begin
    case (exp_708)
      0:exp_712_reg <= exp_699;
      1:exp_712_reg <= exp_710;
      default:exp_712_reg <= exp_711;
    endcase
  end
  assign exp_712 = exp_712_reg;
  assign exp_708 = exp_707 & exp_610;
  assign exp_707 = exp_656 == exp_706;

      reg [31:0] exp_656_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_656_reg <= exp_653;
        end
      end
      assign exp_656 = exp_656_reg;
      assign exp_653 = exp_652 + exp_651;
  assign exp_652 = 0;

  reg [31:0] exp_651_reg;
  always@(*) begin
    case (exp_648)
      0:exp_651_reg <= exp_633;
      1:exp_651_reg <= exp_649;
      default:exp_651_reg <= exp_650;
    endcase
  end
  assign exp_651 = exp_651_reg;
  assign exp_648 = exp_639 & exp_610;
  assign exp_639 = exp_638 + exp_637;
  assign exp_638 = 0;
  assign exp_637 = exp_633[31:31];

      reg [31:0] exp_633_reg = 0;
      always@(posedge clk) begin
        if (exp_631) begin
          exp_633_reg <= exp_355;
        end
      end
      assign exp_633 = exp_633_reg;
      assign exp_631 = exp_613 == exp_630;
  assign exp_630 = 0;
  assign exp_610 = ~exp_609;
  assign exp_609 = exp_576[0:0];
  assign exp_650 = 0;
  assign exp_649 = -exp_633;
  assign exp_641 = exp_613 == exp_640;
  assign exp_640 = 1;
  assign exp_706 = 0;
  assign exp_711 = 0;
  assign exp_699 = exp_698 + exp_697;
  assign exp_698 = 0;

  reg [31:0] exp_697_reg;
  always@(*) begin
    case (exp_694)
      0:exp_697_reg <= exp_692;
      1:exp_697_reg <= exp_695;
      default:exp_697_reg <= exp_696;
    endcase
  end
  assign exp_697 = exp_697_reg;
  assign exp_694 = exp_658 & exp_610;

      reg [0:0] exp_658_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_658_reg <= exp_654;
        end
      end
      assign exp_658 = exp_658_reg;
      assign exp_654 = exp_636 ^ exp_639;
  assign exp_636 = exp_635 + exp_634;
  assign exp_635 = 0;
  assign exp_634 = exp_632[31:31];

      reg [31:0] exp_632_reg = 0;
      always@(posedge clk) begin
        if (exp_631) begin
          exp_632_reg <= exp_354;
        end
      end
      assign exp_632 = exp_632_reg;
      assign exp_696 = 0;

      reg [31:0] exp_692_reg = 0;
      always@(posedge clk) begin
        if (exp_625) begin
          exp_692_reg <= exp_662;
        end
      end
      assign exp_692 = exp_692_reg;
    
      reg [31:0] exp_662_reg = 0;
      always@(posedge clk) begin
        if (exp_661) begin
          exp_662_reg <= exp_689;
        end
      end
      assign exp_662 = exp_662_reg;
    
  reg [31:0] exp_689_reg;
  always@(*) begin
    case (exp_623)
      0:exp_689_reg <= exp_681;
      1:exp_689_reg <= exp_687;
      default:exp_689_reg <= exp_688;
    endcase
  end
  assign exp_689 = exp_689_reg;
  assign exp_623 = exp_613 == exp_622;
  assign exp_622 = 2;
  assign exp_688 = 0;

  reg [31:0] exp_681_reg;
  always@(*) begin
    case (exp_671)
      0:exp_681_reg <= exp_675;
      1:exp_681_reg <= exp_679;
      default:exp_681_reg <= exp_680;
    endcase
  end
  assign exp_681 = exp_681_reg;
  assign exp_671 = ~exp_670;
  assign exp_670 = exp_669[32:32];
  assign exp_669 = exp_668 - exp_656;
  assign exp_668 = exp_667;
  assign exp_667 = {exp_665, exp_666};  assign exp_665 = exp_660[31:0];

      reg [31:0] exp_660_reg = 0;
      always@(posedge clk) begin
        if (exp_659) begin
          exp_660_reg <= exp_686;
        end
      end
      assign exp_660 = exp_660_reg;
    
  reg [32:0] exp_686_reg;
  always@(*) begin
    case (exp_623)
      0:exp_686_reg <= exp_673;
      1:exp_686_reg <= exp_684;
      default:exp_686_reg <= exp_685;
    endcase
  end
  assign exp_686 = exp_686_reg;
  assign exp_685 = 0;

  reg [32:0] exp_673_reg;
  always@(*) begin
    case (exp_671)
      0:exp_673_reg <= exp_667;
      1:exp_673_reg <= exp_669;
      default:exp_673_reg <= exp_672;
    endcase
  end
  assign exp_673 = exp_673_reg;
  assign exp_672 = 0;
  assign exp_684 = 0;
  assign exp_659 = 1;
  assign exp_666 = exp_664[31:31];

      reg [31:0] exp_664_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_664_reg <= exp_691;
        end
      end
      assign exp_664 = exp_664_reg;
    
  reg [31:0] exp_691_reg;
  always@(*) begin
    case (exp_623)
      0:exp_691_reg <= exp_683;
      1:exp_691_reg <= exp_655;
      default:exp_691_reg <= exp_690;
    endcase
  end
  assign exp_691 = exp_691_reg;
  assign exp_690 = 0;
  assign exp_683 = exp_664 << exp_682;
  assign exp_682 = 1;

      reg [31:0] exp_655_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_655_reg <= exp_647;
        end
      end
      assign exp_655 = exp_655_reg;
      assign exp_647 = exp_646 + exp_645;
  assign exp_646 = 0;

  reg [31:0] exp_645_reg;
  always@(*) begin
    case (exp_642)
      0:exp_645_reg <= exp_632;
      1:exp_645_reg <= exp_643;
      default:exp_645_reg <= exp_644;
    endcase
  end
  assign exp_645 = exp_645_reg;
  assign exp_642 = exp_636 & exp_610;
  assign exp_644 = 0;
  assign exp_643 = -exp_632;
  assign exp_663 = 1;
  assign exp_680 = 0;
  assign exp_675 = exp_662 << exp_674;
  assign exp_674 = 1;
  assign exp_679 = exp_677 | exp_678;
  assign exp_677 = exp_662 << exp_676;
  assign exp_676 = 1;
  assign exp_678 = 1;
  assign exp_687 = 0;
  assign exp_661 = 1;
  assign exp_625 = exp_613 == exp_624;
  assign exp_624 = 35;
  assign exp_695 = -exp_692;
  assign exp_710 = $signed(exp_709);
  assign exp_709 = -1;
  assign exp_627 = exp_613 == exp_626;
  assign exp_626 = 36;

      reg [31:0] exp_719_reg = 0;
      always@(posedge clk) begin
        if (exp_627) begin
          exp_719_reg <= exp_717;
        end
      end
      assign exp_719 = exp_719_reg;
    
  reg [31:0] exp_717_reg;
  always@(*) begin
    case (exp_715)
      0:exp_717_reg <= exp_705;
      1:exp_717_reg <= exp_632;
      default:exp_717_reg <= exp_716;
    endcase
  end
  assign exp_717 = exp_717_reg;
  assign exp_715 = exp_714 & exp_610;
  assign exp_714 = exp_656 == exp_713;
  assign exp_713 = 0;
  assign exp_716 = 0;
  assign exp_705 = exp_704 + exp_703;
  assign exp_704 = 0;

  reg [31:0] exp_703_reg;
  always@(*) begin
    case (exp_700)
      0:exp_703_reg <= exp_693;
      1:exp_703_reg <= exp_701;
      default:exp_703_reg <= exp_702;
    endcase
  end
  assign exp_703 = exp_703_reg;
  assign exp_700 = exp_657 & exp_610;

      reg [0:0] exp_657_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_657_reg <= exp_636;
        end
      end
      assign exp_657 = exp_657_reg;
      assign exp_702 = 0;

      reg [31:0] exp_693_reg = 0;
      always@(posedge clk) begin
        if (exp_625) begin
          exp_693_reg <= exp_660;
        end
      end
      assign exp_693 = exp_693_reg;
      assign exp_701 = -exp_693;
  assign exp_288 = $signed(exp_287);
  assign exp_287 = 0;
  assign exp_517 = exp_352 != exp_353;
  assign exp_530 = 0;
  assign exp_531 = 0;
  assign exp_518 = $signed(exp_352) < $signed(exp_353);
  assign exp_519 = $signed(exp_352) >= $signed(exp_353);
  assign exp_524 = exp_521 < exp_523;
  assign exp_521 = exp_520 + exp_352;
  assign exp_520 = 0;
  assign exp_523 = exp_522 + exp_353;
  assign exp_522 = 0;
  assign exp_529 = exp_526 >= exp_528;
  assign exp_526 = exp_525 + exp_352;
  assign exp_525 = 0;
  assign exp_528 = exp_527 + exp_353;
  assign exp_527 = 0;
  assign exp_844 = 0;
  assign exp_843 = exp_242 + exp_842;
  assign exp_842 = 4;

  reg [32:0] exp_574_reg;
  always@(*) begin
    case (exp_375)
      0:exp_574_reg <= exp_564;
      1:exp_574_reg <= exp_572;
      default:exp_574_reg <= exp_573;
    endcase
  end
  assign exp_574 = exp_574_reg;
  assign exp_573 = 0;
  assign exp_564 = exp_563 + exp_361;

  reg [31:0] exp_563_reg;
  always@(*) begin
    case (exp_373)
      0:exp_563_reg <= exp_549;
      1:exp_563_reg <= exp_561;
      default:exp_563_reg <= exp_562;
    endcase
  end
  assign exp_563 = exp_563_reg;
  assign exp_562 = 0;
  assign exp_549 = $signed(exp_548);
  assign exp_548 = exp_547 + exp_546;
  assign exp_547 = 0;
  assign exp_546 = {exp_545, exp_542};  assign exp_545 = {exp_544, exp_541};  assign exp_544 = {exp_543, exp_540};  assign exp_543 = {exp_538, exp_539};  assign exp_538 = exp_360[31:31];
  assign exp_539 = exp_360[7:7];
  assign exp_540 = exp_360[30:25];
  assign exp_541 = exp_360[11:8];
  assign exp_542 = 0;
  assign exp_561 = $signed(exp_560);
  assign exp_560 = exp_559 + exp_558;
  assign exp_559 = 0;
  assign exp_558 = {exp_557, exp_554};  assign exp_557 = {exp_556, exp_553};  assign exp_556 = {exp_555, exp_552};  assign exp_555 = {exp_550, exp_551};  assign exp_550 = exp_360[31:31];
  assign exp_551 = exp_360[19:12];
  assign exp_552 = exp_360[20:20];
  assign exp_553 = exp_360[30:21];
  assign exp_554 = 0;

      reg [31:0] exp_361_reg = 0;
      always@(posedge clk) begin
        if (exp_351) begin
          exp_361_reg <= exp_244;
        end
      end
      assign exp_361 = exp_361_reg;
      assign exp_572 = exp_571 & exp_570;
  assign exp_571 = $signed(exp_569);
  assign exp_569 = exp_352 + exp_568;
  assign exp_568 = $signed(exp_567);
  assign exp_567 = exp_566 + exp_565;
  assign exp_566 = 0;
  assign exp_565 = exp_360[31:20];
  assign exp_570 = 4294967294;
  assign exp_241 = exp_234 & exp_232;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_243;
  assign exp_376 = 3;
  assign exp_222 = ~exp_207;
  assign exp_207 = exp_6;
  assign exp_200 = exp_184 & exp_185;
  assign exp_184 = exp_192;
  assign exp_192 = exp_5 & exp_191;
  assign exp_185 = exp_6;
  assign exp_181 = exp_2;
  assign stdin_ready_out = exp_223;
  assign stdout_valid_out = exp_200;
  assign stdout_out = exp_181;

endmodule