
module soc(clk, stdin_rx, stdout_tx, leds_out);
  input [0:0] stdin_rx;
  input [0:0] clk;
  output [0:0] stdout_tx;
  output [31:0] leds_out;
  wire [0:0] exp_375;
  wire [0:0] exp_372;
  wire [0:0] exp_296;
  wire [0:0] exp_299;
  wire [0:0] exp_294;
  wire [0:0] exp_357;
  wire [0:0] exp_342;
  wire [0:0] exp_356;
  wire [0:0] exp_353;
  wire [0:0] exp_352;
  wire [0:0] exp_316;
  wire [0:0] exp_340;
  wire [0:0] exp_336;
  wire [0:0] exp_301;
  wire [0:0] exp_314;
  wire [0:0] exp_311;
  wire [0:0] exp_293;
  wire [0:0] exp_279;
  wire [0:0] exp_287;
  wire [0:0] exp_11;
  wire [0:0] exp_402;
  wire [0:0] exp_749;
  wire [0:0] exp_686;
  wire [0:0] exp_551;
  wire [6:0] exp_536;
  wire [31:0] exp_534;
  wire [31:0] exp_104;
  wire [31:0] exp_103;
  wire [23:0] exp_102;
  wire [15:0] exp_101;
  wire [7:0] exp_90;
  wire [0:0] exp_89;
  wire [0:0] exp_94;
  wire [12:0] exp_85;
  wire [29:0] exp_93;
  wire [31:0] exp_16;
  wire [31:0] exp_416;
  wire [32:0] exp_1019;
  wire [0:0] exp_1015;
  wire [0:0] exp_711;
  wire [0:0] exp_689;
  wire [0:0] exp_547;
  wire [6:0] exp_546;
  wire [0:0] exp_549;
  wire [6:0] exp_548;
  wire [0:0] exp_710;
  wire [0:0] exp_555;
  wire [6:0] exp_554;
  wire [0:0] exp_709;
  wire [0:0] exp_708;
  wire [0:0] exp_707;
  wire [2:0] exp_537;
  wire [0:0] exp_706;
  wire [0:0] exp_690;
  wire [31:0] exp_526;
  wire [31:0] exp_464;
  wire [0:0] exp_460;
  wire [4:0] exp_440;
  wire [0:0] exp_459;
  wire [0:0] exp_463;
  wire [31:0] exp_456;
  wire [0:0] exp_437;
  wire [0:0] exp_1010;
  wire [0:0] exp_1009;
  wire [0:0] exp_1008;
  wire [0:0] exp_1007;
  wire [4:0] exp_419;
  wire [4:0] exp_1002;
  wire [0:0] exp_1001;
  wire [0:0] exp_593;
  wire [0:0] exp_592;
  wire [0:0] exp_591;
  wire [0:0] exp_590;
  wire [0:0] exp_589;
  wire [0:0] exp_588;
  wire [0:0] exp_539;
  wire [4:0] exp_538;
  wire [0:0] exp_541;
  wire [5:0] exp_540;
  wire [0:0] exp_543;
  wire [5:0] exp_542;
  wire [0:0] exp_545;
  wire [4:0] exp_544;
  wire [0:0] exp_996;
  wire [0:0] exp_995;
  wire [0:0] exp_781;
  wire [0:0] exp_755;
  wire [0:0] exp_753;
  wire [6:0] exp_751;
  wire [5:0] exp_752;
  wire [0:0] exp_754;
  wire [0:0] exp_780;
  wire [2:0] exp_750;
  wire [0:0] exp_994;
  wire [0:0] exp_992;
  wire [0:0] exp_985;
  wire [2:0] exp_900;
  wire [2:0] exp_907;
  wire [0:0] exp_902;
  wire [2:0] exp_901;
  wire [0:0] exp_906;
  wire [2:0] exp_904;
  wire [0:0] exp_903;
  wire [0:0] exp_905;
  wire [0:0] exp_896;
  wire [0:0] exp_895;
  wire [0:0] exp_894;
  wire [2:0] exp_984;
  wire [0:0] exp_993;
  wire [0:0] exp_803;
  wire [5:0] exp_787;
  wire [5:0] exp_794;
  wire [0:0] exp_789;
  wire [5:0] exp_788;
  wire [0:0] exp_793;
  wire [5:0] exp_791;
  wire [0:0] exp_790;
  wire [0:0] exp_792;
  wire [5:0] exp_802;
  wire [0:0] exp_414;
  wire [0:0] exp_413;
  wire [0:0] exp_411;
  wire [0:0] exp_410;
  wire [0:0] exp_408;
  wire [0:0] exp_409;
  wire [0:0] exp_407;
  wire [0:0] exp_1020;
  wire [0:0] exp_406;
  wire [0:0] exp_405;
  wire [0:0] exp_1024;
  wire [0:0] exp_1023;
  wire [0:0] exp_1022;
  wire [0:0] exp_1021;
  wire [0:0] exp_401;
  wire [0:0] exp_393;
  wire [0:0] exp_291;
  wire [0:0] exp_204;
  wire [0:0] exp_163;
  wire [0:0] exp_34;
  wire [0:0] exp_15;
  wire [0:0] exp_33;
  wire [0:0] exp_29;
  wire [0:0] exp_26;
  wire [31:0] exp_9;
  wire [31:0] exp_398;
  wire [31:0] exp_605;
  wire [31:0] exp_604;
  wire [31:0] exp_603;
  wire [31:0] exp_602;
  wire [11:0] exp_601;
  wire [11:0] exp_600;
  wire [11:0] exp_599;
  wire [0:0] exp_553;
  wire [5:0] exp_552;
  wire [0:0] exp_598;
  wire [11:0] exp_594;
  wire [11:0] exp_597;
  wire [6:0] exp_595;
  wire [4:0] exp_596;
  wire [0:0] exp_25;
  wire [0:0] exp_28;
  wire [14:0] exp_27;
  wire [0:0] exp_21;
  wire [0:0] exp_146;
  wire [0:0] exp_23;
  wire [0:0] exp_12;
  wire [0:0] exp_403;
  wire [0:0] exp_688;
  wire [0:0] exp_687;
  wire [0:0] exp_145;
  wire [0:0] exp_140;
  wire [0:0] exp_144;
  wire [0:0] exp_142;
  wire [0:0] exp_22;
  wire [0:0] exp_30;
  wire [0:0] exp_141;
  wire [0:0] exp_143;
  wire [0:0] exp_139;
  wire [0:0] exp_125;
  wire [0:0] exp_162;
  wire [0:0] exp_158;
  wire [0:0] exp_155;
  wire [31:0] exp_154;
  wire [0:0] exp_157;
  wire [31:0] exp_156;
  wire [0:0] exp_150;
  wire [0:0] exp_184;
  wire [0:0] exp_203;
  wire [0:0] exp_199;
  wire [0:0] exp_196;
  wire [31:0] exp_195;
  wire [0:0] exp_198;
  wire [31:0] exp_197;
  wire [0:0] exp_191;
  wire [0:0] exp_261;
  wire [0:0] exp_266;
  wire [0:0] exp_263;
  wire [0:0] exp_262;
  wire [0:0] exp_235;
  wire [0:0] exp_259;
  wire [0:0] exp_255;
  wire [0:0] exp_219;
  wire [0:0] exp_233;
  wire [0:0] exp_230;
  wire [0:0] exp_215;
  wire [0:0] exp_217;
  wire [0:0] exp_213;
  wire [0:0] exp_267;
  wire [0:0] exp_206;
  wire [0:0] exp_192;
  wire [0:0] exp_200;
  wire [0:0] exp_205;
  wire [0:0] exp_193;
  wire [0:0] exp_216;
  wire [0:0] exp_212;
  wire [0:0] exp_210;
  wire [0:0] exp_208;
  wire [0:0] exp_7;
  wire [0:0] exp_207;
  wire [0:0] exp_209;
  wire [0:0] exp_211;
  wire [0:0] exp_214;
  wire [0:0] exp_229;
  wire [0:0] exp_232;
  wire [0:0] exp_231;
  wire [0:0] exp_228;
  wire [0:0] exp_222;
  wire [9:0] exp_220;
  wire [9:0] exp_227;
  wire [0:0] exp_226;
  wire [9:0] exp_224;
  wire [0:0] exp_223;
  wire [0:0] exp_225;
  wire [9:0] exp_221;
  wire [0:0] exp_218;
  wire [0:0] exp_258;
  wire [0:0] exp_257;
  wire [0:0] exp_256;
  wire [0:0] exp_244;
  wire [0:0] exp_238;
  wire [8:0] exp_236;
  wire [8:0] exp_243;
  wire [0:0] exp_242;
  wire [8:0] exp_240;
  wire [0:0] exp_239;
  wire [0:0] exp_241;
  wire [8:0] exp_237;
  wire [0:0] exp_254;
  wire [0:0] exp_248;
  wire [2:0] exp_246;
  wire [2:0] exp_253;
  wire [0:0] exp_252;
  wire [2:0] exp_250;
  wire [0:0] exp_249;
  wire [0:0] exp_251;
  wire [0:0] exp_245;
  wire [2:0] exp_247;
  wire [0:0] exp_234;
  wire [0:0] exp_265;
  wire [0:0] exp_264;
  wire [0:0] exp_260;
  wire [0:0] exp_290;
  wire [0:0] exp_286;
  wire [0:0] exp_283;
  wire [31:0] exp_282;
  wire [0:0] exp_285;
  wire [31:0] exp_284;
  wire [0:0] exp_278;
  wire [0:0] exp_392;
  wire [0:0] exp_388;
  wire [0:0] exp_385;
  wire [31:0] exp_384;
  wire [0:0] exp_387;
  wire [31:0] exp_386;
  wire [0:0] exp_380;
  wire [0:0] exp_397;
  wire [0:0] exp_998;
  wire [0:0] exp_997;
  wire [0:0] exp_412;
  wire [0:0] exp_455;
  wire [31:0] exp_427;
  wire [0:0] exp_426;
  wire [1:0] exp_435;
  wire [4:0] exp_422;
  wire [0:0] exp_425;
  wire [0:0] exp_1004;
  wire [0:0] exp_1003;
  wire [4:0] exp_421;
  wire [31:0] exp_423;
  wire [31:0] exp_1000;
  wire [0:0] exp_999;
  wire [31:0] exp_636;
  wire [0:0] exp_635;
  wire [31:0] exp_587;
  wire [2:0] exp_530;
  wire [2:0] exp_521;
  wire [0:0] exp_518;
  wire [0:0] exp_452;
  wire [6:0] exp_442;
  wire [6:0] exp_451;
  wire [0:0] exp_454;
  wire [6:0] exp_453;
  wire [0:0] exp_520;
  wire [2:0] exp_508;
  wire [0:0] exp_450;
  wire [4:0] exp_449;
  wire [0:0] exp_507;
  wire [2:0] exp_495;
  wire [0:0] exp_448;
  wire [5:0] exp_447;
  wire [0:0] exp_494;
  wire [2:0] exp_444;
  wire [0:0] exp_493;
  wire [0:0] exp_506;
  wire [0:0] exp_519;
  wire [0:0] exp_525;
  wire [0:0] exp_586;
  wire [31:0] exp_566;
  wire [0:0] exp_532;
  wire [0:0] exp_524;
  wire [0:0] exp_510;
  wire [0:0] exp_497;
  wire [0:0] exp_483;
  wire [0:0] exp_481;
  wire [0:0] exp_482;
  wire [0:0] exp_446;
  wire [4:0] exp_445;
  wire [0:0] exp_496;
  wire [0:0] exp_509;
  wire [0:0] exp_523;
  wire [0:0] exp_522;
  wire [0:0] exp_565;
  wire [31:0] exp_563;
  wire [31:0] exp_528;
  wire [31:0] exp_514;
  wire [0:0] exp_511;
  wire [0:0] exp_513;
  wire [31:0] exp_503;
  wire [0:0] exp_502;
  wire [31:0] exp_489;
  wire [0:0] exp_488;
  wire [31:0] exp_487;
  wire [31:0] exp_485;
  wire [19:0] exp_484;
  wire [3:0] exp_486;
  wire [31:0] exp_501;
  wire [31:0] exp_499;
  wire [19:0] exp_498;
  wire [3:0] exp_500;
  wire [31:0] exp_512;
  wire [31:0] exp_529;
  wire [31:0] exp_517;
  wire [0:0] exp_515;
  wire [0:0] exp_516;
  wire [31:0] exp_505;
  wire [0:0] exp_504;
  wire [31:0] exp_492;
  wire [0:0] exp_491;
  wire [31:0] exp_476;
  wire [0:0] exp_475;
  wire [31:0] exp_470;
  wire [0:0] exp_466;
  wire [4:0] exp_441;
  wire [0:0] exp_465;
  wire [0:0] exp_469;
  wire [31:0] exp_458;
  wire [0:0] exp_438;
  wire [0:0] exp_1014;
  wire [0:0] exp_1013;
  wire [0:0] exp_1012;
  wire [0:0] exp_1011;
  wire [4:0] exp_420;
  wire [0:0] exp_457;
  wire [31:0] exp_434;
  wire [0:0] exp_433;
  wire [1:0] exp_436;
  wire [4:0] exp_429;
  wire [0:0] exp_432;
  wire [0:0] exp_1006;
  wire [0:0] exp_1005;
  wire [4:0] exp_428;
  wire [31:0] exp_430;
  wire [31:0] exp_439;
  wire [31:0] exp_468;
  wire [0:0] exp_467;
  wire [31:0] exp_474;
  wire [31:0] exp_471;
  wire [31:0] exp_473;
  wire [11:0] exp_472;
  wire [31:0] exp_490;
  wire [31:0] exp_418;
  wire [0:0] exp_417;
  wire [31:0] exp_564;
  wire [31:0] exp_568;
  wire [31:0] exp_567;
  wire [5:0] exp_562;
  wire [5:0] exp_561;
  wire [5:0] exp_560;
  wire [4:0] exp_531;
  wire [4:0] exp_480;
  wire [0:0] exp_479;
  wire [4:0] exp_478;
  wire [4:0] exp_443;
  wire [31:0] exp_584;
  wire [1:0] exp_570;
  wire [0:0] exp_569;
  wire [31:0] exp_585;
  wire [1:0] exp_576;
  wire [0:0] exp_575;
  wire [31:0] exp_572;
  wire [31:0] exp_571;
  wire [31:0] exp_574;
  wire [31:0] exp_573;
  wire [31:0] exp_577;
  wire [31:0] exp_581;
  wire [32:0] exp_580;
  wire [32:0] exp_578;
  wire [0:0] exp_559;
  wire [0:0] exp_533;
  wire [0:0] exp_477;
  wire [0:0] exp_558;
  wire [0:0] exp_557;
  wire [0:0] exp_556;
  wire [32:0] exp_579;
  wire [31:0] exp_582;
  wire [31:0] exp_583;
  wire [31:0] exp_634;
  wire [0:0] exp_633;
  wire [31:0] exp_624;
  wire [7:0] exp_623;
  wire [7:0] exp_622;
  wire [7:0] exp_617;
  wire [1:0] exp_608;
  wire [1:0] exp_607;
  wire [1:0] exp_606;
  wire [0:0] exp_616;
  wire [7:0] exp_612;
  wire [31:0] exp_400;
  wire [31:0] exp_391;
  wire [0:0] exp_390;
  wire [31:0] exp_289;
  wire [0:0] exp_288;
  wire [31:0] exp_202;
  wire [0:0] exp_201;
  wire [31:0] exp_161;
  wire [0:0] exp_160;
  wire [31:0] exp_32;
  wire [0:0] exp_31;
  wire [31:0] exp_14;
  wire [31:0] exp_20;
  wire [31:0] exp_127;
  wire [31:0] exp_138;
  wire [23:0] exp_137;
  wire [15:0] exp_136;
  wire [7:0] exp_62;
  wire [0:0] exp_61;
  wire [0:0] exp_129;
  wire [12:0] exp_57;
  wire [29:0] exp_128;
  wire [31:0] exp_18;
  wire [0:0] exp_60;
  wire [0:0] exp_124;
  wire [0:0] exp_122;
  wire [0:0] exp_123;
  wire [3:0] exp_24;
  wire [3:0] exp_13;
  wire [3:0] exp_404;
  wire [3:0] exp_685;
  wire [0:0] exp_684;
  wire [3:0] exp_672;
  wire [3:0] exp_668;
  wire [1:0] exp_671;
  wire [1:0] exp_670;
  wire [1:0] exp_669;
  wire [3:0] exp_677;
  wire [3:0] exp_673;
  wire [0:0] exp_676;
  wire [0:0] exp_675;
  wire [0:0] exp_674;
  wire [3:0] exp_678;
  wire [3:0] exp_679;
  wire [3:0] exp_680;
  wire [3:0] exp_681;
  wire [3:0] exp_682;
  wire [3:0] exp_683;
  wire [12:0] exp_56;
  wire [29:0] exp_120;
  wire [7:0] exp_58;
  wire [7:0] exp_121;
  wire [31:0] exp_19;
  wire [31:0] exp_10;
  wire [31:0] exp_399;
  wire [31:0] exp_667;
  wire [0:0] exp_666;
  wire [31:0] exp_654;
  wire [0:0] exp_653;
  wire [31:0] exp_640;
  wire [7:0] exp_639;
  wire [7:0] exp_638;
  wire [7:0] exp_637;
  wire [31:0] exp_527;
  wire [31:0] exp_648;
  wire [3:0] exp_647;
  wire [31:0] exp_650;
  wire [4:0] exp_649;
  wire [31:0] exp_652;
  wire [4:0] exp_651;
  wire [31:0] exp_658;
  wire [0:0] exp_611;
  wire [0:0] exp_610;
  wire [0:0] exp_609;
  wire [0:0] exp_657;
  wire [31:0] exp_644;
  wire [15:0] exp_643;
  wire [15:0] exp_642;
  wire [15:0] exp_641;
  wire [31:0] exp_656;
  wire [4:0] exp_655;
  wire [31:0] exp_660;
  wire [31:0] exp_659;
  wire [31:0] exp_646;
  wire [31:0] exp_645;
  wire [31:0] exp_661;
  wire [31:0] exp_662;
  wire [31:0] exp_663;
  wire [31:0] exp_664;
  wire [31:0] exp_665;
  wire [7:0] exp_55;
  wire [7:0] exp_83;
  wire [0:0] exp_82;
  wire [0:0] exp_96;
  wire [12:0] exp_78;
  wire [29:0] exp_95;
  wire [0:0] exp_81;
  wire [0:0] exp_92;
  wire [12:0] exp_77;
  wire [31:0] exp_91;
  wire [7:0] exp_79;
  wire [0:0] exp_54;
  wire [0:0] exp_131;
  wire [12:0] exp_50;
  wire [29:0] exp_130;
  wire [0:0] exp_53;
  wire [0:0] exp_119;
  wire [0:0] exp_117;
  wire [0:0] exp_118;
  wire [12:0] exp_49;
  wire [29:0] exp_115;
  wire [7:0] exp_51;
  wire [7:0] exp_116;
  wire [7:0] exp_48;
  wire [7:0] exp_76;
  wire [0:0] exp_75;
  wire [0:0] exp_98;
  wire [12:0] exp_71;
  wire [29:0] exp_97;
  wire [0:0] exp_74;
  wire [12:0] exp_70;
  wire [7:0] exp_72;
  wire [0:0] exp_47;
  wire [0:0] exp_133;
  wire [12:0] exp_43;
  wire [29:0] exp_132;
  wire [0:0] exp_46;
  wire [0:0] exp_114;
  wire [0:0] exp_112;
  wire [0:0] exp_113;
  wire [12:0] exp_42;
  wire [29:0] exp_110;
  wire [7:0] exp_44;
  wire [7:0] exp_111;
  wire [7:0] exp_41;
  wire [7:0] exp_69;
  wire [0:0] exp_68;
  wire [0:0] exp_100;
  wire [12:0] exp_64;
  wire [29:0] exp_99;
  wire [0:0] exp_67;
  wire [12:0] exp_63;
  wire [7:0] exp_65;
  wire [0:0] exp_40;
  wire [0:0] exp_135;
  wire [12:0] exp_36;
  wire [29:0] exp_134;
  wire [0:0] exp_39;
  wire [0:0] exp_109;
  wire [0:0] exp_107;
  wire [0:0] exp_108;
  wire [12:0] exp_35;
  wire [29:0] exp_105;
  wire [7:0] exp_37;
  wire [7:0] exp_106;
  wire [0:0] exp_126;
  wire [31:0] exp_149;
  wire [31:0] exp_187;
  wire [0:0] exp_185;
  wire [31:0] exp_147;
  wire [0:0] exp_186;
  wire [31:0] exp_165;
  wire [31:0] exp_172;
  wire [0:0] exp_167;
  wire [31:0] exp_166;
  wire [0:0] exp_171;
  wire [31:0] exp_169;
  wire [0:0] exp_168;
  wire [0:0] exp_170;
  wire [0:0] exp_164;
  wire [31:0] exp_175;
  wire [31:0] exp_182;
  wire [0:0] exp_177;
  wire [31:0] exp_176;
  wire [0:0] exp_181;
  wire [31:0] exp_179;
  wire [0:0] exp_178;
  wire [0:0] exp_180;
  wire [0:0] exp_174;
  wire [0:0] exp_173;
  wire [31:0] exp_190;
  wire [31:0] exp_274;
  wire [7:0] exp_271;
  wire [7:0] exp_273;
  wire [6:0] exp_272;
  wire [0:0] exp_270;
  wire [0:0] exp_269;
  wire [0:0] exp_268;
  wire [31:0] exp_277;
  wire [31:0] exp_376;
  wire [31:0] exp_379;
  wire [31:0] exp_396;
  wire [7:0] exp_613;
  wire [7:0] exp_614;
  wire [7:0] exp_615;
  wire [31:0] exp_627;
  wire [15:0] exp_626;
  wire [15:0] exp_625;
  wire [15:0] exp_621;
  wire [0:0] exp_620;
  wire [15:0] exp_618;
  wire [15:0] exp_619;
  wire [31:0] exp_628;
  wire [31:0] exp_629;
  wire [31:0] exp_630;
  wire [31:0] exp_631;
  wire [31:0] exp_632;
  wire [31:0] exp_991;
  wire [0:0] exp_990;
  wire [31:0] exp_987;
  wire [0:0] exp_758;
  wire [0:0] exp_757;
  wire [0:0] exp_756;
  wire [0:0] exp_986;
  wire [31:0] exp_982;
  wire [63:0] exp_981;
  wire [0:0] exp_978;
  wire [0:0] exp_961;
  wire [0:0] exp_938;
  wire [0:0] exp_935;
  wire [0:0] exp_933;
  wire [0:0] exp_915;
  wire [0:0] exp_914;
  wire [0:0] exp_913;
  wire [31:0] exp_911;
  wire [0:0] exp_910;
  wire [0:0] exp_909;
  wire [0:0] exp_898;
  wire [0:0] exp_897;
  wire [0:0] exp_761;
  wire [0:0] exp_760;
  wire [0:0] exp_759;
  wire [0:0] exp_764;
  wire [0:0] exp_763;
  wire [1:0] exp_762;
  wire [0:0] exp_934;
  wire [0:0] exp_918;
  wire [0:0] exp_917;
  wire [0:0] exp_916;
  wire [31:0] exp_912;
  wire [0:0] exp_899;
  wire [0:0] exp_920;
  wire [0:0] exp_919;
  wire [0:0] exp_940;
  wire [1:0] exp_939;
  wire [0:0] exp_963;
  wire [1:0] exp_962;
  wire [0:0] exp_980;
  wire [63:0] exp_977;
  wire [63:0] exp_976;
  wire [63:0] exp_972;
  wire [63:0] exp_968;
  wire [63:0] exp_964;
  wire [31:0] exp_957;
  wire [31:0] exp_944;
  wire [31:0] exp_942;
  wire [15:0] exp_941;
  wire [31:0] exp_936;
  wire [31:0] exp_926;
  wire [31:0] exp_925;
  wire [31:0] exp_924;
  wire [0:0] exp_921;
  wire [0:0] exp_923;
  wire [31:0] exp_922;
  wire [15:0] exp_943;
  wire [31:0] exp_937;
  wire [31:0] exp_932;
  wire [31:0] exp_931;
  wire [31:0] exp_930;
  wire [0:0] exp_927;
  wire [0:0] exp_929;
  wire [31:0] exp_928;
  wire [63:0] exp_967;
  wire [63:0] exp_965;
  wire [31:0] exp_958;
  wire [31:0] exp_948;
  wire [31:0] exp_946;
  wire [15:0] exp_945;
  wire [15:0] exp_947;
  wire [4:0] exp_966;
  wire [63:0] exp_971;
  wire [63:0] exp_969;
  wire [31:0] exp_959;
  wire [31:0] exp_952;
  wire [31:0] exp_950;
  wire [15:0] exp_949;
  wire [15:0] exp_951;
  wire [4:0] exp_970;
  wire [63:0] exp_975;
  wire [63:0] exp_973;
  wire [31:0] exp_960;
  wire [31:0] exp_956;
  wire [31:0] exp_954;
  wire [15:0] exp_953;
  wire [15:0] exp_955;
  wire [5:0] exp_974;
  wire [63:0] exp_979;
  wire [31:0] exp_983;
  wire [31:0] exp_989;
  wire [0:0] exp_782;
  wire [0:0] exp_988;
  wire [31:0] exp_892;
  wire [31:0] exp_886;
  wire [0:0] exp_882;
  wire [0:0] exp_881;
  wire [31:0] exp_830;
  wire [31:0] exp_827;
  wire [31:0] exp_826;
  wire [31:0] exp_825;
  wire [0:0] exp_822;
  wire [0:0] exp_813;
  wire [0:0] exp_812;
  wire [0:0] exp_811;
  wire [31:0] exp_807;
  wire [0:0] exp_805;
  wire [0:0] exp_804;
  wire [0:0] exp_784;
  wire [0:0] exp_783;
  wire [0:0] exp_824;
  wire [31:0] exp_823;
  wire [0:0] exp_815;
  wire [0:0] exp_814;
  wire [0:0] exp_880;
  wire [0:0] exp_885;
  wire [31:0] exp_873;
  wire [31:0] exp_872;
  wire [31:0] exp_871;
  wire [0:0] exp_868;
  wire [0:0] exp_832;
  wire [0:0] exp_828;
  wire [0:0] exp_810;
  wire [0:0] exp_809;
  wire [0:0] exp_808;
  wire [31:0] exp_806;
  wire [0:0] exp_870;
  wire [31:0] exp_866;
  wire [31:0] exp_836;
  wire [31:0] exp_863;
  wire [0:0] exp_797;
  wire [1:0] exp_796;
  wire [0:0] exp_862;
  wire [31:0] exp_855;
  wire [0:0] exp_845;
  wire [0:0] exp_844;
  wire [32:0] exp_843;
  wire [32:0] exp_842;
  wire [32:0] exp_841;
  wire [31:0] exp_839;
  wire [31:0] exp_834;
  wire [32:0] exp_860;
  wire [0:0] exp_859;
  wire [32:0] exp_847;
  wire [0:0] exp_846;
  wire [0:0] exp_858;
  wire [0:0] exp_833;
  wire [0:0] exp_840;
  wire [31:0] exp_838;
  wire [31:0] exp_865;
  wire [0:0] exp_864;
  wire [31:0] exp_857;
  wire [0:0] exp_856;
  wire [31:0] exp_829;
  wire [31:0] exp_821;
  wire [31:0] exp_820;
  wire [31:0] exp_819;
  wire [0:0] exp_816;
  wire [0:0] exp_818;
  wire [31:0] exp_817;
  wire [0:0] exp_837;
  wire [0:0] exp_854;
  wire [31:0] exp_849;
  wire [0:0] exp_848;
  wire [31:0] exp_853;
  wire [31:0] exp_851;
  wire [0:0] exp_850;
  wire [0:0] exp_852;
  wire [0:0] exp_861;
  wire [0:0] exp_835;
  wire [0:0] exp_799;
  wire [5:0] exp_798;
  wire [31:0] exp_869;
  wire [31:0] exp_884;
  wire [0:0] exp_883;
  wire [0:0] exp_801;
  wire [5:0] exp_800;
  wire [31:0] exp_893;
  wire [31:0] exp_891;
  wire [0:0] exp_889;
  wire [0:0] exp_888;
  wire [0:0] exp_887;
  wire [0:0] exp_890;
  wire [31:0] exp_879;
  wire [31:0] exp_878;
  wire [31:0] exp_877;
  wire [0:0] exp_874;
  wire [0:0] exp_831;
  wire [0:0] exp_876;
  wire [31:0] exp_867;
  wire [31:0] exp_875;
  wire [31:0] exp_462;
  wire [0:0] exp_461;
  wire [0:0] exp_691;
  wire [0:0] exp_704;
  wire [0:0] exp_705;
  wire [0:0] exp_692;
  wire [0:0] exp_693;
  wire [0:0] exp_698;
  wire [31:0] exp_695;
  wire [31:0] exp_694;
  wire [31:0] exp_697;
  wire [31:0] exp_696;
  wire [0:0] exp_703;
  wire [31:0] exp_700;
  wire [31:0] exp_699;
  wire [31:0] exp_702;
  wire [31:0] exp_701;
  wire [0:0] exp_1018;
  wire [31:0] exp_1017;
  wire [2:0] exp_1016;
  wire [32:0] exp_748;
  wire [0:0] exp_747;
  wire [31:0] exp_738;
  wire [31:0] exp_737;
  wire [0:0] exp_736;
  wire [31:0] exp_723;
  wire [12:0] exp_722;
  wire [12:0] exp_721;
  wire [12:0] exp_720;
  wire [11:0] exp_719;
  wire [7:0] exp_718;
  wire [1:0] exp_717;
  wire [0:0] exp_712;
  wire [0:0] exp_713;
  wire [5:0] exp_714;
  wire [3:0] exp_715;
  wire [0:0] exp_716;
  wire [31:0] exp_735;
  wire [20:0] exp_734;
  wire [20:0] exp_733;
  wire [20:0] exp_732;
  wire [19:0] exp_731;
  wire [9:0] exp_730;
  wire [8:0] exp_729;
  wire [0:0] exp_724;
  wire [7:0] exp_725;
  wire [0:0] exp_726;
  wire [9:0] exp_727;
  wire [0:0] exp_728;
  wire [31:0] exp_535;
  wire [32:0] exp_746;
  wire [32:0] exp_745;
  wire [31:0] exp_743;
  wire [31:0] exp_742;
  wire [11:0] exp_741;
  wire [11:0] exp_740;
  wire [11:0] exp_739;
  wire [32:0] exp_744;
  wire [0:0] exp_415;
  wire [0:0] exp_88;
  wire [12:0] exp_84;
  wire [7:0] exp_86;
  wire [0:0] exp_17;
  wire [1:0] exp_550;
  wire [0:0] exp_280;
  wire [0:0] exp_313;
  wire [0:0] exp_312;
  wire [0:0] exp_310;
  wire [0:0] exp_304;
  wire [8:0] exp_302;
  wire [8:0] exp_309;
  wire [0:0] exp_308;
  wire [8:0] exp_306;
  wire [0:0] exp_305;
  wire [0:0] exp_307;
  wire [8:0] exp_303;
  wire [0:0] exp_300;
  wire [0:0] exp_339;
  wire [0:0] exp_338;
  wire [0:0] exp_337;
  wire [0:0] exp_325;
  wire [0:0] exp_319;
  wire [8:0] exp_317;
  wire [8:0] exp_324;
  wire [0:0] exp_323;
  wire [8:0] exp_321;
  wire [0:0] exp_320;
  wire [0:0] exp_322;
  wire [8:0] exp_318;
  wire [0:0] exp_335;
  wire [0:0] exp_329;
  wire [2:0] exp_327;
  wire [2:0] exp_334;
  wire [0:0] exp_333;
  wire [2:0] exp_331;
  wire [0:0] exp_330;
  wire [0:0] exp_332;
  wire [0:0] exp_326;
  wire [2:0] exp_328;
  wire [0:0] exp_315;
  wire [0:0] exp_355;
  wire [0:0] exp_354;
  wire [0:0] exp_351;
  wire [0:0] exp_345;
  wire [8:0] exp_343;
  wire [8:0] exp_350;
  wire [0:0] exp_349;
  wire [8:0] exp_347;
  wire [0:0] exp_346;
  wire [0:0] exp_348;
  wire [8:0] exp_344;
  wire [0:0] exp_341;
  wire [0:0] exp_298;
  wire [0:0] exp_297;
  wire [0:0] exp_295;
  wire [0:0] exp_374;
  wire [0:0] exp_371;
  wire [0:0] exp_370;
  wire [0:0] exp_368;
  wire [7:0] exp_359;
  wire [7:0] exp_367;
  wire [0:0] exp_365;
  wire [0:0] exp_366;
  wire [7:0] exp_364;
  wire [0:0] exp_360;
  wire [0:0] exp_363;
  wire [7:0] exp_362;
  wire [0:0] exp_361;
  wire [7:0] exp_292;
  wire [31:0] exp_276;
  wire [0:0] exp_358;
  wire [0:0] exp_369;
  wire [0:0] exp_373;
  wire [31:0] exp_395;
  wire [31:0] exp_378;
  wire [0:0] exp_394;
  wire [0:0] exp_381;
  wire [0:0] exp_389;
  wire [0:0] exp_382;


  reg [0:0] exp_375_reg;
  always@(*) begin
    case (exp_372)
      0:exp_375_reg <= exp_371;
      1:exp_375_reg <= exp_373;
      default:exp_375_reg <= exp_374;
    endcase
  end
  assign exp_375 = exp_375_reg;
  assign exp_372 = exp_296 | exp_342;

      reg [0:0] exp_296_reg = 1;
      always@(posedge clk) begin
        if (exp_295) begin
          exp_296_reg <= exp_299;
        end
      end
      assign exp_296 = exp_296_reg;
      assign exp_299 = exp_294 | exp_298;
  assign exp_294 = exp_357;
  assign exp_357 = exp_342 & exp_351;

      reg [0:0] exp_342_reg = 0;
      always@(posedge clk) begin
        if (exp_341) begin
          exp_342_reg <= exp_356;
        end
      end
      assign exp_342 = exp_342_reg;
      assign exp_356 = exp_353 | exp_355;
  assign exp_353 = exp_352 & exp_335;
  assign exp_352 = exp_316 & exp_325;

      reg [0:0] exp_316_reg = 0;
      always@(posedge clk) begin
        if (exp_315) begin
          exp_316_reg <= exp_340;
        end
      end
      assign exp_316 = exp_316_reg;
      assign exp_340 = exp_336 | exp_339;
  assign exp_336 = exp_301 & exp_310;

      reg [0:0] exp_301_reg = 0;
      always@(posedge clk) begin
        if (exp_300) begin
          exp_301_reg <= exp_314;
        end
      end
      assign exp_301 = exp_301_reg;
      assign exp_314 = exp_311 | exp_313;
  assign exp_311 = exp_296 & exp_293;
  assign exp_293 = exp_279 & exp_280;
  assign exp_279 = exp_287;
  assign exp_287 = exp_11 & exp_286;
  assign exp_11 = exp_402;
  assign exp_402 = exp_749;
  assign exp_749 = exp_686 & exp_414;
  assign exp_686 = exp_551 | exp_553;
  assign exp_551 = exp_536 == exp_550;
  assign exp_536 = exp_534[6:0];

      reg [31:0] exp_534_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_534_reg <= exp_104;
        end
      end
      assign exp_534 = exp_534_reg;
    
      reg [31:0] exp_104_reg = 0;
      always@(posedge clk) begin
        if (exp_17) begin
          exp_104_reg <= exp_103;
        end
      end
      assign exp_104 = exp_104_reg;
      assign exp_103 = {exp_102, exp_69};  assign exp_102 = {exp_101, exp_76};  assign exp_101 = {exp_90, exp_83};  assign exp_89 = exp_94;
  assign exp_94 = 1;
  assign exp_85 = exp_93;
  assign exp_93 = exp_16[31:2];
  assign exp_16 = exp_416;

      reg [31:0] exp_416_reg = 0;
      always@(posedge clk) begin
        if (exp_415) begin
          exp_416_reg <= exp_1019;
        end
      end
      assign exp_416 = exp_416_reg;
    
  reg [32:0] exp_1019_reg;
  always@(*) begin
    case (exp_1015)
      0:exp_1019_reg <= exp_1017;
      1:exp_1019_reg <= exp_748;
      default:exp_1019_reg <= exp_1018;
    endcase
  end
  assign exp_1019 = exp_1019_reg;
  assign exp_1015 = exp_711 & exp_414;
  assign exp_711 = exp_689 | exp_710;
  assign exp_689 = exp_547 | exp_549;
  assign exp_547 = exp_536 == exp_546;
  assign exp_546 = 111;
  assign exp_549 = exp_536 == exp_548;
  assign exp_548 = 103;

  reg [0:0] exp_710_reg;
  always@(*) begin
    case (exp_555)
      0:exp_710_reg <= exp_708;
      1:exp_710_reg <= exp_707;
      default:exp_710_reg <= exp_709;
    endcase
  end
  assign exp_710 = exp_710_reg;
  assign exp_555 = exp_536 == exp_554;
  assign exp_554 = 99;
  assign exp_709 = 0;
  assign exp_708 = 0;

  reg [0:0] exp_707_reg;
  always@(*) begin
    case (exp_537)
      0:exp_707_reg <= exp_690;
      1:exp_707_reg <= exp_691;
      2:exp_707_reg <= exp_704;
      3:exp_707_reg <= exp_705;
      4:exp_707_reg <= exp_692;
      5:exp_707_reg <= exp_693;
      6:exp_707_reg <= exp_698;
      7:exp_707_reg <= exp_703;
      default:exp_707_reg <= exp_706;
    endcase
  end
  assign exp_707 = exp_707_reg;
  assign exp_537 = exp_534[14:12];
  assign exp_706 = 0;
  assign exp_690 = exp_526 == exp_527;

      reg [31:0] exp_526_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_526_reg <= exp_464;
        end
      end
      assign exp_526 = exp_526_reg;
    
  reg [31:0] exp_464_reg;
  always@(*) begin
    case (exp_460)
      0:exp_464_reg <= exp_456;
      1:exp_464_reg <= exp_462;
      default:exp_464_reg <= exp_463;
    endcase
  end
  assign exp_464 = exp_464_reg;
  assign exp_460 = exp_440 == exp_459;
  assign exp_440 = exp_104[19:15];
  assign exp_459 = 0;
  assign exp_463 = 0;

  reg [31:0] exp_456_reg;
  always@(*) begin
    case (exp_437)
      0:exp_456_reg <= exp_427;
      1:exp_456_reg <= exp_439;
      default:exp_456_reg <= exp_455;
    endcase
  end
  assign exp_456 = exp_456_reg;
  assign exp_437 = exp_1010;
  assign exp_1010 = exp_1009 & exp_406;
  assign exp_1009 = exp_1008 & exp_414;
  assign exp_1008 = exp_1007 & exp_1001;
  assign exp_1007 = exp_419 == exp_1002;
  assign exp_419 = exp_104[19:15];
  assign exp_1002 = exp_534[11:7];
  assign exp_1001 = exp_593 | exp_996;
  assign exp_593 = exp_592 | exp_551;
  assign exp_592 = exp_591 | exp_545;
  assign exp_591 = exp_590 | exp_543;
  assign exp_590 = exp_589 | exp_549;
  assign exp_589 = exp_588 | exp_547;
  assign exp_588 = exp_539 | exp_541;
  assign exp_539 = exp_536 == exp_538;
  assign exp_538 = 19;
  assign exp_541 = exp_536 == exp_540;
  assign exp_540 = 51;
  assign exp_543 = exp_536 == exp_542;
  assign exp_542 = 55;
  assign exp_545 = exp_536 == exp_544;
  assign exp_544 = 23;
  assign exp_996 = exp_995 & exp_755;

  reg [0:0] exp_995_reg;
  always@(*) begin
    case (exp_781)
      0:exp_995_reg <= exp_992;
      1:exp_995_reg <= exp_993;
      default:exp_995_reg <= exp_994;
    endcase
  end
  assign exp_995 = exp_995_reg;
  assign exp_781 = exp_755 & exp_780;
  assign exp_755 = exp_753 & exp_754;
  assign exp_753 = exp_751 == exp_752;
  assign exp_751 = exp_534[6:0];
  assign exp_752 = 51;
  assign exp_754 = exp_534[25:25];
  assign exp_780 = exp_750[2:2];
  assign exp_750 = exp_534[14:12];
  assign exp_994 = 0;
  assign exp_992 = exp_985 & exp_755;
  assign exp_985 = exp_900 == exp_984;

      reg [2:0] exp_900_reg = 0;
      always@(posedge clk) begin
        if (exp_896) begin
          exp_900_reg <= exp_907;
        end
      end
      assign exp_900 = exp_900_reg;
    
  reg [2:0] exp_907_reg;
  always@(*) begin
    case (exp_902)
      0:exp_907_reg <= exp_904;
      1:exp_907_reg <= exp_905;
      default:exp_907_reg <= exp_906;
    endcase
  end
  assign exp_907 = exp_907_reg;
  assign exp_902 = exp_900 == exp_901;
  assign exp_901 = 4;
  assign exp_906 = 0;
  assign exp_904 = exp_900 + exp_903;
  assign exp_903 = 1;
  assign exp_905 = 0;
  assign exp_896 = exp_755 & exp_895;
  assign exp_895 = ~exp_894;
  assign exp_894 = exp_750[2:2];
  assign exp_984 = 4;
  assign exp_993 = exp_803 & exp_755;
  assign exp_803 = exp_787 == exp_802;

      reg [5:0] exp_787_reg = 0;
      always@(posedge clk) begin
        if (exp_781) begin
          exp_787_reg <= exp_794;
        end
      end
      assign exp_787 = exp_787_reg;
    
  reg [5:0] exp_794_reg;
  always@(*) begin
    case (exp_789)
      0:exp_794_reg <= exp_791;
      1:exp_794_reg <= exp_792;
      default:exp_794_reg <= exp_793;
    endcase
  end
  assign exp_794 = exp_794_reg;
  assign exp_789 = exp_787 == exp_788;
  assign exp_788 = 37;
  assign exp_793 = 0;
  assign exp_791 = exp_787 + exp_790;
  assign exp_790 = 1;
  assign exp_792 = 0;
  assign exp_802 = 37;

      reg [0:0] exp_414_reg = 0;
      always@(posedge clk) begin
        if (exp_406) begin
          exp_414_reg <= exp_413;
        end
      end
      assign exp_414 = exp_414_reg;
      assign exp_413 = exp_411 & exp_412;

      reg [0:0] exp_411_reg = 0;
      always@(posedge clk) begin
        if (exp_406) begin
          exp_411_reg <= exp_410;
        end
      end
      assign exp_411 = exp_411_reg;
      assign exp_410 = exp_408 & exp_409;
  assign exp_408 = 1;
  assign exp_409 = ~exp_407;
  assign exp_407 = exp_1020;
  assign exp_1020 = exp_414 & exp_711;
  assign exp_406 = ~exp_405;
  assign exp_405 = exp_1024;
  assign exp_1024 = exp_414 & exp_1023;
  assign exp_1023 = exp_1022 | exp_998;
  assign exp_1022 = exp_402 & exp_1021;
  assign exp_1021 = ~exp_401;
  assign exp_401 = exp_393;
  assign exp_393 = exp_291 | exp_392;
  assign exp_291 = exp_204 | exp_290;
  assign exp_204 = exp_163 | exp_203;
  assign exp_163 = exp_34 | exp_162;
  assign exp_34 = exp_15 | exp_33;
  assign exp_15 = 0;
  assign exp_33 = exp_29 & exp_21;
  assign exp_29 = exp_26 & exp_28;
  assign exp_26 = exp_9 >= exp_25;
  assign exp_9 = exp_398;
  assign exp_398 = exp_605;
  assign exp_605 = exp_604 + exp_603;
  assign exp_604 = 0;
  assign exp_603 = exp_526 + exp_602;
  assign exp_602 = $signed(exp_601);
  assign exp_601 = exp_600 + exp_599;
  assign exp_600 = 0;

  reg [11:0] exp_599_reg;
  always@(*) begin
    case (exp_553)
      0:exp_599_reg <= exp_594;
      1:exp_599_reg <= exp_597;
      default:exp_599_reg <= exp_598;
    endcase
  end
  assign exp_599 = exp_599_reg;
  assign exp_553 = exp_536 == exp_552;
  assign exp_552 = 35;
  assign exp_598 = 0;
  assign exp_594 = exp_534[31:20];
  assign exp_597 = {exp_595, exp_596};  assign exp_595 = exp_534[31:25];
  assign exp_596 = exp_534[11:7];
  assign exp_25 = 0;
  assign exp_28 = exp_9 <= exp_27;
  assign exp_27 = 20476;
  assign exp_21 = exp_146;

  reg [0:0] exp_146_reg;
  always@(*) begin
    case (exp_23)
      0:exp_146_reg <= exp_140;
      1:exp_146_reg <= exp_125;
      default:exp_146_reg <= exp_145;
    endcase
  end
  assign exp_146 = exp_146_reg;
  assign exp_23 = exp_12;
  assign exp_12 = exp_403;
  assign exp_403 = exp_688;
  assign exp_688 = exp_687 + exp_553;
  assign exp_687 = 0;
  assign exp_145 = 0;

      reg [0:0] exp_140_reg = 0;
      always@(posedge clk) begin
        if (exp_139) begin
          exp_140_reg <= exp_144;
        end
      end
      assign exp_140 = exp_140_reg;
      assign exp_144 = exp_142 & exp_143;
  assign exp_142 = exp_22 & exp_141;
  assign exp_22 = exp_30;
  assign exp_30 = exp_11 & exp_29;
  assign exp_141 = ~exp_23;
  assign exp_143 = ~exp_140;
  assign exp_139 = 1;
  assign exp_125 = 1;
  assign exp_162 = exp_158 & exp_150;
  assign exp_158 = exp_155 & exp_157;
  assign exp_155 = exp_9 >= exp_154;
  assign exp_154 = 2147483648;
  assign exp_157 = exp_9 <= exp_156;
  assign exp_156 = 2147483652;
  assign exp_150 = exp_184;
  assign exp_184 = 1;
  assign exp_203 = exp_199 & exp_191;
  assign exp_199 = exp_196 & exp_198;
  assign exp_196 = exp_9 >= exp_195;
  assign exp_195 = 2147483656;
  assign exp_198 = exp_9 <= exp_197;
  assign exp_197 = 2147483656;
  assign exp_191 = exp_261;

      reg [0:0] exp_261_reg = 0;
      always@(posedge clk) begin
        if (exp_260) begin
          exp_261_reg <= exp_266;
        end
      end
      assign exp_261 = exp_261_reg;
      assign exp_266 = exp_263 | exp_265;
  assign exp_263 = exp_262 & exp_254;
  assign exp_262 = exp_235 & exp_244;

      reg [0:0] exp_235_reg = 0;
      always@(posedge clk) begin
        if (exp_234) begin
          exp_235_reg <= exp_259;
        end
      end
      assign exp_235 = exp_235_reg;
      assign exp_259 = exp_255 | exp_258;
  assign exp_255 = exp_219 & exp_228;

      reg [0:0] exp_219_reg = 0;
      always@(posedge clk) begin
        if (exp_218) begin
          exp_219_reg <= exp_233;
        end
      end
      assign exp_219 = exp_219_reg;
      assign exp_233 = exp_230 | exp_232;
  assign exp_230 = exp_215 & exp_229;

      reg [0:0] exp_215_reg = 1;
      always@(posedge clk) begin
        if (exp_214) begin
          exp_215_reg <= exp_217;
        end
      end
      assign exp_215 = exp_215_reg;
      assign exp_217 = exp_213 | exp_216;
  assign exp_213 = exp_267;
  assign exp_267 = exp_261 & exp_206;
  assign exp_206 = exp_192 & exp_205;
  assign exp_192 = exp_200;
  assign exp_200 = exp_11 & exp_199;
  assign exp_205 = ~exp_193;
  assign exp_193 = exp_12;
  assign exp_216 = exp_215 & exp_212;

      reg [0:0] exp_212_reg = 1;
      always@(posedge clk) begin
        if (exp_211) begin
          exp_212_reg <= exp_210;
        end
      end
      assign exp_212 = exp_212_reg;
    
      reg [0:0] exp_210_reg = 1;
      always@(posedge clk) begin
        if (exp_209) begin
          exp_210_reg <= exp_208;
        end
      end
      assign exp_210 = exp_210_reg;
    
      reg [0:0] exp_208_reg = 1;
      always@(posedge clk) begin
        if (exp_207) begin
          exp_208_reg <= exp_7;
        end
      end
      assign exp_208 = exp_208_reg;
      assign exp_7 = stdin_rx;
  assign exp_207 = 1;
  assign exp_209 = 1;
  assign exp_211 = 1;
  assign exp_214 = 1;
  assign exp_229 = ~exp_212;
  assign exp_232 = exp_219 & exp_231;
  assign exp_231 = ~exp_228;
  assign exp_228 = exp_222 & exp_219;
  assign exp_222 = exp_220 == exp_221;

      reg [9:0] exp_220_reg = 0;
      always@(posedge clk) begin
        if (exp_219) begin
          exp_220_reg <= exp_227;
        end
      end
      assign exp_220 = exp_220_reg;
    
  reg [9:0] exp_227_reg;
  always@(*) begin
    case (exp_222)
      0:exp_227_reg <= exp_224;
      1:exp_227_reg <= exp_225;
      default:exp_227_reg <= exp_226;
    endcase
  end
  assign exp_227 = exp_227_reg;
  assign exp_226 = 0;
  assign exp_224 = exp_220 + exp_223;
  assign exp_223 = 1;
  assign exp_225 = 0;
  assign exp_221 = 649;
  assign exp_218 = 1;
  assign exp_258 = exp_235 & exp_257;
  assign exp_257 = ~exp_256;
  assign exp_256 = exp_244 & exp_254;
  assign exp_244 = exp_238 & exp_235;
  assign exp_238 = exp_236 == exp_237;

      reg [8:0] exp_236_reg = 0;
      always@(posedge clk) begin
        if (exp_235) begin
          exp_236_reg <= exp_243;
        end
      end
      assign exp_236 = exp_236_reg;
    
  reg [8:0] exp_243_reg;
  always@(*) begin
    case (exp_238)
      0:exp_243_reg <= exp_240;
      1:exp_243_reg <= exp_241;
      default:exp_243_reg <= exp_242;
    endcase
  end
  assign exp_243 = exp_243_reg;
  assign exp_242 = 0;
  assign exp_240 = exp_236 + exp_239;
  assign exp_239 = 1;
  assign exp_241 = 0;
  assign exp_237 = 433;
  assign exp_254 = exp_248 & exp_245;
  assign exp_248 = exp_246 == exp_247;

      reg [2:0] exp_246_reg = 0;
      always@(posedge clk) begin
        if (exp_245) begin
          exp_246_reg <= exp_253;
        end
      end
      assign exp_246 = exp_246_reg;
    
  reg [2:0] exp_253_reg;
  always@(*) begin
    case (exp_248)
      0:exp_253_reg <= exp_250;
      1:exp_253_reg <= exp_251;
      default:exp_253_reg <= exp_252;
    endcase
  end
  assign exp_253 = exp_253_reg;
  assign exp_252 = 0;
  assign exp_250 = exp_246 + exp_249;
  assign exp_249 = 1;
  assign exp_251 = 0;
  assign exp_245 = exp_235 & exp_244;
  assign exp_247 = 7;
  assign exp_234 = 1;
  assign exp_265 = exp_261 & exp_264;
  assign exp_264 = ~exp_206;
  assign exp_260 = 1;
  assign exp_290 = exp_286 & exp_278;
  assign exp_286 = exp_283 & exp_285;
  assign exp_283 = exp_9 >= exp_282;
  assign exp_282 = 2147483660;
  assign exp_285 = exp_9 <= exp_284;
  assign exp_284 = 2147483660;
  assign exp_278 = exp_296;
  assign exp_392 = exp_388 & exp_380;
  assign exp_388 = exp_385 & exp_387;
  assign exp_385 = exp_9 >= exp_384;
  assign exp_384 = 2147483664;
  assign exp_387 = exp_9 <= exp_386;
  assign exp_386 = 2147483664;
  assign exp_380 = exp_397;
  assign exp_397 = 1;
  assign exp_998 = exp_755 & exp_997;
  assign exp_997 = ~exp_995;
  assign exp_412 = ~exp_407;
  assign exp_455 = 0;

  //Create RAM
  reg [31:0] exp_427_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_425) begin
      exp_427_ram[exp_421] <= exp_423;
    end
  end
  assign exp_427 = exp_427_ram[exp_422];
  assign exp_426 = exp_435;
  assign exp_435 = 1;
  assign exp_422 = exp_419;
  assign exp_425 = exp_1004;
  assign exp_1004 = exp_1003 & exp_406;
  assign exp_1003 = exp_1001 & exp_414;
  assign exp_421 = exp_1002;
  assign exp_423 = exp_1000;

  reg [31:0] exp_1000_reg;
  always@(*) begin
    case (exp_996)
      0:exp_1000_reg <= exp_636;
      1:exp_1000_reg <= exp_991;
      default:exp_1000_reg <= exp_999;
    endcase
  end
  assign exp_1000 = exp_1000_reg;
  assign exp_999 = 0;

  reg [31:0] exp_636_reg;
  always@(*) begin
    case (exp_551)
      0:exp_636_reg <= exp_587;
      1:exp_636_reg <= exp_634;
      default:exp_636_reg <= exp_635;
    endcase
  end
  assign exp_636 = exp_636_reg;
  assign exp_635 = 0;

  reg [31:0] exp_587_reg;
  always@(*) begin
    case (exp_530)
      0:exp_587_reg <= exp_566;
      1:exp_587_reg <= exp_568;
      2:exp_587_reg <= exp_584;
      3:exp_587_reg <= exp_585;
      4:exp_587_reg <= exp_577;
      5:exp_587_reg <= exp_581;
      6:exp_587_reg <= exp_582;
      7:exp_587_reg <= exp_583;
      default:exp_587_reg <= exp_586;
    endcase
  end
  assign exp_587 = exp_587_reg;

      reg [2:0] exp_530_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_530_reg <= exp_521;
        end
      end
      assign exp_530 = exp_530_reg;
    
  reg [2:0] exp_521_reg;
  always@(*) begin
    case (exp_518)
      0:exp_521_reg <= exp_508;
      1:exp_521_reg <= exp_519;
      default:exp_521_reg <= exp_520;
    endcase
  end
  assign exp_521 = exp_521_reg;
  assign exp_518 = exp_452 | exp_454;
  assign exp_452 = exp_442 == exp_451;
  assign exp_442 = exp_104[6:0];
  assign exp_451 = 111;
  assign exp_454 = exp_442 == exp_453;
  assign exp_453 = 103;
  assign exp_520 = 0;

  reg [2:0] exp_508_reg;
  always@(*) begin
    case (exp_450)
      0:exp_508_reg <= exp_495;
      1:exp_508_reg <= exp_506;
      default:exp_508_reg <= exp_507;
    endcase
  end
  assign exp_508 = exp_508_reg;
  assign exp_450 = exp_442 == exp_449;
  assign exp_449 = 23;
  assign exp_507 = 0;

  reg [2:0] exp_495_reg;
  always@(*) begin
    case (exp_448)
      0:exp_495_reg <= exp_444;
      1:exp_495_reg <= exp_493;
      default:exp_495_reg <= exp_494;
    endcase
  end
  assign exp_495 = exp_495_reg;
  assign exp_448 = exp_442 == exp_447;
  assign exp_447 = 55;
  assign exp_494 = 0;
  assign exp_444 = exp_104[14:12];
  assign exp_493 = 0;
  assign exp_506 = 0;
  assign exp_519 = 0;
  assign exp_525 = exp_406 & exp_411;
  assign exp_586 = 0;

  reg [31:0] exp_566_reg;
  always@(*) begin
    case (exp_532)
      0:exp_566_reg <= exp_563;
      1:exp_566_reg <= exp_564;
      default:exp_566_reg <= exp_565;
    endcase
  end
  assign exp_566 = exp_566_reg;

      reg [0:0] exp_532_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_532_reg <= exp_524;
        end
      end
      assign exp_532 = exp_532_reg;
      assign exp_524 = exp_510 & exp_523;
  assign exp_510 = exp_497 & exp_509;
  assign exp_497 = exp_483 & exp_496;
  assign exp_483 = exp_481 & exp_482;
  assign exp_481 = exp_104[30:30];
  assign exp_482 = ~exp_446;
  assign exp_446 = exp_442 == exp_445;
  assign exp_445 = 19;
  assign exp_496 = ~exp_448;
  assign exp_509 = ~exp_450;
  assign exp_523 = ~exp_522;
  assign exp_522 = exp_452 | exp_454;
  assign exp_565 = 0;
  assign exp_563 = exp_528 + exp_529;

      reg [31:0] exp_528_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_528_reg <= exp_514;
        end
      end
      assign exp_528 = exp_528_reg;
    
  reg [31:0] exp_514_reg;
  always@(*) begin
    case (exp_511)
      0:exp_514_reg <= exp_503;
      1:exp_514_reg <= exp_512;
      default:exp_514_reg <= exp_513;
    endcase
  end
  assign exp_514 = exp_514_reg;
  assign exp_511 = exp_452 | exp_454;
  assign exp_513 = 0;

  reg [31:0] exp_503_reg;
  always@(*) begin
    case (exp_450)
      0:exp_503_reg <= exp_489;
      1:exp_503_reg <= exp_501;
      default:exp_503_reg <= exp_502;
    endcase
  end
  assign exp_503 = exp_503_reg;
  assign exp_502 = 0;

  reg [31:0] exp_489_reg;
  always@(*) begin
    case (exp_448)
      0:exp_489_reg <= exp_464;
      1:exp_489_reg <= exp_487;
      default:exp_489_reg <= exp_488;
    endcase
  end
  assign exp_489 = exp_489_reg;
  assign exp_488 = 0;
  assign exp_487 = exp_485 << exp_486;
  assign exp_485 = exp_484;
  assign exp_484 = exp_104[31:12];
  assign exp_486 = 12;
  assign exp_501 = exp_499 << exp_500;
  assign exp_499 = exp_498;
  assign exp_498 = exp_104[31:12];
  assign exp_500 = 12;
  assign exp_512 = 4;

      reg [31:0] exp_529_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_529_reg <= exp_517;
        end
      end
      assign exp_529 = exp_529_reg;
    
  reg [31:0] exp_517_reg;
  always@(*) begin
    case (exp_515)
      0:exp_517_reg <= exp_505;
      1:exp_517_reg <= exp_418;
      default:exp_517_reg <= exp_516;
    endcase
  end
  assign exp_517 = exp_517_reg;
  assign exp_515 = exp_452 | exp_454;
  assign exp_516 = 0;

  reg [31:0] exp_505_reg;
  always@(*) begin
    case (exp_450)
      0:exp_505_reg <= exp_492;
      1:exp_505_reg <= exp_418;
      default:exp_505_reg <= exp_504;
    endcase
  end
  assign exp_505 = exp_505_reg;
  assign exp_504 = 0;

  reg [31:0] exp_492_reg;
  always@(*) begin
    case (exp_448)
      0:exp_492_reg <= exp_476;
      1:exp_492_reg <= exp_490;
      default:exp_492_reg <= exp_491;
    endcase
  end
  assign exp_492 = exp_492_reg;
  assign exp_491 = 0;

  reg [31:0] exp_476_reg;
  always@(*) begin
    case (exp_446)
      0:exp_476_reg <= exp_470;
      1:exp_476_reg <= exp_474;
      default:exp_476_reg <= exp_475;
    endcase
  end
  assign exp_476 = exp_476_reg;
  assign exp_475 = 0;

  reg [31:0] exp_470_reg;
  always@(*) begin
    case (exp_466)
      0:exp_470_reg <= exp_458;
      1:exp_470_reg <= exp_468;
      default:exp_470_reg <= exp_469;
    endcase
  end
  assign exp_470 = exp_470_reg;
  assign exp_466 = exp_441 == exp_465;
  assign exp_441 = exp_104[24:20];
  assign exp_465 = 0;
  assign exp_469 = 0;

  reg [31:0] exp_458_reg;
  always@(*) begin
    case (exp_438)
      0:exp_458_reg <= exp_434;
      1:exp_458_reg <= exp_439;
      default:exp_458_reg <= exp_457;
    endcase
  end
  assign exp_458 = exp_458_reg;
  assign exp_438 = exp_1014;
  assign exp_1014 = exp_1013 & exp_406;
  assign exp_1013 = exp_1012 & exp_414;
  assign exp_1012 = exp_1011 & exp_1001;
  assign exp_1011 = exp_420 == exp_1002;
  assign exp_420 = exp_104[24:20];
  assign exp_457 = 0;

  //Create RAM
  reg [31:0] exp_434_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_432) begin
      exp_434_ram[exp_428] <= exp_430;
    end
  end
  assign exp_434 = exp_434_ram[exp_429];
  assign exp_433 = exp_436;
  assign exp_436 = 1;
  assign exp_429 = exp_420;
  assign exp_432 = exp_1006;
  assign exp_1006 = exp_1005 & exp_406;
  assign exp_1005 = exp_1001 & exp_414;
  assign exp_428 = exp_1002;
  assign exp_430 = exp_1000;
  assign exp_439 = exp_1000;
  assign exp_468 = $signed(exp_467);
  assign exp_467 = 0;
  assign exp_474 = exp_471 + exp_473;
  assign exp_471 = 0;
  assign exp_473 = $signed(exp_472);
  assign exp_472 = exp_104[31:20];
  assign exp_490 = 0;

      reg [31:0] exp_418_reg = 0;
      always@(posedge clk) begin
        if (exp_417) begin
          exp_418_reg <= exp_416;
        end
      end
      assign exp_418 = exp_418_reg;
      assign exp_417 = exp_408 & exp_406;
  assign exp_564 = exp_528 - exp_529;
  assign exp_568 = exp_528 << exp_567;
  assign exp_567 = $signed(exp_562);
  assign exp_562 = exp_561 + exp_560;
  assign exp_561 = 0;
  assign exp_560 = exp_531;

      reg [4:0] exp_531_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_531_reg <= exp_480;
        end
      end
      assign exp_531 = exp_531_reg;
    
  reg [4:0] exp_480_reg;
  always@(*) begin
    case (exp_446)
      0:exp_480_reg <= exp_478;
      1:exp_480_reg <= exp_443;
      default:exp_480_reg <= exp_479;
    endcase
  end
  assign exp_480 = exp_480_reg;
  assign exp_479 = 0;
  assign exp_478 = exp_476[4:0];
  assign exp_443 = exp_104[24:20];
  assign exp_584 = $signed(exp_570);
  assign exp_570 = exp_569;
  assign exp_569 = $signed(exp_528) < $signed(exp_529);
  assign exp_585 = $signed(exp_576);
  assign exp_576 = exp_575;
  assign exp_575 = exp_572 < exp_574;
  assign exp_572 = exp_571 + exp_528;
  assign exp_571 = 0;
  assign exp_574 = exp_573 + exp_529;
  assign exp_573 = 0;
  assign exp_577 = exp_528 ^ exp_529;
  assign exp_581 = exp_580[31:0];
  assign exp_580 = $signed(exp_578) >>> $signed(exp_579);
  assign exp_578 = {exp_559, exp_528};
  reg [0:0] exp_559_reg;
  always@(*) begin
    case (exp_533)
      0:exp_559_reg <= exp_557;
      1:exp_559_reg <= exp_556;
      default:exp_559_reg <= exp_558;
    endcase
  end
  assign exp_559 = exp_559_reg;

      reg [0:0] exp_533_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_533_reg <= exp_477;
        end
      end
      assign exp_533 = exp_533_reg;
      assign exp_477 = exp_104[30:30];
  assign exp_558 = 0;
  assign exp_557 = 0;
  assign exp_556 = exp_528[31:31];
  assign exp_579 = $signed(exp_562);
  assign exp_582 = exp_528 | exp_529;
  assign exp_583 = exp_528 & exp_529;

  reg [31:0] exp_634_reg;
  always@(*) begin
    case (exp_537)
      0:exp_634_reg <= exp_624;
      1:exp_634_reg <= exp_627;
      2:exp_634_reg <= exp_400;
      3:exp_634_reg <= exp_628;
      4:exp_634_reg <= exp_629;
      5:exp_634_reg <= exp_630;
      6:exp_634_reg <= exp_631;
      7:exp_634_reg <= exp_632;
      default:exp_634_reg <= exp_633;
    endcase
  end
  assign exp_634 = exp_634_reg;
  assign exp_633 = 0;
  assign exp_624 = $signed(exp_623);
  assign exp_623 = exp_622 + exp_617;
  assign exp_622 = 0;

  reg [7:0] exp_617_reg;
  always@(*) begin
    case (exp_608)
      0:exp_617_reg <= exp_612;
      1:exp_617_reg <= exp_613;
      2:exp_617_reg <= exp_614;
      3:exp_617_reg <= exp_615;
      default:exp_617_reg <= exp_616;
    endcase
  end
  assign exp_617 = exp_617_reg;
  assign exp_608 = exp_607 + exp_606;
  assign exp_607 = 0;
  assign exp_606 = exp_605[1:0];
  assign exp_616 = 0;
  assign exp_612 = exp_400[7:0];
  assign exp_400 = exp_391;

  reg [31:0] exp_391_reg;
  always@(*) begin
    case (exp_388)
      0:exp_391_reg <= exp_289;
      1:exp_391_reg <= exp_379;
      default:exp_391_reg <= exp_390;
    endcase
  end
  assign exp_391 = exp_391_reg;
  assign exp_390 = 0;

  reg [31:0] exp_289_reg;
  always@(*) begin
    case (exp_286)
      0:exp_289_reg <= exp_202;
      1:exp_289_reg <= exp_277;
      default:exp_289_reg <= exp_288;
    endcase
  end
  assign exp_289 = exp_289_reg;
  assign exp_288 = 0;

  reg [31:0] exp_202_reg;
  always@(*) begin
    case (exp_199)
      0:exp_202_reg <= exp_161;
      1:exp_202_reg <= exp_190;
      default:exp_202_reg <= exp_201;
    endcase
  end
  assign exp_202 = exp_202_reg;
  assign exp_201 = 0;

  reg [31:0] exp_161_reg;
  always@(*) begin
    case (exp_158)
      0:exp_161_reg <= exp_32;
      1:exp_161_reg <= exp_149;
      default:exp_161_reg <= exp_160;
    endcase
  end
  assign exp_161 = exp_161_reg;
  assign exp_160 = 0;

  reg [31:0] exp_32_reg;
  always@(*) begin
    case (exp_29)
      0:exp_32_reg <= exp_14;
      1:exp_32_reg <= exp_20;
      default:exp_32_reg <= exp_31;
    endcase
  end
  assign exp_32 = exp_32_reg;
  assign exp_31 = 0;
  assign exp_14 = 0;
  assign exp_20 = exp_127;

      reg [31:0] exp_127_reg = 0;
      always@(posedge clk) begin
        if (exp_126) begin
          exp_127_reg <= exp_138;
        end
      end
      assign exp_127 = exp_127_reg;
      assign exp_138 = {exp_137, exp_41};  assign exp_137 = {exp_136, exp_48};  assign exp_136 = {exp_62, exp_55};
  //Create RAM
  reg [7:0] exp_62_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_62_ram[0] = 0;
    exp_62_ram[1] = 0;
    exp_62_ram[2] = 0;
    exp_62_ram[3] = 0;
    exp_62_ram[4] = 0;
    exp_62_ram[5] = 0;
    exp_62_ram[6] = 0;
    exp_62_ram[7] = 0;
    exp_62_ram[8] = 0;
    exp_62_ram[9] = 0;
    exp_62_ram[10] = 0;
    exp_62_ram[11] = 0;
    exp_62_ram[12] = 0;
    exp_62_ram[13] = 0;
    exp_62_ram[14] = 0;
    exp_62_ram[15] = 0;
    exp_62_ram[16] = 0;
    exp_62_ram[17] = 0;
    exp_62_ram[18] = 0;
    exp_62_ram[19] = 0;
    exp_62_ram[20] = 0;
    exp_62_ram[21] = 0;
    exp_62_ram[22] = 0;
    exp_62_ram[23] = 0;
    exp_62_ram[24] = 0;
    exp_62_ram[25] = 0;
    exp_62_ram[26] = 0;
    exp_62_ram[27] = 0;
    exp_62_ram[28] = 0;
    exp_62_ram[29] = 0;
    exp_62_ram[30] = 0;
    exp_62_ram[31] = 0;
    exp_62_ram[32] = 252;
    exp_62_ram[33] = 113;
    exp_62_ram[34] = 0;
    exp_62_ram[35] = 0;
    exp_62_ram[36] = 0;
    exp_62_ram[37] = 0;
    exp_62_ram[38] = 0;
    exp_62_ram[39] = 0;
    exp_62_ram[40] = 40;
    exp_62_ram[41] = 0;
    exp_62_ram[42] = 165;
    exp_62_ram[43] = 14;
    exp_62_ram[44] = 0;
    exp_62_ram[45] = 12;
    exp_62_ram[46] = 15;
    exp_62_ram[47] = 0;
    exp_62_ram[48] = 0;
    exp_62_ram[49] = 0;
    exp_62_ram[50] = 0;
    exp_62_ram[51] = 0;
    exp_62_ram[52] = 2;
    exp_62_ram[53] = 0;
    exp_62_ram[54] = 64;
    exp_62_ram[55] = 0;
    exp_62_ram[56] = 0;
    exp_62_ram[57] = 0;
    exp_62_ram[58] = 0;
    exp_62_ram[59] = 0;
    exp_62_ram[60] = 0;
    exp_62_ram[61] = 1;
    exp_62_ram[62] = 3;
    exp_62_ram[63] = 1;
    exp_62_ram[64] = 1;
    exp_62_ram[65] = 1;
    exp_62_ram[66] = 3;
    exp_62_ram[67] = 0;
    exp_62_ram[68] = 2;
    exp_62_ram[69] = 1;
    exp_62_ram[70] = 0;
    exp_62_ram[71] = 0;
    exp_62_ram[72] = 1;
    exp_62_ram[73] = 255;
    exp_62_ram[74] = 1;
    exp_62_ram[75] = 0;
    exp_62_ram[76] = 255;
    exp_62_ram[77] = 1;
    exp_62_ram[78] = 64;
    exp_62_ram[79] = 3;
    exp_62_ram[80] = 1;
    exp_62_ram[81] = 1;
    exp_62_ram[82] = 3;
    exp_62_ram[83] = 1;
    exp_62_ram[84] = 0;
    exp_62_ram[85] = 2;
    exp_62_ram[86] = 0;
    exp_62_ram[87] = 0;
    exp_62_ram[88] = 0;
    exp_62_ram[89] = 255;
    exp_62_ram[90] = 1;
    exp_62_ram[91] = 0;
    exp_62_ram[92] = 255;
    exp_62_ram[93] = 1;
    exp_62_ram[94] = 0;
    exp_62_ram[95] = 0;
    exp_62_ram[96] = 14;
    exp_62_ram[97] = 1;
    exp_62_ram[98] = 1;
    exp_62_ram[99] = 242;
    exp_62_ram[100] = 1;
    exp_62_ram[101] = 243;
    exp_62_ram[102] = 0;
    exp_62_ram[103] = 0;
    exp_62_ram[104] = 2;
    exp_62_ram[105] = 0;
    exp_62_ram[106] = 12;
    exp_62_ram[107] = 15;
    exp_62_ram[108] = 1;
    exp_62_ram[109] = 0;
    exp_62_ram[110] = 0;
    exp_62_ram[111] = 0;
    exp_62_ram[112] = 0;
    exp_62_ram[113] = 2;
    exp_62_ram[114] = 0;
    exp_62_ram[115] = 64;
    exp_62_ram[116] = 10;
    exp_62_ram[117] = 65;
    exp_62_ram[118] = 0;
    exp_62_ram[119] = 1;
    exp_62_ram[120] = 1;
    exp_62_ram[121] = 1;
    exp_62_ram[122] = 1;
    exp_62_ram[123] = 3;
    exp_62_ram[124] = 3;
    exp_62_ram[125] = 1;
    exp_62_ram[126] = 0;
    exp_62_ram[127] = 2;
    exp_62_ram[128] = 0;
    exp_62_ram[129] = 1;
    exp_62_ram[130] = 1;
    exp_62_ram[131] = 255;
    exp_62_ram[132] = 1;
    exp_62_ram[133] = 1;
    exp_62_ram[134] = 255;
    exp_62_ram[135] = 1;
    exp_62_ram[136] = 65;
    exp_62_ram[137] = 3;
    exp_62_ram[138] = 1;
    exp_62_ram[139] = 1;
    exp_62_ram[140] = 3;
    exp_62_ram[141] = 1;
    exp_62_ram[142] = 0;
    exp_62_ram[143] = 2;
    exp_62_ram[144] = 0;
    exp_62_ram[145] = 0;
    exp_62_ram[146] = 0;
    exp_62_ram[147] = 255;
    exp_62_ram[148] = 1;
    exp_62_ram[149] = 0;
    exp_62_ram[150] = 255;
    exp_62_ram[151] = 1;
    exp_62_ram[152] = 0;
    exp_62_ram[153] = 0;
    exp_62_ram[154] = 1;
    exp_62_ram[155] = 1;
    exp_62_ram[156] = 244;
    exp_62_ram[157] = 1;
    exp_62_ram[158] = 244;
    exp_62_ram[159] = 0;
    exp_62_ram[160] = 0;
    exp_62_ram[161] = 0;
    exp_62_ram[162] = 0;
    exp_62_ram[163] = 0;
    exp_62_ram[164] = 1;
    exp_62_ram[165] = 0;
    exp_62_ram[166] = 3;
    exp_62_ram[167] = 1;
    exp_62_ram[168] = 1;
    exp_62_ram[169] = 1;
    exp_62_ram[170] = 3;
    exp_62_ram[171] = 1;
    exp_62_ram[172] = 0;
    exp_62_ram[173] = 2;
    exp_62_ram[174] = 0;
    exp_62_ram[175] = 0;
    exp_62_ram[176] = 1;
    exp_62_ram[177] = 255;
    exp_62_ram[178] = 1;
    exp_62_ram[179] = 0;
    exp_62_ram[180] = 255;
    exp_62_ram[181] = 1;
    exp_62_ram[182] = 64;
    exp_62_ram[183] = 3;
    exp_62_ram[184] = 1;
    exp_62_ram[185] = 1;
    exp_62_ram[186] = 3;
    exp_62_ram[187] = 1;
    exp_62_ram[188] = 2;
    exp_62_ram[189] = 0;
    exp_62_ram[190] = 0;
    exp_62_ram[191] = 0;
    exp_62_ram[192] = 1;
    exp_62_ram[193] = 255;
    exp_62_ram[194] = 1;
    exp_62_ram[195] = 0;
    exp_62_ram[196] = 255;
    exp_62_ram[197] = 1;
    exp_62_ram[198] = 1;
    exp_62_ram[199] = 64;
    exp_62_ram[200] = 0;
    exp_62_ram[201] = 235;
    exp_62_ram[202] = 24;
    exp_62_ram[203] = 0;
    exp_62_ram[204] = 4;
    exp_62_ram[205] = 15;
    exp_62_ram[206] = 0;
    exp_62_ram[207] = 0;
    exp_62_ram[208] = 0;
    exp_62_ram[209] = 0;
    exp_62_ram[210] = 165;
    exp_62_ram[211] = 0;
    exp_62_ram[212] = 0;
    exp_62_ram[213] = 2;
    exp_62_ram[214] = 0;
    exp_62_ram[215] = 64;
    exp_62_ram[216] = 2;
    exp_62_ram[217] = 0;
    exp_62_ram[218] = 238;
    exp_62_ram[219] = 0;
    exp_62_ram[220] = 0;
    exp_62_ram[221] = 239;
    exp_62_ram[222] = 1;
    exp_62_ram[223] = 1;
    exp_62_ram[224] = 252;
    exp_62_ram[225] = 1;
    exp_62_ram[226] = 251;
    exp_62_ram[227] = 0;
    exp_62_ram[228] = 0;
    exp_62_ram[229] = 0;
    exp_62_ram[230] = 0;
    exp_62_ram[231] = 1;
    exp_62_ram[232] = 3;
    exp_62_ram[233] = 0;
    exp_62_ram[234] = 0;
    exp_62_ram[235] = 0;
    exp_62_ram[236] = 0;
    exp_62_ram[237] = 1;
    exp_62_ram[238] = 1;
    exp_62_ram[239] = 1;
    exp_62_ram[240] = 3;
    exp_62_ram[241] = 1;
    exp_62_ram[242] = 0;
    exp_62_ram[243] = 3;
    exp_62_ram[244] = 0;
    exp_62_ram[245] = 1;
    exp_62_ram[246] = 1;
    exp_62_ram[247] = 255;
    exp_62_ram[248] = 1;
    exp_62_ram[249] = 1;
    exp_62_ram[250] = 255;
    exp_62_ram[251] = 1;
    exp_62_ram[252] = 65;
    exp_62_ram[253] = 3;
    exp_62_ram[254] = 3;
    exp_62_ram[255] = 1;
    exp_62_ram[256] = 2;
    exp_62_ram[257] = 1;
    exp_62_ram[258] = 1;
    exp_62_ram[259] = 0;
    exp_62_ram[260] = 0;
    exp_62_ram[261] = 1;
    exp_62_ram[262] = 1;
    exp_62_ram[263] = 255;
    exp_62_ram[264] = 1;
    exp_62_ram[265] = 1;
    exp_62_ram[266] = 255;
    exp_62_ram[267] = 1;
    exp_62_ram[268] = 1;
    exp_62_ram[269] = 0;
    exp_62_ram[270] = 0;
    exp_62_ram[271] = 255;
    exp_62_ram[272] = 0;
    exp_62_ram[273] = 1;
    exp_62_ram[274] = 0;
    exp_62_ram[275] = 1;
    exp_62_ram[276] = 65;
    exp_62_ram[277] = 2;
    exp_62_ram[278] = 2;
    exp_62_ram[279] = 1;
    exp_62_ram[280] = 2;
    exp_62_ram[281] = 0;
    exp_62_ram[282] = 1;
    exp_62_ram[283] = 2;
    exp_62_ram[284] = 0;
    exp_62_ram[285] = 1;
    exp_62_ram[286] = 1;
    exp_62_ram[287] = 0;
    exp_62_ram[288] = 2;
    exp_62_ram[289] = 206;
    exp_62_ram[290] = 0;
    exp_62_ram[291] = 255;
    exp_62_ram[292] = 0;
    exp_62_ram[293] = 1;
    exp_62_ram[294] = 0;
    exp_62_ram[295] = 0;
    exp_62_ram[296] = 1;
    exp_62_ram[297] = 0;
    exp_62_ram[298] = 218;
    exp_62_ram[299] = 255;
    exp_62_ram[300] = 204;
    exp_62_ram[301] = 0;
    exp_62_ram[302] = 0;
    exp_62_ram[303] = 218;
    exp_62_ram[304] = 0;
    exp_62_ram[305] = 255;
    exp_62_ram[306] = 1;
    exp_62_ram[307] = 0;
    exp_62_ram[308] = 0;
    exp_62_ram[309] = 0;
    exp_62_ram[310] = 127;
    exp_62_ram[311] = 1;
    exp_62_ram[312] = 127;
    exp_62_ram[313] = 1;
    exp_62_ram[314] = 0;
    exp_62_ram[315] = 0;
    exp_62_ram[316] = 127;
    exp_62_ram[317] = 1;
    exp_62_ram[318] = 1;
    exp_62_ram[319] = 0;
    exp_62_ram[320] = 8;
    exp_62_ram[321] = 0;
    exp_62_ram[322] = 0;
    exp_62_ram[323] = 1;
    exp_62_ram[324] = 0;
    exp_62_ram[325] = 254;
    exp_62_ram[326] = 8;
    exp_62_ram[327] = 0;
    exp_62_ram[328] = 0;
    exp_62_ram[329] = 0;
    exp_62_ram[330] = 0;
    exp_62_ram[331] = 4;
    exp_62_ram[332] = 0;
    exp_62_ram[333] = 0;
    exp_62_ram[334] = 3;
    exp_62_ram[335] = 4;
    exp_62_ram[336] = 255;
    exp_62_ram[337] = 0;
    exp_62_ram[338] = 255;
    exp_62_ram[339] = 0;
    exp_62_ram[340] = 0;
    exp_62_ram[341] = 0;
    exp_62_ram[342] = 0;
    exp_62_ram[343] = 254;
    exp_62_ram[344] = 0;
    exp_62_ram[345] = 253;
    exp_62_ram[346] = 2;
    exp_62_ram[347] = 252;
    exp_62_ram[348] = 255;
    exp_62_ram[349] = 0;
    exp_62_ram[350] = 0;
    exp_62_ram[351] = 0;
    exp_62_ram[352] = 0;
    exp_62_ram[353] = 254;
    exp_62_ram[354] = 251;
    exp_62_ram[355] = 252;
    exp_62_ram[356] = 254;
    exp_62_ram[357] = 247;
    exp_62_ram[358] = 248;
    exp_62_ram[359] = 0;
    exp_62_ram[360] = 248;
    exp_62_ram[361] = 255;
    exp_62_ram[362] = 0;
    exp_62_ram[363] = 0;
    exp_62_ram[364] = 0;
    exp_62_ram[365] = 6;
    exp_62_ram[366] = 42;
    exp_62_ram[367] = 65;
    exp_62_ram[368] = 0;
    exp_62_ram[369] = 64;
    exp_62_ram[370] = 4;
    exp_62_ram[371] = 0;
    exp_62_ram[372] = 64;
    exp_62_ram[373] = 1;
    exp_62_ram[374] = 0;
    exp_62_ram[375] = 0;
    exp_62_ram[376] = 0;
    exp_62_ram[377] = 0;
    exp_62_ram[378] = 0;
    exp_62_ram[379] = 0;
    exp_62_ram[380] = 1;
    exp_62_ram[381] = 0;
    exp_62_ram[382] = 0;
    exp_62_ram[383] = 0;
    exp_62_ram[384] = 1;
    exp_62_ram[385] = 0;
    exp_62_ram[386] = 255;
    exp_62_ram[387] = 0;
    exp_62_ram[388] = 0;
    exp_62_ram[389] = 252;
    exp_62_ram[390] = 0;
    exp_62_ram[391] = 0;
    exp_62_ram[392] = 252;
    exp_62_ram[393] = 254;
    exp_62_ram[394] = 0;
    exp_62_ram[395] = 0;
    exp_62_ram[396] = 0;
    exp_62_ram[397] = 1;
    exp_62_ram[398] = 1;
    exp_62_ram[399] = 1;
    exp_62_ram[400] = 0;
    exp_62_ram[401] = 24;
    exp_62_ram[402] = 0;
    exp_62_ram[403] = 0;
    exp_62_ram[404] = 0;
    exp_62_ram[405] = 8;
    exp_62_ram[406] = 0;
    exp_62_ram[407] = 32;
    exp_62_ram[408] = 0;
    exp_62_ram[409] = 67;
    exp_62_ram[410] = 65;
    exp_62_ram[411] = 67;
    exp_62_ram[412] = 9;
    exp_62_ram[413] = 0;
    exp_62_ram[414] = 0;
    exp_62_ram[415] = 3;
    exp_62_ram[416] = 2;
    exp_62_ram[417] = 7;
    exp_62_ram[418] = 2;
    exp_62_ram[419] = 255;
    exp_62_ram[420] = 65;
    exp_62_ram[421] = 0;
    exp_62_ram[422] = 0;
    exp_62_ram[423] = 0;
    exp_62_ram[424] = 0;
    exp_62_ram[425] = 1;
    exp_62_ram[426] = 1;
    exp_62_ram[427] = 0;
    exp_62_ram[428] = 1;
    exp_62_ram[429] = 0;
    exp_62_ram[430] = 0;
    exp_62_ram[431] = 1;
    exp_62_ram[432] = 1;
    exp_62_ram[433] = 0;
    exp_62_ram[434] = 0;
    exp_62_ram[435] = 0;
    exp_62_ram[436] = 0;
    exp_62_ram[437] = 2;
    exp_62_ram[438] = 0;
    exp_62_ram[439] = 24;
    exp_62_ram[440] = 2;
    exp_62_ram[441] = 248;
    exp_62_ram[442] = 253;
    exp_62_ram[443] = 0;
    exp_62_ram[444] = 0;
    exp_62_ram[445] = 251;
    exp_62_ram[446] = 67;
    exp_62_ram[447] = 3;
    exp_62_ram[448] = 3;
    exp_62_ram[449] = 0;
    exp_62_ram[450] = 0;
    exp_62_ram[451] = 17;
    exp_62_ram[452] = 0;
    exp_62_ram[453] = 0;
    exp_62_ram[454] = 0;
    exp_62_ram[455] = 0;
    exp_62_ram[456] = 0;
    exp_62_ram[457] = 65;
    exp_62_ram[458] = 12;
    exp_62_ram[459] = 0;
    exp_62_ram[460] = 0;
    exp_62_ram[461] = 0;
    exp_62_ram[462] = 0;
    exp_62_ram[463] = 0;
    exp_62_ram[464] = 3;
    exp_62_ram[465] = 2;
    exp_62_ram[466] = 9;
    exp_62_ram[467] = 255;
    exp_62_ram[468] = 0;
    exp_62_ram[469] = 2;
    exp_62_ram[470] = 65;
    exp_62_ram[471] = 1;
    exp_62_ram[472] = 0;
    exp_62_ram[473] = 0;
    exp_62_ram[474] = 255;
    exp_62_ram[475] = 255;
    exp_62_ram[476] = 0;
    exp_62_ram[477] = 0;
    exp_62_ram[478] = 2;
    exp_62_ram[479] = 0;
    exp_62_ram[480] = 0;
    exp_62_ram[481] = 0;
    exp_62_ram[482] = 0;
    exp_62_ram[483] = 0;
    exp_62_ram[484] = 0;
    exp_62_ram[485] = 0;
    exp_62_ram[486] = 0;
    exp_62_ram[487] = 0;
    exp_62_ram[488] = 0;
    exp_62_ram[489] = 255;
    exp_62_ram[490] = 255;
    exp_62_ram[491] = 67;
    exp_62_ram[492] = 0;
    exp_62_ram[493] = 65;
    exp_62_ram[494] = 0;
    exp_62_ram[495] = 1;
    exp_62_ram[496] = 0;
    exp_62_ram[497] = 0;
    exp_62_ram[498] = 237;
    exp_62_ram[499] = 253;
    exp_62_ram[500] = 0;
    exp_62_ram[501] = 0;
    exp_62_ram[502] = 249;
    exp_62_ram[503] = 0;
    exp_62_ram[504] = 0;
    exp_62_ram[505] = 0;
    exp_62_ram[506] = 235;
    exp_62_ram[507] = 2;
    exp_62_ram[508] = 2;
    exp_62_ram[509] = 64;
    exp_62_ram[510] = 0;
    exp_62_ram[511] = 254;
    exp_62_ram[512] = 0;
    exp_62_ram[513] = 0;
    exp_62_ram[514] = 0;
    exp_62_ram[515] = 0;
    exp_62_ram[516] = 0;
    exp_62_ram[517] = 0;
    exp_62_ram[518] = 0;
    exp_62_ram[519] = 0;
    exp_62_ram[520] = 254;
    exp_62_ram[521] = 2;
    exp_62_ram[522] = 2;
    exp_62_ram[523] = 64;
    exp_62_ram[524] = 0;
    exp_62_ram[525] = 254;
    exp_62_ram[526] = 0;
    exp_62_ram[527] = 0;
    exp_62_ram[528] = 0;
    exp_62_ram[529] = 0;
    exp_62_ram[530] = 0;
    exp_62_ram[531] = 0;
    exp_62_ram[532] = 0;
    exp_62_ram[533] = 0;
    exp_62_ram[534] = 254;
    exp_62_ram[535] = 0;
    exp_62_ram[536] = 2;
    exp_62_ram[537] = 15;
    exp_62_ram[538] = 0;
    exp_62_ram[539] = 0;
    exp_62_ram[540] = 0;
    exp_62_ram[541] = 2;
    exp_62_ram[542] = 64;
    exp_62_ram[543] = 0;
    exp_62_ram[544] = 165;
    exp_62_ram[545] = 0;
    exp_62_ram[546] = 0;
    exp_62_ram[547] = 64;
    exp_62_ram[548] = 0;
    exp_62_ram[549] = 1;
    exp_62_ram[550] = 1;
    exp_62_ram[551] = 252;
    exp_62_ram[552] = 1;
    exp_62_ram[553] = 252;
    exp_62_ram[554] = 77;
    exp_62_ram[555] = 117;
    exp_62_ram[556] = 100;
    exp_62_ram[557] = 70;
    exp_62_ram[558] = 97;
    exp_62_ram[559] = 0;
    exp_62_ram[560] = 70;
    exp_62_ram[561] = 97;
    exp_62_ram[562] = 114;
    exp_62_ram[563] = 74;
    exp_62_ram[564] = 117;
    exp_62_ram[565] = 103;
    exp_62_ram[566] = 79;
    exp_62_ram[567] = 111;
    exp_62_ram[568] = 99;
    exp_62_ram[569] = 0;
    exp_62_ram[570] = 108;
    exp_62_ram[571] = 111;
    exp_62_ram[572] = 33;
    exp_62_ram[573] = 0;
    exp_62_ram[574] = 110;
    exp_62_ram[575] = 32;
    exp_62_ram[576] = 103;
    exp_62_ram[577] = 114;
    exp_62_ram[578] = 114;
    exp_62_ram[579] = 109;
    exp_62_ram[580] = 46;
    exp_62_ram[581] = 0;
    exp_62_ram[582] = 0;
    exp_62_ram[583] = 51;
    exp_62_ram[584] = 105;
    exp_62_ram[585] = 110;
    exp_62_ram[586] = 101;
    exp_62_ram[587] = 117;
    exp_62_ram[588] = 112;
    exp_62_ram[589] = 115;
    exp_62_ram[590] = 32;
    exp_62_ram[591] = 101;
    exp_62_ram[592] = 100;
    exp_62_ram[593] = 0;
    exp_62_ram[594] = 54;
    exp_62_ram[595] = 105;
    exp_62_ram[596] = 110;
    exp_62_ram[597] = 101;
    exp_62_ram[598] = 117;
    exp_62_ram[599] = 112;
    exp_62_ram[600] = 115;
    exp_62_ram[601] = 32;
    exp_62_ram[602] = 101;
    exp_62_ram[603] = 100;
    exp_62_ram[604] = 0;
    exp_62_ram[605] = 51;
    exp_62_ram[606] = 105;
    exp_62_ram[607] = 110;
    exp_62_ram[608] = 101;
    exp_62_ram[609] = 105;
    exp_62_ram[610] = 101;
    exp_62_ram[611] = 110;
    exp_62_ram[612] = 115;
    exp_62_ram[613] = 110;
    exp_62_ram[614] = 0;
    exp_62_ram[615] = 54;
    exp_62_ram[616] = 105;
    exp_62_ram[617] = 110;
    exp_62_ram[618] = 101;
    exp_62_ram[619] = 105;
    exp_62_ram[620] = 101;
    exp_62_ram[621] = 110;
    exp_62_ram[622] = 115;
    exp_62_ram[623] = 110;
    exp_62_ram[624] = 0;
    exp_62_ram[625] = 114;
    exp_62_ram[626] = 0;
    exp_62_ram[627] = 116;
    exp_62_ram[628] = 0;
    exp_62_ram[629] = 58;
    exp_62_ram[630] = 0;
    exp_62_ram[631] = 114;
    exp_62_ram[632] = 0;
    exp_62_ram[633] = 117;
    exp_62_ram[634] = 10;
    exp_62_ram[635] = 0;
    exp_62_ram[636] = 105;
    exp_62_ram[637] = 86;
    exp_62_ram[638] = 109;
    exp_62_ram[639] = 0;
    exp_62_ram[640] = 32;
    exp_62_ram[641] = 108;
    exp_62_ram[642] = 111;
    exp_62_ram[643] = 10;
    exp_62_ram[644] = 0;
    exp_62_ram[645] = 75;
    exp_62_ram[646] = 104;
    exp_62_ram[647] = 105;
    exp_62_ram[648] = 10;
    exp_62_ram[649] = 0;
    exp_62_ram[650] = 84;
    exp_62_ram[651] = 32;
    exp_62_ram[652] = 116;
    exp_62_ram[653] = 105;
    exp_62_ram[654] = 105;
    exp_62_ram[655] = 0;
    exp_62_ram[656] = 87;
    exp_62_ram[657] = 32;
    exp_62_ram[658] = 99;
    exp_62_ram[659] = 0;
    exp_62_ram[660] = 2;
    exp_62_ram[661] = 3;
    exp_62_ram[662] = 4;
    exp_62_ram[663] = 4;
    exp_62_ram[664] = 5;
    exp_62_ram[665] = 5;
    exp_62_ram[666] = 5;
    exp_62_ram[667] = 5;
    exp_62_ram[668] = 6;
    exp_62_ram[669] = 6;
    exp_62_ram[670] = 6;
    exp_62_ram[671] = 6;
    exp_62_ram[672] = 6;
    exp_62_ram[673] = 6;
    exp_62_ram[674] = 6;
    exp_62_ram[675] = 6;
    exp_62_ram[676] = 7;
    exp_62_ram[677] = 7;
    exp_62_ram[678] = 7;
    exp_62_ram[679] = 7;
    exp_62_ram[680] = 7;
    exp_62_ram[681] = 7;
    exp_62_ram[682] = 7;
    exp_62_ram[683] = 7;
    exp_62_ram[684] = 7;
    exp_62_ram[685] = 7;
    exp_62_ram[686] = 7;
    exp_62_ram[687] = 7;
    exp_62_ram[688] = 7;
    exp_62_ram[689] = 7;
    exp_62_ram[690] = 7;
    exp_62_ram[691] = 7;
    exp_62_ram[692] = 8;
    exp_62_ram[693] = 8;
    exp_62_ram[694] = 8;
    exp_62_ram[695] = 8;
    exp_62_ram[696] = 8;
    exp_62_ram[697] = 8;
    exp_62_ram[698] = 8;
    exp_62_ram[699] = 8;
    exp_62_ram[700] = 8;
    exp_62_ram[701] = 8;
    exp_62_ram[702] = 8;
    exp_62_ram[703] = 8;
    exp_62_ram[704] = 8;
    exp_62_ram[705] = 8;
    exp_62_ram[706] = 8;
    exp_62_ram[707] = 8;
    exp_62_ram[708] = 8;
    exp_62_ram[709] = 8;
    exp_62_ram[710] = 8;
    exp_62_ram[711] = 8;
    exp_62_ram[712] = 8;
    exp_62_ram[713] = 8;
    exp_62_ram[714] = 8;
    exp_62_ram[715] = 8;
    exp_62_ram[716] = 8;
    exp_62_ram[717] = 8;
    exp_62_ram[718] = 8;
    exp_62_ram[719] = 8;
    exp_62_ram[720] = 8;
    exp_62_ram[721] = 8;
    exp_62_ram[722] = 8;
    exp_62_ram[723] = 8;
    exp_62_ram[724] = 253;
    exp_62_ram[725] = 2;
    exp_62_ram[726] = 3;
    exp_62_ram[727] = 252;
    exp_62_ram[728] = 253;
    exp_62_ram[729] = 254;
    exp_62_ram[730] = 254;
    exp_62_ram[731] = 0;
    exp_62_ram[732] = 0;
    exp_62_ram[733] = 2;
    exp_62_ram[734] = 3;
    exp_62_ram[735] = 0;
    exp_62_ram[736] = 253;
    exp_62_ram[737] = 2;
    exp_62_ram[738] = 3;
    exp_62_ram[739] = 252;
    exp_62_ram[740] = 252;
    exp_62_ram[741] = 253;
    exp_62_ram[742] = 254;
    exp_62_ram[743] = 253;
    exp_62_ram[744] = 254;
    exp_62_ram[745] = 0;
    exp_62_ram[746] = 253;
    exp_62_ram[747] = 0;
    exp_62_ram[748] = 2;
    exp_62_ram[749] = 3;
    exp_62_ram[750] = 0;
    exp_62_ram[751] = 255;
    exp_62_ram[752] = 0;
    exp_62_ram[753] = 0;
    exp_62_ram[754] = 1;
    exp_62_ram[755] = 0;
    exp_62_ram[756] = 9;
    exp_62_ram[757] = 0;
    exp_62_ram[758] = 247;
    exp_62_ram[759] = 0;
    exp_62_ram[760] = 0;
    exp_62_ram[761] = 0;
    exp_62_ram[762] = 0;
    exp_62_ram[763] = 1;
    exp_62_ram[764] = 0;
    exp_62_ram[765] = 253;
    exp_62_ram[766] = 2;
    exp_62_ram[767] = 2;
    exp_62_ram[768] = 3;
    exp_62_ram[769] = 252;
    exp_62_ram[770] = 252;
    exp_62_ram[771] = 254;
    exp_62_ram[772] = 2;
    exp_62_ram[773] = 254;
    exp_62_ram[774] = 0;
    exp_62_ram[775] = 254;
    exp_62_ram[776] = 253;
    exp_62_ram[777] = 0;
    exp_62_ram[778] = 0;
    exp_62_ram[779] = 253;
    exp_62_ram[780] = 0;
    exp_62_ram[781] = 244;
    exp_62_ram[782] = 253;
    exp_62_ram[783] = 254;
    exp_62_ram[784] = 0;
    exp_62_ram[785] = 0;
    exp_62_ram[786] = 252;
    exp_62_ram[787] = 254;
    exp_62_ram[788] = 0;
    exp_62_ram[789] = 2;
    exp_62_ram[790] = 2;
    exp_62_ram[791] = 3;
    exp_62_ram[792] = 0;
    exp_62_ram[793] = 254;
    exp_62_ram[794] = 0;
    exp_62_ram[795] = 0;
    exp_62_ram[796] = 2;
    exp_62_ram[797] = 254;
    exp_62_ram[798] = 0;
    exp_62_ram[799] = 9;
    exp_62_ram[800] = 0;
    exp_62_ram[801] = 254;
    exp_62_ram[802] = 246;
    exp_62_ram[803] = 0;
    exp_62_ram[804] = 9;
    exp_62_ram[805] = 0;
    exp_62_ram[806] = 0;
    exp_62_ram[807] = 238;
    exp_62_ram[808] = 0;
    exp_62_ram[809] = 0;
    exp_62_ram[810] = 1;
    exp_62_ram[811] = 1;
    exp_62_ram[812] = 2;
    exp_62_ram[813] = 0;
    exp_62_ram[814] = 254;
    exp_62_ram[815] = 0;
    exp_62_ram[816] = 2;
    exp_62_ram[817] = 0;
    exp_62_ram[818] = 254;
    exp_62_ram[819] = 254;
    exp_62_ram[820] = 254;
    exp_62_ram[821] = 254;
    exp_62_ram[822] = 0;
    exp_62_ram[823] = 1;
    exp_62_ram[824] = 2;
    exp_62_ram[825] = 0;
    exp_62_ram[826] = 254;
    exp_62_ram[827] = 0;
    exp_62_ram[828] = 0;
    exp_62_ram[829] = 2;
    exp_62_ram[830] = 0;
    exp_62_ram[831] = 254;
    exp_62_ram[832] = 254;
    exp_62_ram[833] = 254;
    exp_62_ram[834] = 254;
    exp_62_ram[835] = 254;
    exp_62_ram[836] = 0;
    exp_62_ram[837] = 254;
    exp_62_ram[838] = 0;
    exp_62_ram[839] = 31;
    exp_62_ram[840] = 0;
    exp_62_ram[841] = 1;
    exp_62_ram[842] = 1;
    exp_62_ram[843] = 2;
    exp_62_ram[844] = 0;
    exp_62_ram[845] = 253;
    exp_62_ram[846] = 2;
    exp_62_ram[847] = 3;
    exp_62_ram[848] = 252;
    exp_62_ram[849] = 252;
    exp_62_ram[850] = 253;
    exp_62_ram[851] = 254;
    exp_62_ram[852] = 1;
    exp_62_ram[853] = 254;
    exp_62_ram[854] = 0;
    exp_62_ram[855] = 254;
    exp_62_ram[856] = 254;
    exp_62_ram[857] = 0;
    exp_62_ram[858] = 0;
    exp_62_ram[859] = 253;
    exp_62_ram[860] = 255;
    exp_62_ram[861] = 252;
    exp_62_ram[862] = 252;
    exp_62_ram[863] = 254;
    exp_62_ram[864] = 253;
    exp_62_ram[865] = 64;
    exp_62_ram[866] = 0;
    exp_62_ram[867] = 2;
    exp_62_ram[868] = 3;
    exp_62_ram[869] = 0;
    exp_62_ram[870] = 254;
    exp_62_ram[871] = 0;
    exp_62_ram[872] = 2;
    exp_62_ram[873] = 0;
    exp_62_ram[874] = 254;
    exp_62_ram[875] = 254;
    exp_62_ram[876] = 2;
    exp_62_ram[877] = 0;
    exp_62_ram[878] = 254;
    exp_62_ram[879] = 3;
    exp_62_ram[880] = 0;
    exp_62_ram[881] = 0;
    exp_62_ram[882] = 0;
    exp_62_ram[883] = 0;
    exp_62_ram[884] = 0;
    exp_62_ram[885] = 15;
    exp_62_ram[886] = 0;
    exp_62_ram[887] = 1;
    exp_62_ram[888] = 2;
    exp_62_ram[889] = 0;
    exp_62_ram[890] = 253;
    exp_62_ram[891] = 2;
    exp_62_ram[892] = 2;
    exp_62_ram[893] = 3;
    exp_62_ram[894] = 252;
    exp_62_ram[895] = 254;
    exp_62_ram[896] = 4;
    exp_62_ram[897] = 254;
    exp_62_ram[898] = 0;
    exp_62_ram[899] = 0;
    exp_62_ram[900] = 0;
    exp_62_ram[901] = 0;
    exp_62_ram[902] = 0;
    exp_62_ram[903] = 253;
    exp_62_ram[904] = 0;
    exp_62_ram[905] = 0;
    exp_62_ram[906] = 253;
    exp_62_ram[907] = 0;
    exp_62_ram[908] = 0;
    exp_62_ram[909] = 0;
    exp_62_ram[910] = 253;
    exp_62_ram[911] = 254;
    exp_62_ram[912] = 253;
    exp_62_ram[913] = 0;
    exp_62_ram[914] = 0;
    exp_62_ram[915] = 0;
    exp_62_ram[916] = 244;
    exp_62_ram[917] = 0;
    exp_62_ram[918] = 250;
    exp_62_ram[919] = 254;
    exp_62_ram[920] = 0;
    exp_62_ram[921] = 2;
    exp_62_ram[922] = 2;
    exp_62_ram[923] = 3;
    exp_62_ram[924] = 0;
    exp_62_ram[925] = 252;
    exp_62_ram[926] = 2;
    exp_62_ram[927] = 2;
    exp_62_ram[928] = 4;
    exp_62_ram[929] = 252;
    exp_62_ram[930] = 252;
    exp_62_ram[931] = 252;
    exp_62_ram[932] = 252;
    exp_62_ram[933] = 252;
    exp_62_ram[934] = 252;
    exp_62_ram[935] = 253;
    exp_62_ram[936] = 253;
    exp_62_ram[937] = 253;
    exp_62_ram[938] = 254;
    exp_62_ram[939] = 252;
    exp_62_ram[940] = 0;
    exp_62_ram[941] = 8;
    exp_62_ram[942] = 252;
    exp_62_ram[943] = 0;
    exp_62_ram[944] = 8;
    exp_62_ram[945] = 252;
    exp_62_ram[946] = 254;
    exp_62_ram[947] = 3;
    exp_62_ram[948] = 253;
    exp_62_ram[949] = 0;
    exp_62_ram[950] = 252;
    exp_62_ram[951] = 253;
    exp_62_ram[952] = 253;
    exp_62_ram[953] = 0;
    exp_62_ram[954] = 253;
    exp_62_ram[955] = 2;
    exp_62_ram[956] = 0;
    exp_62_ram[957] = 254;
    exp_62_ram[958] = 0;
    exp_62_ram[959] = 254;
    exp_62_ram[960] = 254;
    exp_62_ram[961] = 252;
    exp_62_ram[962] = 252;
    exp_62_ram[963] = 4;
    exp_62_ram[964] = 252;
    exp_62_ram[965] = 255;
    exp_62_ram[966] = 252;
    exp_62_ram[967] = 252;
    exp_62_ram[968] = 252;
    exp_62_ram[969] = 0;
    exp_62_ram[970] = 0;
    exp_62_ram[971] = 253;
    exp_62_ram[972] = 0;
    exp_62_ram[973] = 252;
    exp_62_ram[974] = 253;
    exp_62_ram[975] = 253;
    exp_62_ram[976] = 0;
    exp_62_ram[977] = 253;
    exp_62_ram[978] = 0;
    exp_62_ram[979] = 252;
    exp_62_ram[980] = 252;
    exp_62_ram[981] = 252;
    exp_62_ram[982] = 0;
    exp_62_ram[983] = 4;
    exp_62_ram[984] = 2;
    exp_62_ram[985] = 253;
    exp_62_ram[986] = 0;
    exp_62_ram[987] = 252;
    exp_62_ram[988] = 253;
    exp_62_ram[989] = 253;
    exp_62_ram[990] = 0;
    exp_62_ram[991] = 253;
    exp_62_ram[992] = 2;
    exp_62_ram[993] = 0;
    exp_62_ram[994] = 253;
    exp_62_ram[995] = 254;
    exp_62_ram[996] = 64;
    exp_62_ram[997] = 252;
    exp_62_ram[998] = 252;
    exp_62_ram[999] = 253;
    exp_62_ram[1000] = 0;
    exp_62_ram[1001] = 3;
    exp_62_ram[1002] = 3;
    exp_62_ram[1003] = 4;
    exp_62_ram[1004] = 0;
    exp_62_ram[1005] = 253;
    exp_62_ram[1006] = 2;
    exp_62_ram[1007] = 2;
    exp_62_ram[1008] = 3;
    exp_62_ram[1009] = 254;
    exp_62_ram[1010] = 254;
    exp_62_ram[1011] = 254;
    exp_62_ram[1012] = 254;
    exp_62_ram[1013] = 252;
    exp_62_ram[1014] = 252;
    exp_62_ram[1015] = 0;
    exp_62_ram[1016] = 253;
    exp_62_ram[1017] = 252;
    exp_62_ram[1018] = 0;
    exp_62_ram[1019] = 0;
    exp_62_ram[1020] = 10;
    exp_62_ram[1021] = 0;
    exp_62_ram[1022] = 4;
    exp_62_ram[1023] = 0;
    exp_62_ram[1024] = 0;
    exp_62_ram[1025] = 4;
    exp_62_ram[1026] = 253;
    exp_62_ram[1027] = 0;
    exp_62_ram[1028] = 0;
    exp_62_ram[1029] = 0;
    exp_62_ram[1030] = 2;
    exp_62_ram[1031] = 0;
    exp_62_ram[1032] = 255;
    exp_62_ram[1033] = 0;
    exp_62_ram[1034] = 2;
    exp_62_ram[1035] = 253;
    exp_62_ram[1036] = 0;
    exp_62_ram[1037] = 252;
    exp_62_ram[1038] = 253;
    exp_62_ram[1039] = 0;
    exp_62_ram[1040] = 3;
    exp_62_ram[1041] = 0;
    exp_62_ram[1042] = 253;
    exp_62_ram[1043] = 0;
    exp_62_ram[1044] = 2;
    exp_62_ram[1045] = 253;
    exp_62_ram[1046] = 1;
    exp_62_ram[1047] = 252;
    exp_62_ram[1048] = 2;
    exp_62_ram[1049] = 253;
    exp_62_ram[1050] = 0;
    exp_62_ram[1051] = 252;
    exp_62_ram[1052] = 253;
    exp_62_ram[1053] = 0;
    exp_62_ram[1054] = 3;
    exp_62_ram[1055] = 0;
    exp_62_ram[1056] = 0;
    exp_62_ram[1057] = 0;
    exp_62_ram[1058] = 0;
    exp_62_ram[1059] = 253;
    exp_62_ram[1060] = 0;
    exp_62_ram[1061] = 0;
    exp_62_ram[1062] = 253;
    exp_62_ram[1063] = 1;
    exp_62_ram[1064] = 252;
    exp_62_ram[1065] = 0;
    exp_62_ram[1066] = 1;
    exp_62_ram[1067] = 20;
    exp_62_ram[1068] = 0;
    exp_62_ram[1069] = 64;
    exp_62_ram[1070] = 4;
    exp_62_ram[1071] = 253;
    exp_62_ram[1072] = 4;
    exp_62_ram[1073] = 253;
    exp_62_ram[1074] = 0;
    exp_62_ram[1075] = 0;
    exp_62_ram[1076] = 253;
    exp_62_ram[1077] = 0;
    exp_62_ram[1078] = 2;
    exp_62_ram[1079] = 253;
    exp_62_ram[1080] = 255;
    exp_62_ram[1081] = 252;
    exp_62_ram[1082] = 253;
    exp_62_ram[1083] = 0;
    exp_62_ram[1084] = 253;
    exp_62_ram[1085] = 1;
    exp_62_ram[1086] = 0;
    exp_62_ram[1087] = 253;
    exp_62_ram[1088] = 255;
    exp_62_ram[1089] = 252;
    exp_62_ram[1090] = 253;
    exp_62_ram[1091] = 1;
    exp_62_ram[1092] = 2;
    exp_62_ram[1093] = 0;
    exp_62_ram[1094] = 2;
    exp_62_ram[1095] = 2;
    exp_62_ram[1096] = 253;
    exp_62_ram[1097] = 1;
    exp_62_ram[1098] = 2;
    exp_62_ram[1099] = 253;
    exp_62_ram[1100] = 0;
    exp_62_ram[1101] = 252;
    exp_62_ram[1102] = 253;
    exp_62_ram[1103] = 0;
    exp_62_ram[1104] = 7;
    exp_62_ram[1105] = 0;
    exp_62_ram[1106] = 7;
    exp_62_ram[1107] = 253;
    exp_62_ram[1108] = 1;
    exp_62_ram[1109] = 2;
    exp_62_ram[1110] = 0;
    exp_62_ram[1111] = 2;
    exp_62_ram[1112] = 2;
    exp_62_ram[1113] = 253;
    exp_62_ram[1114] = 1;
    exp_62_ram[1115] = 2;
    exp_62_ram[1116] = 253;
    exp_62_ram[1117] = 0;
    exp_62_ram[1118] = 252;
    exp_62_ram[1119] = 253;
    exp_62_ram[1120] = 0;
    exp_62_ram[1121] = 5;
    exp_62_ram[1122] = 0;
    exp_62_ram[1123] = 3;
    exp_62_ram[1124] = 253;
    exp_62_ram[1125] = 0;
    exp_62_ram[1126] = 2;
    exp_62_ram[1127] = 253;
    exp_62_ram[1128] = 1;
    exp_62_ram[1129] = 2;
    exp_62_ram[1130] = 253;
    exp_62_ram[1131] = 0;
    exp_62_ram[1132] = 252;
    exp_62_ram[1133] = 253;
    exp_62_ram[1134] = 0;
    exp_62_ram[1135] = 6;
    exp_62_ram[1136] = 0;
    exp_62_ram[1137] = 253;
    exp_62_ram[1138] = 1;
    exp_62_ram[1139] = 2;
    exp_62_ram[1140] = 253;
    exp_62_ram[1141] = 0;
    exp_62_ram[1142] = 252;
    exp_62_ram[1143] = 253;
    exp_62_ram[1144] = 0;
    exp_62_ram[1145] = 3;
    exp_62_ram[1146] = 0;
    exp_62_ram[1147] = 253;
    exp_62_ram[1148] = 1;
    exp_62_ram[1149] = 8;
    exp_62_ram[1150] = 253;
    exp_62_ram[1151] = 2;
    exp_62_ram[1152] = 253;
    exp_62_ram[1153] = 0;
    exp_62_ram[1154] = 252;
    exp_62_ram[1155] = 253;
    exp_62_ram[1156] = 0;
    exp_62_ram[1157] = 2;
    exp_62_ram[1158] = 0;
    exp_62_ram[1159] = 5;
    exp_62_ram[1160] = 0;
    exp_62_ram[1161] = 0;
    exp_62_ram[1162] = 2;
    exp_62_ram[1163] = 253;
    exp_62_ram[1164] = 0;
    exp_62_ram[1165] = 252;
    exp_62_ram[1166] = 253;
    exp_62_ram[1167] = 0;
    exp_62_ram[1168] = 2;
    exp_62_ram[1169] = 0;
    exp_62_ram[1170] = 2;
    exp_62_ram[1171] = 0;
    exp_62_ram[1172] = 0;
    exp_62_ram[1173] = 2;
    exp_62_ram[1174] = 253;
    exp_62_ram[1175] = 0;
    exp_62_ram[1176] = 252;
    exp_62_ram[1177] = 253;
    exp_62_ram[1178] = 0;
    exp_62_ram[1179] = 2;
    exp_62_ram[1180] = 0;
    exp_62_ram[1181] = 0;
    exp_62_ram[1182] = 0;
    exp_62_ram[1183] = 253;
    exp_62_ram[1184] = 253;
    exp_62_ram[1185] = 254;
    exp_62_ram[1186] = 254;
    exp_62_ram[1187] = 254;
    exp_62_ram[1188] = 254;
    exp_62_ram[1189] = 190;
    exp_62_ram[1190] = 0;
    exp_62_ram[1191] = 0;
    exp_62_ram[1192] = 2;
    exp_62_ram[1193] = 2;
    exp_62_ram[1194] = 3;
    exp_62_ram[1195] = 0;
    exp_62_ram[1196] = 249;
    exp_62_ram[1197] = 6;
    exp_62_ram[1198] = 6;
    exp_62_ram[1199] = 7;
    exp_62_ram[1200] = 250;
    exp_62_ram[1201] = 250;
    exp_62_ram[1202] = 250;
    exp_62_ram[1203] = 250;
    exp_62_ram[1204] = 250;
    exp_62_ram[1205] = 251;
    exp_62_ram[1206] = 251;
    exp_62_ram[1207] = 250;
    exp_62_ram[1208] = 254;
    exp_62_ram[1209] = 250;
    exp_62_ram[1210] = 0;
    exp_62_ram[1211] = 0;
    exp_62_ram[1212] = 254;
    exp_62_ram[1213] = 0;
    exp_62_ram[1214] = 0;
    exp_62_ram[1215] = 64;
    exp_62_ram[1216] = 0;
    exp_62_ram[1217] = 250;
    exp_62_ram[1218] = 8;
    exp_62_ram[1219] = 250;
    exp_62_ram[1220] = 250;
    exp_62_ram[1221] = 2;
    exp_62_ram[1222] = 254;
    exp_62_ram[1223] = 254;
    exp_62_ram[1224] = 0;
    exp_62_ram[1225] = 0;
    exp_62_ram[1226] = 254;
    exp_62_ram[1227] = 3;
    exp_62_ram[1228] = 15;
    exp_62_ram[1229] = 3;
    exp_62_ram[1230] = 0;
    exp_62_ram[1231] = 2;
    exp_62_ram[1232] = 0;
    exp_62_ram[1233] = 4;
    exp_62_ram[1234] = 0;
    exp_62_ram[1235] = 6;
    exp_62_ram[1236] = 254;
    exp_62_ram[1237] = 0;
    exp_62_ram[1238] = 15;
    exp_62_ram[1239] = 255;
    exp_62_ram[1240] = 15;
    exp_62_ram[1241] = 254;
    exp_62_ram[1242] = 0;
    exp_62_ram[1243] = 254;
    exp_62_ram[1244] = 255;
    exp_62_ram[1245] = 0;
    exp_62_ram[1246] = 252;
    exp_62_ram[1247] = 250;
    exp_62_ram[1248] = 250;
    exp_62_ram[1249] = 2;
    exp_62_ram[1250] = 250;
    exp_62_ram[1251] = 250;
    exp_62_ram[1252] = 0;
    exp_62_ram[1253] = 254;
    exp_62_ram[1254] = 1;
    exp_62_ram[1255] = 246;
    exp_62_ram[1256] = 250;
    exp_62_ram[1257] = 252;
    exp_62_ram[1258] = 0;
    exp_62_ram[1259] = 0;
    exp_62_ram[1260] = 0;
    exp_62_ram[1261] = 0;
    exp_62_ram[1262] = 250;
    exp_62_ram[1263] = 0;
    exp_62_ram[1264] = 250;
    exp_62_ram[1265] = 0;
    exp_62_ram[1266] = 254;
    exp_62_ram[1267] = 251;
    exp_62_ram[1268] = 251;
    exp_62_ram[1269] = 251;
    exp_62_ram[1270] = 251;
    exp_62_ram[1271] = 189;
    exp_62_ram[1272] = 0;
    exp_62_ram[1273] = 0;
    exp_62_ram[1274] = 6;
    exp_62_ram[1275] = 6;
    exp_62_ram[1276] = 7;
    exp_62_ram[1277] = 0;
    exp_62_ram[1278] = 248;
    exp_62_ram[1279] = 6;
    exp_62_ram[1280] = 6;
    exp_62_ram[1281] = 8;
    exp_62_ram[1282] = 250;
    exp_62_ram[1283] = 250;
    exp_62_ram[1284] = 250;
    exp_62_ram[1285] = 250;
    exp_62_ram[1286] = 248;
    exp_62_ram[1287] = 252;
    exp_62_ram[1288] = 250;
    exp_62_ram[1289] = 32;
    exp_62_ram[1290] = 0;
    exp_62_ram[1291] = 203;
    exp_62_ram[1292] = 250;
    exp_62_ram[1293] = 32;
    exp_62_ram[1294] = 250;
    exp_62_ram[1295] = 0;
    exp_62_ram[1296] = 2;
    exp_62_ram[1297] = 2;
    exp_62_ram[1298] = 250;
    exp_62_ram[1299] = 0;
    exp_62_ram[1300] = 253;
    exp_62_ram[1301] = 0;
    exp_62_ram[1302] = 252;
    exp_62_ram[1303] = 250;
    exp_62_ram[1304] = 250;
    exp_62_ram[1305] = 0;
    exp_62_ram[1306] = 250;
    exp_62_ram[1307] = 0;
    exp_62_ram[1308] = 250;
    exp_62_ram[1309] = 0;
    exp_62_ram[1310] = 250;
    exp_62_ram[1311] = 28;
    exp_62_ram[1312] = 250;
    exp_62_ram[1313] = 0;
    exp_62_ram[1314] = 250;
    exp_62_ram[1315] = 254;
    exp_62_ram[1316] = 250;
    exp_62_ram[1317] = 0;
    exp_62_ram[1318] = 254;
    exp_62_ram[1319] = 1;
    exp_62_ram[1320] = 12;
    exp_62_ram[1321] = 0;
    exp_62_ram[1322] = 0;
    exp_62_ram[1323] = 10;
    exp_62_ram[1324] = 0;
    exp_62_ram[1325] = 0;
    exp_62_ram[1326] = 0;
    exp_62_ram[1327] = 254;
    exp_62_ram[1328] = 0;
    exp_62_ram[1329] = 254;
    exp_62_ram[1330] = 250;
    exp_62_ram[1331] = 0;
    exp_62_ram[1332] = 250;
    exp_62_ram[1333] = 0;
    exp_62_ram[1334] = 254;
    exp_62_ram[1335] = 9;
    exp_62_ram[1336] = 254;
    exp_62_ram[1337] = 0;
    exp_62_ram[1338] = 254;
    exp_62_ram[1339] = 250;
    exp_62_ram[1340] = 0;
    exp_62_ram[1341] = 250;
    exp_62_ram[1342] = 0;
    exp_62_ram[1343] = 254;
    exp_62_ram[1344] = 7;
    exp_62_ram[1345] = 254;
    exp_62_ram[1346] = 0;
    exp_62_ram[1347] = 254;
    exp_62_ram[1348] = 250;
    exp_62_ram[1349] = 0;
    exp_62_ram[1350] = 250;
    exp_62_ram[1351] = 0;
    exp_62_ram[1352] = 254;
    exp_62_ram[1353] = 5;
    exp_62_ram[1354] = 254;
    exp_62_ram[1355] = 0;
    exp_62_ram[1356] = 254;
    exp_62_ram[1357] = 250;
    exp_62_ram[1358] = 0;
    exp_62_ram[1359] = 250;
    exp_62_ram[1360] = 0;
    exp_62_ram[1361] = 254;
    exp_62_ram[1362] = 3;
    exp_62_ram[1363] = 254;
    exp_62_ram[1364] = 1;
    exp_62_ram[1365] = 254;
    exp_62_ram[1366] = 250;
    exp_62_ram[1367] = 0;
    exp_62_ram[1368] = 250;
    exp_62_ram[1369] = 0;
    exp_62_ram[1370] = 254;
    exp_62_ram[1371] = 0;
    exp_62_ram[1372] = 254;
    exp_62_ram[1373] = 0;
    exp_62_ram[1374] = 254;
    exp_62_ram[1375] = 240;
    exp_62_ram[1376] = 254;
    exp_62_ram[1377] = 250;
    exp_62_ram[1378] = 0;
    exp_62_ram[1379] = 0;
    exp_62_ram[1380] = 128;
    exp_62_ram[1381] = 0;
    exp_62_ram[1382] = 0;
    exp_62_ram[1383] = 250;
    exp_62_ram[1384] = 0;
    exp_62_ram[1385] = 132;
    exp_62_ram[1386] = 254;
    exp_62_ram[1387] = 6;
    exp_62_ram[1388] = 250;
    exp_62_ram[1389] = 0;
    exp_62_ram[1390] = 2;
    exp_62_ram[1391] = 4;
    exp_62_ram[1392] = 249;
    exp_62_ram[1393] = 0;
    exp_62_ram[1394] = 248;
    exp_62_ram[1395] = 0;
    exp_62_ram[1396] = 252;
    exp_62_ram[1397] = 252;
    exp_62_ram[1398] = 2;
    exp_62_ram[1399] = 254;
    exp_62_ram[1400] = 0;
    exp_62_ram[1401] = 254;
    exp_62_ram[1402] = 252;
    exp_62_ram[1403] = 64;
    exp_62_ram[1404] = 254;
    exp_62_ram[1405] = 0;
    exp_62_ram[1406] = 252;
    exp_62_ram[1407] = 254;
    exp_62_ram[1408] = 250;
    exp_62_ram[1409] = 0;
    exp_62_ram[1410] = 250;
    exp_62_ram[1411] = 254;
    exp_62_ram[1412] = 250;
    exp_62_ram[1413] = 0;
    exp_62_ram[1414] = 2;
    exp_62_ram[1415] = 8;
    exp_62_ram[1416] = 254;
    exp_62_ram[1417] = 64;
    exp_62_ram[1418] = 254;
    exp_62_ram[1419] = 250;
    exp_62_ram[1420] = 0;
    exp_62_ram[1421] = 250;
    exp_62_ram[1422] = 250;
    exp_62_ram[1423] = 0;
    exp_62_ram[1424] = 0;
    exp_62_ram[1425] = 245;
    exp_62_ram[1426] = 0;
    exp_62_ram[1427] = 0;
    exp_62_ram[1428] = 250;
    exp_62_ram[1429] = 0;
    exp_62_ram[1430] = 249;
    exp_62_ram[1431] = 254;
    exp_62_ram[1432] = 4;
    exp_62_ram[1433] = 250;
    exp_62_ram[1434] = 0;
    exp_62_ram[1435] = 2;
    exp_62_ram[1436] = 2;
    exp_62_ram[1437] = 249;
    exp_62_ram[1438] = 0;
    exp_62_ram[1439] = 248;
    exp_62_ram[1440] = 0;
    exp_62_ram[1441] = 252;
    exp_62_ram[1442] = 252;
    exp_62_ram[1443] = 0;
    exp_62_ram[1444] = 0;
    exp_62_ram[1445] = 254;
    exp_62_ram[1446] = 250;
    exp_62_ram[1447] = 0;
    exp_62_ram[1448] = 250;
    exp_62_ram[1449] = 250;
    exp_62_ram[1450] = 0;
    exp_62_ram[1451] = 249;
    exp_62_ram[1452] = 1;
    exp_62_ram[1453] = 14;
    exp_62_ram[1454] = 0;
    exp_62_ram[1455] = 0;
    exp_62_ram[1456] = 14;
    exp_62_ram[1457] = 0;
    exp_62_ram[1458] = 0;
    exp_62_ram[1459] = 0;
    exp_62_ram[1460] = 254;
    exp_62_ram[1461] = 16;
    exp_62_ram[1462] = 254;
    exp_62_ram[1463] = 250;
    exp_62_ram[1464] = 0;
    exp_62_ram[1465] = 250;
    exp_62_ram[1466] = 250;
    exp_62_ram[1467] = 0;
    exp_62_ram[1468] = 6;
    exp_62_ram[1469] = 12;
    exp_62_ram[1470] = 254;
    exp_62_ram[1471] = 32;
    exp_62_ram[1472] = 254;
    exp_62_ram[1473] = 250;
    exp_62_ram[1474] = 0;
    exp_62_ram[1475] = 250;
    exp_62_ram[1476] = 10;
    exp_62_ram[1477] = 254;
    exp_62_ram[1478] = 8;
    exp_62_ram[1479] = 254;
    exp_62_ram[1480] = 250;
    exp_62_ram[1481] = 0;
    exp_62_ram[1482] = 250;
    exp_62_ram[1483] = 250;
    exp_62_ram[1484] = 0;
    exp_62_ram[1485] = 6;
    exp_62_ram[1486] = 8;
    exp_62_ram[1487] = 254;
    exp_62_ram[1488] = 4;
    exp_62_ram[1489] = 254;
    exp_62_ram[1490] = 250;
    exp_62_ram[1491] = 0;
    exp_62_ram[1492] = 250;
    exp_62_ram[1493] = 6;
    exp_62_ram[1494] = 254;
    exp_62_ram[1495] = 16;
    exp_62_ram[1496] = 254;
    exp_62_ram[1497] = 250;
    exp_62_ram[1498] = 0;
    exp_62_ram[1499] = 250;
    exp_62_ram[1500] = 5;
    exp_62_ram[1501] = 254;
    exp_62_ram[1502] = 32;
    exp_62_ram[1503] = 254;
    exp_62_ram[1504] = 250;
    exp_62_ram[1505] = 0;
    exp_62_ram[1506] = 250;
    exp_62_ram[1507] = 3;
    exp_62_ram[1508] = 254;
    exp_62_ram[1509] = 16;
    exp_62_ram[1510] = 254;
    exp_62_ram[1511] = 250;
    exp_62_ram[1512] = 0;
    exp_62_ram[1513] = 250;
    exp_62_ram[1514] = 1;
    exp_62_ram[1515] = 0;
    exp_62_ram[1516] = 1;
    exp_62_ram[1517] = 0;
    exp_62_ram[1518] = 0;
    exp_62_ram[1519] = 0;
    exp_62_ram[1520] = 250;
    exp_62_ram[1521] = 0;
    exp_62_ram[1522] = 253;
    exp_62_ram[1523] = 5;
    exp_62_ram[1524] = 98;
    exp_62_ram[1525] = 0;
    exp_62_ram[1526] = 0;
    exp_62_ram[1527] = 19;
    exp_62_ram[1528] = 0;
    exp_62_ram[1529] = 0;
    exp_62_ram[1530] = 0;
    exp_62_ram[1531] = 250;
    exp_62_ram[1532] = 0;
    exp_62_ram[1533] = 7;
    exp_62_ram[1534] = 0;
    exp_62_ram[1535] = 250;
    exp_62_ram[1536] = 0;
    exp_62_ram[1537] = 5;
    exp_62_ram[1538] = 0;
    exp_62_ram[1539] = 1;
    exp_62_ram[1540] = 252;
    exp_62_ram[1541] = 5;
    exp_62_ram[1542] = 250;
    exp_62_ram[1543] = 0;
    exp_62_ram[1544] = 6;
    exp_62_ram[1545] = 0;
    exp_62_ram[1546] = 0;
    exp_62_ram[1547] = 252;
    exp_62_ram[1548] = 3;
    exp_62_ram[1549] = 250;
    exp_62_ram[1550] = 0;
    exp_62_ram[1551] = 6;
    exp_62_ram[1552] = 0;
    exp_62_ram[1553] = 0;
    exp_62_ram[1554] = 252;
    exp_62_ram[1555] = 1;
    exp_62_ram[1556] = 0;
    exp_62_ram[1557] = 252;
    exp_62_ram[1558] = 254;
    exp_62_ram[1559] = 254;
    exp_62_ram[1560] = 254;
    exp_62_ram[1561] = 250;
    exp_62_ram[1562] = 0;
    exp_62_ram[1563] = 5;
    exp_62_ram[1564] = 0;
    exp_62_ram[1565] = 254;
    exp_62_ram[1566] = 2;
    exp_62_ram[1567] = 254;
    exp_62_ram[1568] = 250;
    exp_62_ram[1569] = 0;
    exp_62_ram[1570] = 6;
    exp_62_ram[1571] = 2;
    exp_62_ram[1572] = 250;
    exp_62_ram[1573] = 0;
    exp_62_ram[1574] = 6;
    exp_62_ram[1575] = 0;
    exp_62_ram[1576] = 254;
    exp_62_ram[1577] = 255;
    exp_62_ram[1578] = 254;
    exp_62_ram[1579] = 254;
    exp_62_ram[1580] = 64;
    exp_62_ram[1581] = 0;
    exp_62_ram[1582] = 254;
    exp_62_ram[1583] = 255;
    exp_62_ram[1584] = 254;
    exp_62_ram[1585] = 250;
    exp_62_ram[1586] = 0;
    exp_62_ram[1587] = 6;
    exp_62_ram[1588] = 0;
    exp_62_ram[1589] = 250;
    exp_62_ram[1590] = 0;
    exp_62_ram[1591] = 6;
    exp_62_ram[1592] = 20;
    exp_62_ram[1593] = 254;
    exp_62_ram[1594] = 32;
    exp_62_ram[1595] = 34;
    exp_62_ram[1596] = 254;
    exp_62_ram[1597] = 16;
    exp_62_ram[1598] = 6;
    exp_62_ram[1599] = 249;
    exp_62_ram[1600] = 0;
    exp_62_ram[1601] = 248;
    exp_62_ram[1602] = 0;
    exp_62_ram[1603] = 250;
    exp_62_ram[1604] = 251;
    exp_62_ram[1605] = 65;
    exp_62_ram[1606] = 251;
    exp_62_ram[1607] = 0;
    exp_62_ram[1608] = 64;
    exp_62_ram[1609] = 0;
    exp_62_ram[1610] = 251;
    exp_62_ram[1611] = 1;
    exp_62_ram[1612] = 15;
    exp_62_ram[1613] = 254;
    exp_62_ram[1614] = 0;
    exp_62_ram[1615] = 254;
    exp_62_ram[1616] = 0;
    exp_62_ram[1617] = 254;
    exp_62_ram[1618] = 253;
    exp_62_ram[1619] = 0;
    exp_62_ram[1620] = 0;
    exp_62_ram[1621] = 250;
    exp_62_ram[1622] = 253;
    exp_62_ram[1623] = 250;
    exp_62_ram[1624] = 250;
    exp_62_ram[1625] = 148;
    exp_62_ram[1626] = 252;
    exp_62_ram[1627] = 27;
    exp_62_ram[1628] = 254;
    exp_62_ram[1629] = 4;
    exp_62_ram[1630] = 0;
    exp_62_ram[1631] = 249;
    exp_62_ram[1632] = 0;
    exp_62_ram[1633] = 248;
    exp_62_ram[1634] = 0;
    exp_62_ram[1635] = 15;
    exp_62_ram[1636] = 3;
    exp_62_ram[1637] = 254;
    exp_62_ram[1638] = 8;
    exp_62_ram[1639] = 2;
    exp_62_ram[1640] = 249;
    exp_62_ram[1641] = 0;
    exp_62_ram[1642] = 248;
    exp_62_ram[1643] = 0;
    exp_62_ram[1644] = 1;
    exp_62_ram[1645] = 65;
    exp_62_ram[1646] = 1;
    exp_62_ram[1647] = 249;
    exp_62_ram[1648] = 0;
    exp_62_ram[1649] = 248;
    exp_62_ram[1650] = 0;
    exp_62_ram[1651] = 250;
    exp_62_ram[1652] = 251;
    exp_62_ram[1653] = 65;
    exp_62_ram[1654] = 251;
    exp_62_ram[1655] = 0;
    exp_62_ram[1656] = 64;
    exp_62_ram[1657] = 0;
    exp_62_ram[1658] = 251;
    exp_62_ram[1659] = 1;
    exp_62_ram[1660] = 15;
    exp_62_ram[1661] = 254;
    exp_62_ram[1662] = 0;
    exp_62_ram[1663] = 254;
    exp_62_ram[1664] = 0;
    exp_62_ram[1665] = 254;
    exp_62_ram[1666] = 253;
    exp_62_ram[1667] = 0;
    exp_62_ram[1668] = 0;
    exp_62_ram[1669] = 250;
    exp_62_ram[1670] = 253;
    exp_62_ram[1671] = 250;
    exp_62_ram[1672] = 250;
    exp_62_ram[1673] = 136;
    exp_62_ram[1674] = 252;
    exp_62_ram[1675] = 15;
    exp_62_ram[1676] = 254;
    exp_62_ram[1677] = 32;
    exp_62_ram[1678] = 14;
    exp_62_ram[1679] = 254;
    exp_62_ram[1680] = 16;
    exp_62_ram[1681] = 4;
    exp_62_ram[1682] = 249;
    exp_62_ram[1683] = 0;
    exp_62_ram[1684] = 248;
    exp_62_ram[1685] = 0;
    exp_62_ram[1686] = 254;
    exp_62_ram[1687] = 0;
    exp_62_ram[1688] = 254;
    exp_62_ram[1689] = 0;
    exp_62_ram[1690] = 254;
    exp_62_ram[1691] = 253;
    exp_62_ram[1692] = 0;
    exp_62_ram[1693] = 250;
    exp_62_ram[1694] = 253;
    exp_62_ram[1695] = 250;
    exp_62_ram[1696] = 250;
    exp_62_ram[1697] = 130;
    exp_62_ram[1698] = 252;
    exp_62_ram[1699] = 9;
    exp_62_ram[1700] = 254;
    exp_62_ram[1701] = 4;
    exp_62_ram[1702] = 0;
    exp_62_ram[1703] = 249;
    exp_62_ram[1704] = 0;
    exp_62_ram[1705] = 248;
    exp_62_ram[1706] = 0;
    exp_62_ram[1707] = 15;
    exp_62_ram[1708] = 3;
    exp_62_ram[1709] = 254;
    exp_62_ram[1710] = 8;
    exp_62_ram[1711] = 2;
    exp_62_ram[1712] = 249;
    exp_62_ram[1713] = 0;
    exp_62_ram[1714] = 248;
    exp_62_ram[1715] = 0;
    exp_62_ram[1716] = 1;
    exp_62_ram[1717] = 1;
    exp_62_ram[1718] = 1;
    exp_62_ram[1719] = 249;
    exp_62_ram[1720] = 0;
    exp_62_ram[1721] = 248;
    exp_62_ram[1722] = 0;
    exp_62_ram[1723] = 252;
    exp_62_ram[1724] = 254;
    exp_62_ram[1725] = 0;
    exp_62_ram[1726] = 254;
    exp_62_ram[1727] = 0;
    exp_62_ram[1728] = 254;
    exp_62_ram[1729] = 253;
    exp_62_ram[1730] = 0;
    exp_62_ram[1731] = 252;
    exp_62_ram[1732] = 250;
    exp_62_ram[1733] = 253;
    exp_62_ram[1734] = 250;
    exp_62_ram[1735] = 250;
    exp_62_ram[1736] = 249;
    exp_62_ram[1737] = 252;
    exp_62_ram[1738] = 250;
    exp_62_ram[1739] = 0;
    exp_62_ram[1740] = 250;
    exp_62_ram[1741] = 48;
    exp_62_ram[1742] = 0;
    exp_62_ram[1743] = 252;
    exp_62_ram[1744] = 254;
    exp_62_ram[1745] = 0;
    exp_62_ram[1746] = 4;
    exp_62_ram[1747] = 2;
    exp_62_ram[1748] = 253;
    exp_62_ram[1749] = 0;
    exp_62_ram[1750] = 252;
    exp_62_ram[1751] = 250;
    exp_62_ram[1752] = 250;
    exp_62_ram[1753] = 0;
    exp_62_ram[1754] = 250;
    exp_62_ram[1755] = 2;
    exp_62_ram[1756] = 0;
    exp_62_ram[1757] = 253;
    exp_62_ram[1758] = 0;
    exp_62_ram[1759] = 252;
    exp_62_ram[1760] = 254;
    exp_62_ram[1761] = 252;
    exp_62_ram[1762] = 249;
    exp_62_ram[1763] = 0;
    exp_62_ram[1764] = 248;
    exp_62_ram[1765] = 0;
    exp_62_ram[1766] = 15;
    exp_62_ram[1767] = 253;
    exp_62_ram[1768] = 0;
    exp_62_ram[1769] = 252;
    exp_62_ram[1770] = 250;
    exp_62_ram[1771] = 250;
    exp_62_ram[1772] = 0;
    exp_62_ram[1773] = 250;
    exp_62_ram[1774] = 0;
    exp_62_ram[1775] = 254;
    exp_62_ram[1776] = 0;
    exp_62_ram[1777] = 4;
    exp_62_ram[1778] = 2;
    exp_62_ram[1779] = 253;
    exp_62_ram[1780] = 0;
    exp_62_ram[1781] = 252;
    exp_62_ram[1782] = 250;
    exp_62_ram[1783] = 250;
    exp_62_ram[1784] = 0;
    exp_62_ram[1785] = 250;
    exp_62_ram[1786] = 2;
    exp_62_ram[1787] = 0;
    exp_62_ram[1788] = 253;
    exp_62_ram[1789] = 0;
    exp_62_ram[1790] = 252;
    exp_62_ram[1791] = 254;
    exp_62_ram[1792] = 252;
    exp_62_ram[1793] = 250;
    exp_62_ram[1794] = 0;
    exp_62_ram[1795] = 250;
    exp_62_ram[1796] = 35;
    exp_62_ram[1797] = 249;
    exp_62_ram[1798] = 0;
    exp_62_ram[1799] = 248;
    exp_62_ram[1800] = 0;
    exp_62_ram[1801] = 252;
    exp_62_ram[1802] = 254;
    exp_62_ram[1803] = 0;
    exp_62_ram[1804] = 254;
    exp_62_ram[1805] = 0;
    exp_62_ram[1806] = 255;
    exp_62_ram[1807] = 0;
    exp_62_ram[1808] = 253;
    exp_62_ram[1809] = 143;
    exp_62_ram[1810] = 252;
    exp_62_ram[1811] = 254;
    exp_62_ram[1812] = 64;
    exp_62_ram[1813] = 0;
    exp_62_ram[1814] = 252;
    exp_62_ram[1815] = 254;
    exp_62_ram[1816] = 0;
    exp_62_ram[1817] = 0;
    exp_62_ram[1818] = 252;
    exp_62_ram[1819] = 254;
    exp_62_ram[1820] = 0;
    exp_62_ram[1821] = 6;
    exp_62_ram[1822] = 2;
    exp_62_ram[1823] = 253;
    exp_62_ram[1824] = 0;
    exp_62_ram[1825] = 252;
    exp_62_ram[1826] = 250;
    exp_62_ram[1827] = 250;
    exp_62_ram[1828] = 0;
    exp_62_ram[1829] = 250;
    exp_62_ram[1830] = 2;
    exp_62_ram[1831] = 0;
    exp_62_ram[1832] = 252;
    exp_62_ram[1833] = 0;
    exp_62_ram[1834] = 252;
    exp_62_ram[1835] = 254;
    exp_62_ram[1836] = 252;
    exp_62_ram[1837] = 3;
    exp_62_ram[1838] = 253;
    exp_62_ram[1839] = 0;
    exp_62_ram[1840] = 252;
    exp_62_ram[1841] = 0;
    exp_62_ram[1842] = 253;
    exp_62_ram[1843] = 0;
    exp_62_ram[1844] = 252;
    exp_62_ram[1845] = 250;
    exp_62_ram[1846] = 250;
    exp_62_ram[1847] = 0;
    exp_62_ram[1848] = 250;
    exp_62_ram[1849] = 0;
    exp_62_ram[1850] = 253;
    exp_62_ram[1851] = 0;
    exp_62_ram[1852] = 2;
    exp_62_ram[1853] = 254;
    exp_62_ram[1854] = 64;
    exp_62_ram[1855] = 250;
    exp_62_ram[1856] = 254;
    exp_62_ram[1857] = 255;
    exp_62_ram[1858] = 254;
    exp_62_ram[1859] = 250;
    exp_62_ram[1860] = 254;
    exp_62_ram[1861] = 0;
    exp_62_ram[1862] = 4;
    exp_62_ram[1863] = 2;
    exp_62_ram[1864] = 253;
    exp_62_ram[1865] = 0;
    exp_62_ram[1866] = 252;
    exp_62_ram[1867] = 250;
    exp_62_ram[1868] = 250;
    exp_62_ram[1869] = 0;
    exp_62_ram[1870] = 250;
    exp_62_ram[1871] = 2;
    exp_62_ram[1872] = 0;
    exp_62_ram[1873] = 252;
    exp_62_ram[1874] = 0;
    exp_62_ram[1875] = 252;
    exp_62_ram[1876] = 254;
    exp_62_ram[1877] = 252;
    exp_62_ram[1878] = 250;
    exp_62_ram[1879] = 0;
    exp_62_ram[1880] = 250;
    exp_62_ram[1881] = 13;
    exp_62_ram[1882] = 0;
    exp_62_ram[1883] = 254;
    exp_62_ram[1884] = 254;
    exp_62_ram[1885] = 2;
    exp_62_ram[1886] = 254;
    exp_62_ram[1887] = 249;
    exp_62_ram[1888] = 0;
    exp_62_ram[1889] = 248;
    exp_62_ram[1890] = 0;
    exp_62_ram[1891] = 0;
    exp_62_ram[1892] = 254;
    exp_62_ram[1893] = 0;
    exp_62_ram[1894] = 254;
    exp_62_ram[1895] = 0;
    exp_62_ram[1896] = 254;
    exp_62_ram[1897] = 1;
    exp_62_ram[1898] = 0;
    exp_62_ram[1899] = 250;
    exp_62_ram[1900] = 253;
    exp_62_ram[1901] = 250;
    exp_62_ram[1902] = 250;
    exp_62_ram[1903] = 207;
    exp_62_ram[1904] = 252;
    exp_62_ram[1905] = 250;
    exp_62_ram[1906] = 0;
    exp_62_ram[1907] = 250;
    exp_62_ram[1908] = 7;
    exp_62_ram[1909] = 253;
    exp_62_ram[1910] = 0;
    exp_62_ram[1911] = 252;
    exp_62_ram[1912] = 250;
    exp_62_ram[1913] = 250;
    exp_62_ram[1914] = 0;
    exp_62_ram[1915] = 250;
    exp_62_ram[1916] = 2;
    exp_62_ram[1917] = 0;
    exp_62_ram[1918] = 250;
    exp_62_ram[1919] = 0;
    exp_62_ram[1920] = 250;
    exp_62_ram[1921] = 3;
    exp_62_ram[1922] = 250;
    exp_62_ram[1923] = 0;
    exp_62_ram[1924] = 253;
    exp_62_ram[1925] = 0;
    exp_62_ram[1926] = 252;
    exp_62_ram[1927] = 250;
    exp_62_ram[1928] = 250;
    exp_62_ram[1929] = 0;
    exp_62_ram[1930] = 250;
    exp_62_ram[1931] = 0;
    exp_62_ram[1932] = 250;
    exp_62_ram[1933] = 0;
    exp_62_ram[1934] = 250;
    exp_62_ram[1935] = 0;
    exp_62_ram[1936] = 250;
    exp_62_ram[1937] = 0;
    exp_62_ram[1938] = 222;
    exp_62_ram[1939] = 253;
    exp_62_ram[1940] = 250;
    exp_62_ram[1941] = 0;
    exp_62_ram[1942] = 250;
    exp_62_ram[1943] = 255;
    exp_62_ram[1944] = 0;
    exp_62_ram[1945] = 253;
    exp_62_ram[1946] = 250;
    exp_62_ram[1947] = 250;
    exp_62_ram[1948] = 0;
    exp_62_ram[1949] = 250;
    exp_62_ram[1950] = 0;
    exp_62_ram[1951] = 0;
    exp_62_ram[1952] = 253;
    exp_62_ram[1953] = 0;
    exp_62_ram[1954] = 7;
    exp_62_ram[1955] = 7;
    exp_62_ram[1956] = 8;
    exp_62_ram[1957] = 0;
    exp_62_ram[1958] = 251;
    exp_62_ram[1959] = 2;
    exp_62_ram[1960] = 2;
    exp_62_ram[1961] = 3;
    exp_62_ram[1962] = 252;
    exp_62_ram[1963] = 0;
    exp_62_ram[1964] = 0;
    exp_62_ram[1965] = 0;
    exp_62_ram[1966] = 0;
    exp_62_ram[1967] = 0;
    exp_62_ram[1968] = 1;
    exp_62_ram[1969] = 1;
    exp_62_ram[1970] = 2;
    exp_62_ram[1971] = 252;
    exp_62_ram[1972] = 253;
    exp_62_ram[1973] = 254;
    exp_62_ram[1974] = 254;
    exp_62_ram[1975] = 254;
    exp_62_ram[1976] = 254;
    exp_62_ram[1977] = 253;
    exp_62_ram[1978] = 255;
    exp_62_ram[1979] = 0;
    exp_62_ram[1980] = 0;
    exp_62_ram[1981] = 206;
    exp_62_ram[1982] = 208;
    exp_62_ram[1983] = 254;
    exp_62_ram[1984] = 254;
    exp_62_ram[1985] = 0;
    exp_62_ram[1986] = 2;
    exp_62_ram[1987] = 2;
    exp_62_ram[1988] = 5;
    exp_62_ram[1989] = 0;
    exp_62_ram[1990] = 254;
    exp_62_ram[1991] = 0;
    exp_62_ram[1992] = 0;
    exp_62_ram[1993] = 2;
    exp_62_ram[1994] = 0;
    exp_62_ram[1995] = 254;
    exp_62_ram[1996] = 254;
    exp_62_ram[1997] = 0;
    exp_62_ram[1998] = 9;
    exp_62_ram[1999] = 0;
    exp_62_ram[2000] = 0;
    exp_62_ram[2001] = 195;
    exp_62_ram[2002] = 0;
    exp_62_ram[2003] = 1;
    exp_62_ram[2004] = 1;
    exp_62_ram[2005] = 2;
    exp_62_ram[2006] = 0;
    exp_62_ram[2007] = 246;
    exp_62_ram[2008] = 8;
    exp_62_ram[2009] = 8;
    exp_62_ram[2010] = 8;
    exp_62_ram[2011] = 10;
    exp_62_ram[2012] = 0;
    exp_62_ram[2013] = 1;
    exp_62_ram[2014] = 252;
    exp_62_ram[2015] = 0;
    exp_62_ram[2016] = 252;
    exp_62_ram[2017] = 1;
    exp_62_ram[2018] = 252;
    exp_62_ram[2019] = 0;
    exp_62_ram[2020] = 250;
    exp_62_ram[2021] = 250;
    exp_62_ram[2022] = 250;
    exp_62_ram[2023] = 252;
    exp_62_ram[2024] = 251;
    exp_62_ram[2025] = 251;
    exp_62_ram[2026] = 251;
    exp_62_ram[2027] = 252;
    exp_62_ram[2028] = 252;
    exp_62_ram[2029] = 252;
    exp_62_ram[2030] = 252;
    exp_62_ram[2031] = 253;
    exp_62_ram[2032] = 253;
    exp_62_ram[2033] = 246;
    exp_62_ram[2034] = 247;
    exp_62_ram[2035] = 247;
    exp_62_ram[2036] = 246;
    exp_62_ram[2037] = 246;
    exp_62_ram[2038] = 246;
    exp_62_ram[2039] = 246;
    exp_62_ram[2040] = 246;
    exp_62_ram[2041] = 248;
    exp_62_ram[2042] = 246;
    exp_62_ram[2043] = 0;
    exp_62_ram[2044] = 82;
    exp_62_ram[2045] = 254;
    exp_62_ram[2046] = 254;
    exp_62_ram[2047] = 251;
    exp_62_ram[2048] = 254;
    exp_62_ram[2049] = 254;
    exp_62_ram[2050] = 0;
    exp_62_ram[2051] = 14;
    exp_62_ram[2052] = 252;
    exp_62_ram[2053] = 252;
    exp_62_ram[2054] = 64;
    exp_62_ram[2055] = 252;
    exp_62_ram[2056] = 251;
    exp_62_ram[2057] = 251;
    exp_62_ram[2058] = 251;
    exp_62_ram[2059] = 252;
    exp_62_ram[2060] = 252;
    exp_62_ram[2061] = 252;
    exp_62_ram[2062] = 252;
    exp_62_ram[2063] = 253;
    exp_62_ram[2064] = 253;
    exp_62_ram[2065] = 246;
    exp_62_ram[2066] = 247;
    exp_62_ram[2067] = 247;
    exp_62_ram[2068] = 246;
    exp_62_ram[2069] = 246;
    exp_62_ram[2070] = 246;
    exp_62_ram[2071] = 246;
    exp_62_ram[2072] = 246;
    exp_62_ram[2073] = 248;
    exp_62_ram[2074] = 246;
    exp_62_ram[2075] = 0;
    exp_62_ram[2076] = 74;
    exp_62_ram[2077] = 254;
    exp_62_ram[2078] = 254;
    exp_62_ram[2079] = 1;
    exp_62_ram[2080] = 250;
    exp_62_ram[2081] = 0;
    exp_62_ram[2082] = 250;
    exp_62_ram[2083] = 1;
    exp_62_ram[2084] = 248;
    exp_62_ram[2085] = 0;
    exp_62_ram[2086] = 248;
    exp_62_ram[2087] = 248;
    exp_62_ram[2088] = 248;
    exp_62_ram[2089] = 252;
    exp_62_ram[2090] = 249;
    exp_62_ram[2091] = 249;
    exp_62_ram[2092] = 249;
    exp_62_ram[2093] = 249;
    exp_62_ram[2094] = 250;
    exp_62_ram[2095] = 250;
    exp_62_ram[2096] = 250;
    exp_62_ram[2097] = 250;
    exp_62_ram[2098] = 251;
    exp_62_ram[2099] = 246;
    exp_62_ram[2100] = 247;
    exp_62_ram[2101] = 247;
    exp_62_ram[2102] = 246;
    exp_62_ram[2103] = 246;
    exp_62_ram[2104] = 246;
    exp_62_ram[2105] = 246;
    exp_62_ram[2106] = 246;
    exp_62_ram[2107] = 248;
    exp_62_ram[2108] = 246;
    exp_62_ram[2109] = 0;
    exp_62_ram[2110] = 65;
    exp_62_ram[2111] = 254;
    exp_62_ram[2112] = 254;
    exp_62_ram[2113] = 249;
    exp_62_ram[2114] = 254;
    exp_62_ram[2115] = 254;
    exp_62_ram[2116] = 0;
    exp_62_ram[2117] = 125;
    exp_62_ram[2118] = 249;
    exp_62_ram[2119] = 250;
    exp_62_ram[2120] = 64;
    exp_62_ram[2121] = 248;
    exp_62_ram[2122] = 249;
    exp_62_ram[2123] = 249;
    exp_62_ram[2124] = 249;
    exp_62_ram[2125] = 249;
    exp_62_ram[2126] = 250;
    exp_62_ram[2127] = 250;
    exp_62_ram[2128] = 250;
    exp_62_ram[2129] = 250;
    exp_62_ram[2130] = 251;
    exp_62_ram[2131] = 246;
    exp_62_ram[2132] = 247;
    exp_62_ram[2133] = 247;
    exp_62_ram[2134] = 246;
    exp_62_ram[2135] = 246;
    exp_62_ram[2136] = 246;
    exp_62_ram[2137] = 246;
    exp_62_ram[2138] = 246;
    exp_62_ram[2139] = 248;
    exp_62_ram[2140] = 246;
    exp_62_ram[2141] = 0;
    exp_62_ram[2142] = 57;
    exp_62_ram[2143] = 254;
    exp_62_ram[2144] = 254;
    exp_62_ram[2145] = 0;
    exp_62_ram[2146] = 0;
    exp_62_ram[2147] = 0;
    exp_62_ram[2148] = 0;
    exp_62_ram[2149] = 1;
    exp_62_ram[2150] = 1;
    exp_62_ram[2151] = 1;
    exp_62_ram[2152] = 1;
    exp_62_ram[2153] = 2;
    exp_62_ram[2154] = 246;
    exp_62_ram[2155] = 247;
    exp_62_ram[2156] = 247;
    exp_62_ram[2157] = 246;
    exp_62_ram[2158] = 246;
    exp_62_ram[2159] = 246;
    exp_62_ram[2160] = 246;
    exp_62_ram[2161] = 246;
    exp_62_ram[2162] = 248;
    exp_62_ram[2163] = 246;
    exp_62_ram[2164] = 0;
    exp_62_ram[2165] = 52;
    exp_62_ram[2166] = 252;
    exp_62_ram[2167] = 252;
    exp_62_ram[2168] = 254;
    exp_62_ram[2169] = 253;
    exp_62_ram[2170] = 4;
    exp_62_ram[2171] = 254;
    exp_62_ram[2172] = 253;
    exp_62_ram[2173] = 0;
    exp_62_ram[2174] = 254;
    exp_62_ram[2175] = 253;
    exp_62_ram[2176] = 2;
    exp_62_ram[2177] = 254;
    exp_62_ram[2178] = 253;
    exp_62_ram[2179] = 0;
    exp_62_ram[2180] = 254;
    exp_62_ram[2181] = 253;
    exp_62_ram[2182] = 0;
    exp_62_ram[2183] = 254;
    exp_62_ram[2184] = 253;
    exp_62_ram[2185] = 0;
    exp_62_ram[2186] = 0;
    exp_62_ram[2187] = 0;
    exp_62_ram[2188] = 0;
    exp_62_ram[2189] = 0;
    exp_62_ram[2190] = 9;
    exp_62_ram[2191] = 9;
    exp_62_ram[2192] = 9;
    exp_62_ram[2193] = 10;
    exp_62_ram[2194] = 0;
    exp_62_ram[2195] = 248;
    exp_62_ram[2196] = 6;
    exp_62_ram[2197] = 6;
    exp_62_ram[2198] = 8;
    exp_62_ram[2199] = 250;
    exp_62_ram[2200] = 250;
    exp_62_ram[2201] = 252;
    exp_62_ram[2202] = 251;
    exp_62_ram[2203] = 251;
    exp_62_ram[2204] = 0;
    exp_62_ram[2205] = 103;
    exp_62_ram[2206] = 252;
    exp_62_ram[2207] = 253;
    exp_62_ram[2208] = 253;
    exp_62_ram[2209] = 253;
    exp_62_ram[2210] = 253;
    exp_62_ram[2211] = 254;
    exp_62_ram[2212] = 254;
    exp_62_ram[2213] = 254;
    exp_62_ram[2214] = 254;
    exp_62_ram[2215] = 248;
    exp_62_ram[2216] = 249;
    exp_62_ram[2217] = 249;
    exp_62_ram[2218] = 248;
    exp_62_ram[2219] = 248;
    exp_62_ram[2220] = 248;
    exp_62_ram[2221] = 248;
    exp_62_ram[2222] = 248;
    exp_62_ram[2223] = 250;
    exp_62_ram[2224] = 248;
    exp_62_ram[2225] = 0;
    exp_62_ram[2226] = 201;
    exp_62_ram[2227] = 0;
    exp_62_ram[2228] = 0;
    exp_62_ram[2229] = 7;
    exp_62_ram[2230] = 7;
    exp_62_ram[2231] = 8;
    exp_62_ram[2232] = 0;
    exp_62_ram[2233] = 254;
    exp_62_ram[2234] = 0;
    exp_62_ram[2235] = 2;
    exp_62_ram[2236] = 128;
    exp_62_ram[2237] = 254;
    exp_62_ram[2238] = 128;
    exp_62_ram[2239] = 0;
    exp_62_ram[2240] = 254;
    exp_62_ram[2241] = 254;
    exp_62_ram[2242] = 0;
    exp_62_ram[2243] = 254;
    exp_62_ram[2244] = 254;
    exp_62_ram[2245] = 254;
    exp_62_ram[2246] = 0;
    exp_62_ram[2247] = 254;
    exp_62_ram[2248] = 254;
    exp_62_ram[2249] = 254;
    exp_62_ram[2250] = 0;
    exp_62_ram[2251] = 0;
    exp_62_ram[2252] = 0;
    exp_62_ram[2253] = 254;
    exp_62_ram[2254] = 0;
    exp_62_ram[2255] = 254;
    exp_62_ram[2256] = 254;
    exp_62_ram[2257] = 0;
    exp_62_ram[2258] = 254;
    exp_62_ram[2259] = 254;
    exp_62_ram[2260] = 254;
    exp_62_ram[2261] = 0;
    exp_62_ram[2262] = 0;
    exp_62_ram[2263] = 1;
    exp_62_ram[2264] = 2;
    exp_62_ram[2265] = 0;
    exp_62_ram[2266] = 254;
    exp_62_ram[2267] = 0;
    exp_62_ram[2268] = 0;
    exp_62_ram[2269] = 2;
    exp_62_ram[2270] = 254;
    exp_62_ram[2271] = 254;
    exp_62_ram[2272] = 254;
    exp_62_ram[2273] = 254;
    exp_62_ram[2274] = 254;
    exp_62_ram[2275] = 254;
    exp_62_ram[2276] = 254;
    exp_62_ram[2277] = 254;
    exp_62_ram[2278] = 64;
    exp_62_ram[2279] = 0;
    exp_62_ram[2280] = 1;
    exp_62_ram[2281] = 64;
    exp_62_ram[2282] = 65;
    exp_62_ram[2283] = 0;
    exp_62_ram[2284] = 0;
    exp_62_ram[2285] = 0;
    exp_62_ram[2286] = 0;
    exp_62_ram[2287] = 0;
    exp_62_ram[2288] = 166;
    exp_62_ram[2289] = 0;
    exp_62_ram[2290] = 0;
    exp_62_ram[2291] = 0;
    exp_62_ram[2292] = 0;
    exp_62_ram[2293] = 1;
    exp_62_ram[2294] = 1;
    exp_62_ram[2295] = 2;
    exp_62_ram[2296] = 0;
    exp_62_ram[2297] = 254;
    exp_62_ram[2298] = 0;
    exp_62_ram[2299] = 2;
    exp_62_ram[2300] = 254;
    exp_62_ram[2301] = 254;
    exp_62_ram[2302] = 0;
    exp_62_ram[2303] = 2;
    exp_62_ram[2304] = 254;
    exp_62_ram[2305] = 6;
    exp_62_ram[2306] = 2;
    exp_62_ram[2307] = 0;
    exp_62_ram[2308] = 254;
    exp_62_ram[2309] = 25;
    exp_62_ram[2310] = 2;
    exp_62_ram[2311] = 0;
    exp_62_ram[2312] = 0;
    exp_62_ram[2313] = 0;
    exp_62_ram[2314] = 0;
    exp_62_ram[2315] = 0;
    exp_62_ram[2316] = 1;
    exp_62_ram[2317] = 2;
    exp_62_ram[2318] = 0;
    exp_62_ram[2319] = 254;
    exp_62_ram[2320] = 0;
    exp_62_ram[2321] = 0;
    exp_62_ram[2322] = 2;
    exp_62_ram[2323] = 254;
    exp_62_ram[2324] = 254;
    exp_62_ram[2325] = 249;
    exp_62_ram[2326] = 0;
    exp_62_ram[2327] = 0;
    exp_62_ram[2328] = 22;
    exp_62_ram[2329] = 0;
    exp_62_ram[2330] = 22;
    exp_62_ram[2331] = 0;
    exp_62_ram[2332] = 1;
    exp_62_ram[2333] = 1;
    exp_62_ram[2334] = 2;
    exp_62_ram[2335] = 0;
    exp_62_ram[2336] = 254;
    exp_62_ram[2337] = 0;
    exp_62_ram[2338] = 0;
    exp_62_ram[2339] = 2;
    exp_62_ram[2340] = 254;
    exp_62_ram[2341] = 254;
    exp_62_ram[2342] = 254;
    exp_62_ram[2343] = 0;
    exp_62_ram[2344] = 2;
    exp_62_ram[2345] = 254;
    exp_62_ram[2346] = 0;
    exp_62_ram[2347] = 0;
    exp_62_ram[2348] = 254;
    exp_62_ram[2349] = 0;
    exp_62_ram[2350] = 0;
    exp_62_ram[2351] = 254;
    exp_62_ram[2352] = 0;
    exp_62_ram[2353] = 0;
    exp_62_ram[2354] = 1;
    exp_62_ram[2355] = 3;
    exp_62_ram[2356] = 254;
    exp_62_ram[2357] = 0;
    exp_62_ram[2358] = 2;
    exp_62_ram[2359] = 254;
    exp_62_ram[2360] = 240;
    exp_62_ram[2361] = 0;
    exp_62_ram[2362] = 0;
    exp_62_ram[2363] = 1;
    exp_62_ram[2364] = 1;
    exp_62_ram[2365] = 1;
    exp_62_ram[2366] = 0;
    exp_62_ram[2367] = 1;
    exp_62_ram[2368] = 0;
    exp_62_ram[2369] = 1;
    exp_62_ram[2370] = 1;
    exp_62_ram[2371] = 2;
    exp_62_ram[2372] = 0;
    exp_62_ram[2373] = 249;
    exp_62_ram[2374] = 6;
    exp_62_ram[2375] = 6;
    exp_62_ram[2376] = 6;
    exp_62_ram[2377] = 7;
    exp_62_ram[2378] = 5;
    exp_62_ram[2379] = 5;
    exp_62_ram[2380] = 5;
    exp_62_ram[2381] = 5;
    exp_62_ram[2382] = 5;
    exp_62_ram[2383] = 5;
    exp_62_ram[2384] = 5;
    exp_62_ram[2385] = 5;
    exp_62_ram[2386] = 3;
    exp_62_ram[2387] = 7;
    exp_62_ram[2388] = 0;
    exp_62_ram[2389] = 0;
    exp_62_ram[2390] = 0;
    exp_62_ram[2391] = 250;
    exp_62_ram[2392] = 251;
    exp_62_ram[2393] = 123;
    exp_62_ram[2394] = 250;
    exp_62_ram[2395] = 1;
    exp_62_ram[2396] = 250;
    exp_62_ram[2397] = 250;
    exp_62_ram[2398] = 118;
    exp_62_ram[2399] = 251;
    exp_62_ram[2400] = 6;
    exp_62_ram[2401] = 251;
    exp_62_ram[2402] = 235;
    exp_62_ram[2403] = 0;
    exp_62_ram[2404] = 0;
    exp_62_ram[2405] = 24;
    exp_62_ram[2406] = 2;
    exp_62_ram[2407] = 248;
    exp_62_ram[2408] = 248;
    exp_62_ram[2409] = 251;
    exp_62_ram[2410] = 251;
    exp_62_ram[2411] = 249;
    exp_62_ram[2412] = 249;
    exp_62_ram[2413] = 0;
    exp_62_ram[2414] = 0;
    exp_62_ram[2415] = 0;
    exp_62_ram[2416] = 0;
    exp_62_ram[2417] = 0;
    exp_62_ram[2418] = 0;
    exp_62_ram[2419] = 0;
    exp_62_ram[2420] = 0;
    exp_62_ram[2421] = 250;
    exp_62_ram[2422] = 250;
    exp_62_ram[2423] = 251;
    exp_62_ram[2424] = 0;
    exp_62_ram[2425] = 250;
    exp_62_ram[2426] = 248;
    exp_62_ram[2427] = 0;
    exp_62_ram[2428] = 250;
    exp_62_ram[2429] = 1;
    exp_62_ram[2430] = 0;
    exp_62_ram[2431] = 251;
    exp_62_ram[2432] = 6;
    exp_62_ram[2433] = 251;
    exp_62_ram[2434] = 251;
    exp_62_ram[2435] = 231;
    exp_62_ram[2436] = 0;
    exp_62_ram[2437] = 0;
    exp_62_ram[2438] = 24;
    exp_62_ram[2439] = 2;
    exp_62_ram[2440] = 0;
    exp_62_ram[2441] = 0;
    exp_62_ram[2442] = 251;
    exp_62_ram[2443] = 251;
    exp_62_ram[2444] = 1;
    exp_62_ram[2445] = 0;
    exp_62_ram[2446] = 0;
    exp_62_ram[2447] = 1;
    exp_62_ram[2448] = 0;
    exp_62_ram[2449] = 0;
    exp_62_ram[2450] = 250;
    exp_62_ram[2451] = 250;
    exp_62_ram[2452] = 251;
    exp_62_ram[2453] = 0;
    exp_62_ram[2454] = 250;
    exp_62_ram[2455] = 249;
    exp_62_ram[2456] = 0;
    exp_62_ram[2457] = 0;
    exp_62_ram[2458] = 255;
    exp_62_ram[2459] = 0;
    exp_62_ram[2460] = 24;
    exp_62_ram[2461] = 2;
    exp_62_ram[2462] = 0;
    exp_62_ram[2463] = 65;
    exp_62_ram[2464] = 0;
    exp_62_ram[2465] = 251;
    exp_62_ram[2466] = 251;
    exp_62_ram[2467] = 1;
    exp_62_ram[2468] = 0;
    exp_62_ram[2469] = 0;
    exp_62_ram[2470] = 1;
    exp_62_ram[2471] = 0;
    exp_62_ram[2472] = 0;
    exp_62_ram[2473] = 250;
    exp_62_ram[2474] = 250;
    exp_62_ram[2475] = 0;
    exp_62_ram[2476] = 0;
    exp_62_ram[2477] = 225;
    exp_62_ram[2478] = 2;
    exp_62_ram[2479] = 0;
    exp_62_ram[2480] = 65;
    exp_62_ram[2481] = 0;
    exp_62_ram[2482] = 251;
    exp_62_ram[2483] = 251;
    exp_62_ram[2484] = 1;
    exp_62_ram[2485] = 0;
    exp_62_ram[2486] = 0;
    exp_62_ram[2487] = 1;
    exp_62_ram[2488] = 0;
    exp_62_ram[2489] = 0;
    exp_62_ram[2490] = 250;
    exp_62_ram[2491] = 250;
    exp_62_ram[2492] = 0;
    exp_62_ram[2493] = 0;
    exp_62_ram[2494] = 0;
    exp_62_ram[2495] = 64;
    exp_62_ram[2496] = 0;
    exp_62_ram[2497] = 0;
    exp_62_ram[2498] = 65;
    exp_62_ram[2499] = 0;
    exp_62_ram[2500] = 251;
    exp_62_ram[2501] = 251;
    exp_62_ram[2502] = 1;
    exp_62_ram[2503] = 0;
    exp_62_ram[2504] = 0;
    exp_62_ram[2505] = 1;
    exp_62_ram[2506] = 0;
    exp_62_ram[2507] = 0;
    exp_62_ram[2508] = 250;
    exp_62_ram[2509] = 250;
    exp_62_ram[2510] = 0;
    exp_62_ram[2511] = 0;
    exp_62_ram[2512] = 65;
    exp_62_ram[2513] = 0;
    exp_62_ram[2514] = 251;
    exp_62_ram[2515] = 251;
    exp_62_ram[2516] = 1;
    exp_62_ram[2517] = 0;
    exp_62_ram[2518] = 0;
    exp_62_ram[2519] = 1;
    exp_62_ram[2520] = 0;
    exp_62_ram[2521] = 0;
    exp_62_ram[2522] = 250;
    exp_62_ram[2523] = 250;
    exp_62_ram[2524] = 251;
    exp_62_ram[2525] = 251;
    exp_62_ram[2526] = 0;
    exp_62_ram[2527] = 0;
    exp_62_ram[2528] = 6;
    exp_62_ram[2529] = 6;
    exp_62_ram[2530] = 6;
    exp_62_ram[2531] = 6;
    exp_62_ram[2532] = 5;
    exp_62_ram[2533] = 5;
    exp_62_ram[2534] = 5;
    exp_62_ram[2535] = 5;
    exp_62_ram[2536] = 4;
    exp_62_ram[2537] = 4;
    exp_62_ram[2538] = 4;
    exp_62_ram[2539] = 4;
    exp_62_ram[2540] = 3;
    exp_62_ram[2541] = 7;
    exp_62_ram[2542] = 0;
    exp_62_ram[2543] = 246;
    exp_62_ram[2544] = 8;
    exp_62_ram[2545] = 8;
    exp_62_ram[2546] = 8;
    exp_62_ram[2547] = 9;
    exp_62_ram[2548] = 9;
    exp_62_ram[2549] = 10;
    exp_62_ram[2550] = 248;
    exp_62_ram[2551] = 249;
    exp_62_ram[2552] = 0;
    exp_62_ram[2553] = 0;
    exp_62_ram[2554] = 0;
    exp_62_ram[2555] = 0;
    exp_62_ram[2556] = 1;
    exp_62_ram[2557] = 1;
    exp_62_ram[2558] = 1;
    exp_62_ram[2559] = 1;
    exp_62_ram[2560] = 2;
    exp_62_ram[2561] = 250;
    exp_62_ram[2562] = 251;
    exp_62_ram[2563] = 251;
    exp_62_ram[2564] = 250;
    exp_62_ram[2565] = 250;
    exp_62_ram[2566] = 252;
    exp_62_ram[2567] = 252;
    exp_62_ram[2568] = 252;
    exp_62_ram[2569] = 252;
    exp_62_ram[2570] = 250;
    exp_62_ram[2571] = 251;
    exp_62_ram[2572] = 251;
    exp_62_ram[2573] = 251;
    exp_62_ram[2574] = 251;
    exp_62_ram[2575] = 252;
    exp_62_ram[2576] = 252;
    exp_62_ram[2577] = 252;
    exp_62_ram[2578] = 252;
    exp_62_ram[2579] = 246;
    exp_62_ram[2580] = 247;
    exp_62_ram[2581] = 247;
    exp_62_ram[2582] = 246;
    exp_62_ram[2583] = 246;
    exp_62_ram[2584] = 246;
    exp_62_ram[2585] = 246;
    exp_62_ram[2586] = 246;
    exp_62_ram[2587] = 248;
    exp_62_ram[2588] = 246;
    exp_62_ram[2589] = 0;
    exp_62_ram[2590] = 201;
    exp_62_ram[2591] = 252;
    exp_62_ram[2592] = 252;
    exp_62_ram[2593] = 252;
    exp_62_ram[2594] = 2;
    exp_62_ram[2595] = 253;
    exp_62_ram[2596] = 253;
    exp_62_ram[2597] = 255;
    exp_62_ram[2598] = 31;
    exp_62_ram[2599] = 255;
    exp_62_ram[2600] = 0;
    exp_62_ram[2601] = 0;
    exp_62_ram[2602] = 0;
    exp_62_ram[2603] = 0;
    exp_62_ram[2604] = 0;
    exp_62_ram[2605] = 0;
    exp_62_ram[2606] = 252;
    exp_62_ram[2607] = 252;
    exp_62_ram[2608] = 11;
    exp_62_ram[2609] = 252;
    exp_62_ram[2610] = 10;
    exp_62_ram[2611] = 250;
    exp_62_ram[2612] = 251;
    exp_62_ram[2613] = 251;
    exp_62_ram[2614] = 251;
    exp_62_ram[2615] = 251;
    exp_62_ram[2616] = 252;
    exp_62_ram[2617] = 252;
    exp_62_ram[2618] = 252;
    exp_62_ram[2619] = 252;
    exp_62_ram[2620] = 246;
    exp_62_ram[2621] = 247;
    exp_62_ram[2622] = 247;
    exp_62_ram[2623] = 246;
    exp_62_ram[2624] = 246;
    exp_62_ram[2625] = 246;
    exp_62_ram[2626] = 246;
    exp_62_ram[2627] = 246;
    exp_62_ram[2628] = 248;
    exp_62_ram[2629] = 246;
    exp_62_ram[2630] = 0;
    exp_62_ram[2631] = 228;
    exp_62_ram[2632] = 0;
    exp_62_ram[2633] = 0;
    exp_62_ram[2634] = 0;
    exp_62_ram[2635] = 225;
    exp_62_ram[2636] = 0;
    exp_62_ram[2637] = 0;
    exp_62_ram[2638] = 0;
    exp_62_ram[2639] = 0;
    exp_62_ram[2640] = 253;
    exp_62_ram[2641] = 253;
    exp_62_ram[2642] = 64;
    exp_62_ram[2643] = 0;
    exp_62_ram[2644] = 1;
    exp_62_ram[2645] = 64;
    exp_62_ram[2646] = 65;
    exp_62_ram[2647] = 0;
    exp_62_ram[2648] = 252;
    exp_62_ram[2649] = 252;
    exp_62_ram[2650] = 1;
    exp_62_ram[2651] = 253;
    exp_62_ram[2652] = 253;
    exp_62_ram[2653] = 252;
    exp_62_ram[2654] = 252;
    exp_62_ram[2655] = 0;
    exp_62_ram[2656] = 40;
    exp_62_ram[2657] = 0;
    exp_62_ram[2658] = 65;
    exp_62_ram[2659] = 0;
    exp_62_ram[2660] = 253;
    exp_62_ram[2661] = 253;
    exp_62_ram[2662] = 65;
    exp_62_ram[2663] = 0;
    exp_62_ram[2664] = 0;
    exp_62_ram[2665] = 65;
    exp_62_ram[2666] = 64;
    exp_62_ram[2667] = 0;
    exp_62_ram[2668] = 252;
    exp_62_ram[2669] = 252;
    exp_62_ram[2670] = 249;
    exp_62_ram[2671] = 246;
    exp_62_ram[2672] = 253;
    exp_62_ram[2673] = 253;
    exp_62_ram[2674] = 0;
    exp_62_ram[2675] = 114;
    exp_62_ram[2676] = 246;
    exp_62_ram[2677] = 246;
    exp_62_ram[2678] = 246;
    exp_62_ram[2679] = 246;
    exp_62_ram[2680] = 247;
    exp_62_ram[2681] = 247;
    exp_62_ram[2682] = 247;
    exp_62_ram[2683] = 247;
    exp_62_ram[2684] = 248;
    exp_62_ram[2685] = 0;
    exp_62_ram[2686] = 1;
    exp_62_ram[2687] = 1;
    exp_62_ram[2688] = 0;
    exp_62_ram[2689] = 0;
    exp_62_ram[2690] = 0;
    exp_62_ram[2691] = 0;
    exp_62_ram[2692] = 0;
    exp_62_ram[2693] = 2;
    exp_62_ram[2694] = 252;
    exp_62_ram[2695] = 0;
    exp_62_ram[2696] = 249;
    exp_62_ram[2697] = 0;
    exp_62_ram[2698] = 2;
    exp_62_ram[2699] = 7;
    exp_62_ram[2700] = 252;
    exp_62_ram[2701] = 6;
    exp_62_ram[2702] = 250;
    exp_62_ram[2703] = 251;
    exp_62_ram[2704] = 251;
    exp_62_ram[2705] = 251;
    exp_62_ram[2706] = 251;
    exp_62_ram[2707] = 252;
    exp_62_ram[2708] = 252;
    exp_62_ram[2709] = 252;
    exp_62_ram[2710] = 252;
    exp_62_ram[2711] = 246;
    exp_62_ram[2712] = 247;
    exp_62_ram[2713] = 247;
    exp_62_ram[2714] = 246;
    exp_62_ram[2715] = 246;
    exp_62_ram[2716] = 246;
    exp_62_ram[2717] = 246;
    exp_62_ram[2718] = 246;
    exp_62_ram[2719] = 248;
    exp_62_ram[2720] = 246;
    exp_62_ram[2721] = 0;
    exp_62_ram[2722] = 205;
    exp_62_ram[2723] = 0;
    exp_62_ram[2724] = 249;
    exp_62_ram[2725] = 2;
    exp_62_ram[2726] = 0;
    exp_62_ram[2727] = 249;
    exp_62_ram[2728] = 2;
    exp_62_ram[2729] = 253;
    exp_62_ram[2730] = 253;
    exp_62_ram[2731] = 0;
    exp_62_ram[2732] = 0;
    exp_62_ram[2733] = 9;
    exp_62_ram[2734] = 9;
    exp_62_ram[2735] = 9;
    exp_62_ram[2736] = 9;
    exp_62_ram[2737] = 8;
    exp_62_ram[2738] = 10;
    exp_62_ram[2739] = 0;
    exp_62_ram[2740] = 252;
    exp_62_ram[2741] = 2;
    exp_62_ram[2742] = 2;
    exp_62_ram[2743] = 3;
    exp_62_ram[2744] = 3;
    exp_62_ram[2745] = 3;
    exp_62_ram[2746] = 3;
    exp_62_ram[2747] = 3;
    exp_62_ram[2748] = 3;
    exp_62_ram[2749] = 4;
    exp_62_ram[2750] = 252;
    exp_62_ram[2751] = 254;
    exp_62_ram[2752] = 0;
    exp_62_ram[2753] = 0;
    exp_62_ram[2754] = 0;
    exp_62_ram[2755] = 9;
    exp_62_ram[2756] = 0;
    exp_62_ram[2757] = 0;
    exp_62_ram[2758] = 0;
    exp_62_ram[2759] = 0;
    exp_62_ram[2760] = 0;
    exp_62_ram[2761] = 0;
    exp_62_ram[2762] = 214;
    exp_62_ram[2763] = 0;
    exp_62_ram[2764] = 0;
    exp_62_ram[2765] = 252;
    exp_62_ram[2766] = 0;
    exp_62_ram[2767] = 40;
    exp_62_ram[2768] = 40;
    exp_62_ram[2769] = 253;
    exp_62_ram[2770] = 0;
    exp_62_ram[2771] = 252;
    exp_62_ram[2772] = 252;
    exp_62_ram[2773] = 0;
    exp_62_ram[2774] = 253;
    exp_62_ram[2775] = 0;
    exp_62_ram[2776] = 0;
    exp_62_ram[2777] = 252;
    exp_62_ram[2778] = 1;
    exp_62_ram[2779] = 1;
    exp_62_ram[2780] = 253;
    exp_62_ram[2781] = 0;
    exp_62_ram[2782] = 0;
    exp_62_ram[2783] = 0;
    exp_62_ram[2784] = 0;
    exp_62_ram[2785] = 0;
    exp_62_ram[2786] = 0;
    exp_62_ram[2787] = 3;
    exp_62_ram[2788] = 3;
    exp_62_ram[2789] = 3;
    exp_62_ram[2790] = 3;
    exp_62_ram[2791] = 2;
    exp_62_ram[2792] = 2;
    exp_62_ram[2793] = 2;
    exp_62_ram[2794] = 2;
    exp_62_ram[2795] = 4;
    exp_62_ram[2796] = 0;
    exp_62_ram[2797] = 253;
    exp_62_ram[2798] = 2;
    exp_62_ram[2799] = 2;
    exp_62_ram[2800] = 3;
    exp_62_ram[2801] = 3;
    exp_62_ram[2802] = 3;
    exp_62_ram[2803] = 252;
    exp_62_ram[2804] = 252;
    exp_62_ram[2805] = 241;
    exp_62_ram[2806] = 0;
    exp_62_ram[2807] = 0;
    exp_62_ram[2808] = 0;
    exp_62_ram[2809] = 9;
    exp_62_ram[2810] = 0;
    exp_62_ram[2811] = 0;
    exp_62_ram[2812] = 0;
    exp_62_ram[2813] = 0;
    exp_62_ram[2814] = 0;
    exp_62_ram[2815] = 0;
    exp_62_ram[2816] = 200;
    exp_62_ram[2817] = 0;
    exp_62_ram[2818] = 0;
    exp_62_ram[2819] = 254;
    exp_62_ram[2820] = 254;
    exp_62_ram[2821] = 253;
    exp_62_ram[2822] = 253;
    exp_62_ram[2823] = 254;
    exp_62_ram[2824] = 254;
    exp_62_ram[2825] = 64;
    exp_62_ram[2826] = 0;
    exp_62_ram[2827] = 1;
    exp_62_ram[2828] = 64;
    exp_62_ram[2829] = 65;
    exp_62_ram[2830] = 0;
    exp_62_ram[2831] = 0;
    exp_62_ram[2832] = 0;
    exp_62_ram[2833] = 0;
    exp_62_ram[2834] = 40;
    exp_62_ram[2835] = 40;
    exp_62_ram[2836] = 0;
    exp_62_ram[2837] = 2;
    exp_62_ram[2838] = 2;
    exp_62_ram[2839] = 2;
    exp_62_ram[2840] = 2;
    exp_62_ram[2841] = 3;
    exp_62_ram[2842] = 0;
    exp_62_ram[2843] = 249;
    exp_62_ram[2844] = 6;
    exp_62_ram[2845] = 6;
    exp_62_ram[2846] = 7;
    exp_62_ram[2847] = 248;
    exp_62_ram[2848] = 0;
    exp_62_ram[2849] = 138;
    exp_62_ram[2850] = 0;
    exp_62_ram[2851] = 0;
    exp_62_ram[2852] = 0;
    exp_62_ram[2853] = 0;
    exp_62_ram[2854] = 1;
    exp_62_ram[2855] = 252;
    exp_62_ram[2856] = 252;
    exp_62_ram[2857] = 252;
    exp_62_ram[2858] = 254;
    exp_62_ram[2859] = 254;
    exp_62_ram[2860] = 1;
    exp_62_ram[2861] = 254;
    exp_62_ram[2862] = 0;
    exp_62_ram[2863] = 140;
    exp_62_ram[2864] = 0;
    exp_62_ram[2865] = 0;
    exp_62_ram[2866] = 0;
    exp_62_ram[2867] = 0;
    exp_62_ram[2868] = 1;
    exp_62_ram[2869] = 1;
    exp_62_ram[2870] = 1;
    exp_62_ram[2871] = 1;
    exp_62_ram[2872] = 2;
    exp_62_ram[2873] = 251;
    exp_62_ram[2874] = 250;
    exp_62_ram[2875] = 251;
    exp_62_ram[2876] = 251;
    exp_62_ram[2877] = 250;
    exp_62_ram[2878] = 252;
    exp_62_ram[2879] = 252;
    exp_62_ram[2880] = 252;
    exp_62_ram[2881] = 252;
    exp_62_ram[2882] = 2;
    exp_62_ram[2883] = 252;
    exp_62_ram[2884] = 254;
    exp_62_ram[2885] = 4;
    exp_62_ram[2886] = 249;
    exp_62_ram[2887] = 1;
    exp_62_ram[2888] = 0;
    exp_62_ram[2889] = 0;
    exp_62_ram[2890] = 0;
    exp_62_ram[2891] = 254;
    exp_62_ram[2892] = 0;
    exp_62_ram[2893] = 255;
    exp_62_ram[2894] = 0;
    exp_62_ram[2895] = 254;
    exp_62_ram[2896] = 0;
    exp_62_ram[2897] = 41;
    exp_62_ram[2898] = 254;
    exp_62_ram[2899] = 0;
    exp_62_ram[2900] = 0;
    exp_62_ram[2901] = 254;
    exp_62_ram[2902] = 0;
    exp_62_ram[2903] = 254;
    exp_62_ram[2904] = 254;
    exp_62_ram[2905] = 0;
    exp_62_ram[2906] = 250;
    exp_62_ram[2907] = 0;
    exp_62_ram[2908] = 41;
    exp_62_ram[2909] = 2;
    exp_62_ram[2910] = 0;
    exp_62_ram[2911] = 254;
    exp_62_ram[2912] = 5;
    exp_62_ram[2913] = 249;
    exp_62_ram[2914] = 1;
    exp_62_ram[2915] = 0;
    exp_62_ram[2916] = 0;
    exp_62_ram[2917] = 0;
    exp_62_ram[2918] = 254;
    exp_62_ram[2919] = 0;
    exp_62_ram[2920] = 254;
    exp_62_ram[2921] = 0;
    exp_62_ram[2922] = 255;
    exp_62_ram[2923] = 0;
    exp_62_ram[2924] = 251;
    exp_62_ram[2925] = 0;
    exp_62_ram[2926] = 41;
    exp_62_ram[2927] = 0;
    exp_62_ram[2928] = 0;
    exp_62_ram[2929] = 254;
    exp_62_ram[2930] = 0;
    exp_62_ram[2931] = 254;
    exp_62_ram[2932] = 254;
    exp_62_ram[2933] = 0;
    exp_62_ram[2934] = 250;
    exp_62_ram[2935] = 0;
    exp_62_ram[2936] = 41;
    exp_62_ram[2937] = 2;
    exp_62_ram[2938] = 0;
    exp_62_ram[2939] = 249;
    exp_62_ram[2940] = 0;
    exp_62_ram[2941] = 0;
    exp_62_ram[2942] = 0;
    exp_62_ram[2943] = 37;
    exp_62_ram[2944] = 0;
    exp_62_ram[2945] = 0;
    exp_62_ram[2946] = 250;
    exp_62_ram[2947] = 250;
    exp_62_ram[2948] = 250;
    exp_62_ram[2949] = 15;
    exp_62_ram[2950] = 3;
    exp_62_ram[2951] = 15;
    exp_62_ram[2952] = 0;
    exp_62_ram[2953] = 41;
    exp_62_ram[2954] = 0;
    exp_62_ram[2955] = 250;
    exp_62_ram[2956] = 15;
    exp_62_ram[2957] = 3;
    exp_62_ram[2958] = 15;
    exp_62_ram[2959] = 0;
    exp_62_ram[2960] = 41;
    exp_62_ram[2961] = 0;
    exp_62_ram[2962] = 0;
    exp_62_ram[2963] = 41;
    exp_62_ram[2964] = 2;
    exp_62_ram[2965] = 0;
    exp_62_ram[2966] = 249;
    exp_62_ram[2967] = 0;
    exp_62_ram[2968] = 0;
    exp_62_ram[2969] = 0;
    exp_62_ram[2970] = 30;
    exp_62_ram[2971] = 0;
    exp_62_ram[2972] = 0;
    exp_62_ram[2973] = 250;
    exp_62_ram[2974] = 250;
    exp_62_ram[2975] = 250;
    exp_62_ram[2976] = 15;
    exp_62_ram[2977] = 3;
    exp_62_ram[2978] = 15;
    exp_62_ram[2979] = 0;
    exp_62_ram[2980] = 41;
    exp_62_ram[2981] = 0;
    exp_62_ram[2982] = 250;
    exp_62_ram[2983] = 15;
    exp_62_ram[2984] = 3;
    exp_62_ram[2985] = 15;
    exp_62_ram[2986] = 0;
    exp_62_ram[2987] = 41;
    exp_62_ram[2988] = 0;
    exp_62_ram[2989] = 0;
    exp_62_ram[2990] = 41;
    exp_62_ram[2991] = 3;
    exp_62_ram[2992] = 0;
    exp_62_ram[2993] = 249;
    exp_62_ram[2994] = 0;
    exp_62_ram[2995] = 0;
    exp_62_ram[2996] = 0;
    exp_62_ram[2997] = 24;
    exp_62_ram[2998] = 0;
    exp_62_ram[2999] = 0;
    exp_62_ram[3000] = 250;
    exp_62_ram[3001] = 250;
    exp_62_ram[3002] = 250;
    exp_62_ram[3003] = 15;
    exp_62_ram[3004] = 3;
    exp_62_ram[3005] = 15;
    exp_62_ram[3006] = 0;
    exp_62_ram[3007] = 41;
    exp_62_ram[3008] = 0;
    exp_62_ram[3009] = 250;
    exp_62_ram[3010] = 15;
    exp_62_ram[3011] = 3;
    exp_62_ram[3012] = 15;
    exp_62_ram[3013] = 0;
    exp_62_ram[3014] = 41;
    exp_62_ram[3015] = 0;
    exp_62_ram[3016] = 0;
    exp_62_ram[3017] = 41;
    exp_62_ram[3018] = 3;
    exp_62_ram[3019] = 0;
    exp_62_ram[3020] = 249;
    exp_62_ram[3021] = 0;
    exp_62_ram[3022] = 0;
    exp_62_ram[3023] = 0;
    exp_62_ram[3024] = 17;
    exp_62_ram[3025] = 0;
    exp_62_ram[3026] = 0;
    exp_62_ram[3027] = 250;
    exp_62_ram[3028] = 250;
    exp_62_ram[3029] = 250;
    exp_62_ram[3030] = 15;
    exp_62_ram[3031] = 3;
    exp_62_ram[3032] = 15;
    exp_62_ram[3033] = 0;
    exp_62_ram[3034] = 41;
    exp_62_ram[3035] = 0;
    exp_62_ram[3036] = 250;
    exp_62_ram[3037] = 15;
    exp_62_ram[3038] = 3;
    exp_62_ram[3039] = 15;
    exp_62_ram[3040] = 0;
    exp_62_ram[3041] = 41;
    exp_62_ram[3042] = 0;
    exp_62_ram[3043] = 0;
    exp_62_ram[3044] = 41;
    exp_62_ram[3045] = 2;
    exp_62_ram[3046] = 0;
    exp_62_ram[3047] = 249;
    exp_62_ram[3048] = 1;
    exp_62_ram[3049] = 118;
    exp_62_ram[3050] = 62;
    exp_62_ram[3051] = 0;
    exp_62_ram[3052] = 10;
    exp_62_ram[3053] = 0;
    exp_62_ram[3054] = 0;
    exp_62_ram[3055] = 250;
    exp_62_ram[3056] = 250;
    exp_62_ram[3057] = 250;
    exp_62_ram[3058] = 15;
    exp_62_ram[3059] = 3;
    exp_62_ram[3060] = 15;
    exp_62_ram[3061] = 0;
    exp_62_ram[3062] = 41;
    exp_62_ram[3063] = 0;
    exp_62_ram[3064] = 250;
    exp_62_ram[3065] = 6;
    exp_62_ram[3066] = 0;
    exp_62_ram[3067] = 6;
    exp_62_ram[3068] = 0;
    exp_62_ram[3069] = 0;
    exp_62_ram[3070] = 250;
    exp_62_ram[3071] = 250;
    exp_62_ram[3072] = 250;
    exp_62_ram[3073] = 15;
    exp_62_ram[3074] = 3;
    exp_62_ram[3075] = 15;
    exp_62_ram[3076] = 0;
    exp_62_ram[3077] = 41;
    exp_62_ram[3078] = 0;
    exp_62_ram[3079] = 250;
    exp_62_ram[3080] = 0;
    exp_62_ram[3081] = 0;
    exp_62_ram[3082] = 2;
    exp_62_ram[3083] = 0;
    exp_62_ram[3084] = 0;
    exp_62_ram[3085] = 250;
    exp_62_ram[3086] = 250;
    exp_62_ram[3087] = 250;
    exp_62_ram[3088] = 15;
    exp_62_ram[3089] = 3;
    exp_62_ram[3090] = 15;
    exp_62_ram[3091] = 0;
    exp_62_ram[3092] = 41;
    exp_62_ram[3093] = 0;
    exp_62_ram[3094] = 250;
    exp_62_ram[3095] = 15;
    exp_62_ram[3096] = 3;
    exp_62_ram[3097] = 15;
    exp_62_ram[3098] = 0;
    exp_62_ram[3099] = 41;
    exp_62_ram[3100] = 0;
    exp_62_ram[3101] = 0;
    exp_62_ram[3102] = 41;
    exp_62_ram[3103] = 0;
    exp_62_ram[3104] = 0;
    exp_62_ram[3105] = 0;
    exp_62_ram[3106] = 41;
    exp_62_ram[3107] = 0;
    exp_62_ram[3108] = 0;
    exp_62_ram[3109] = 41;
    exp_62_ram[3110] = 0;
    exp_62_ram[3111] = 6;
    exp_62_ram[3112] = 6;
    exp_62_ram[3113] = 7;
    exp_62_ram[3114] = 0;
    exp_62_ram[3115] = 254;
    exp_62_ram[3116] = 0;
    exp_62_ram[3117] = 0;
    exp_62_ram[3118] = 2;
    exp_62_ram[3119] = 254;
    exp_62_ram[3120] = 254;
    exp_62_ram[3121] = 55;
    exp_62_ram[3122] = 0;
    exp_62_ram[3123] = 0;
    exp_62_ram[3124] = 185;
    exp_62_ram[3125] = 0;
    exp_62_ram[3126] = 0;
    exp_62_ram[3127] = 1;
    exp_62_ram[3128] = 1;
    exp_62_ram[3129] = 2;
    exp_62_ram[3130] = 0;
    exp_62_ram[3131] = 248;
    exp_62_ram[3132] = 6;
    exp_62_ram[3133] = 6;
    exp_62_ram[3134] = 7;
    exp_62_ram[3135] = 7;
    exp_62_ram[3136] = 7;
    exp_62_ram[3137] = 7;
    exp_62_ram[3138] = 7;
    exp_62_ram[3139] = 7;
    exp_62_ram[3140] = 5;
    exp_62_ram[3141] = 5;
    exp_62_ram[3142] = 8;
    exp_62_ram[3143] = 248;
    exp_62_ram[3144] = 248;
    exp_62_ram[3145] = 248;
    exp_62_ram[3146] = 123;
    exp_62_ram[3147] = 250;
    exp_62_ram[3148] = 0;
    exp_62_ram[3149] = 250;
    exp_62_ram[3150] = 251;
    exp_62_ram[3151] = 0;
    exp_62_ram[3152] = 175;
    exp_62_ram[3153] = 252;
    exp_62_ram[3154] = 252;
    exp_62_ram[3155] = 0;
    exp_62_ram[3156] = 24;
    exp_62_ram[3157] = 2;
    exp_62_ram[3158] = 252;
    exp_62_ram[3159] = 252;
    exp_62_ram[3160] = 0;
    exp_62_ram[3161] = 0;
    exp_62_ram[3162] = 248;
    exp_62_ram[3163] = 0;
    exp_62_ram[3164] = 6;
    exp_62_ram[3165] = 248;
    exp_62_ram[3166] = 0;
    exp_62_ram[3167] = 0;
    exp_62_ram[3168] = 248;
    exp_62_ram[3169] = 0;
    exp_62_ram[3170] = 4;
    exp_62_ram[3171] = 251;
    exp_62_ram[3172] = 0;
    exp_62_ram[3173] = 250;
    exp_62_ram[3174] = 251;
    exp_62_ram[3175] = 0;
    exp_62_ram[3176] = 252;
    exp_62_ram[3177] = 0;
    exp_62_ram[3178] = 250;
    exp_62_ram[3179] = 252;
    exp_62_ram[3180] = 0;
    exp_62_ram[3181] = 0;
    exp_62_ram[3182] = 248;
    exp_62_ram[3183] = 248;
    exp_62_ram[3184] = 65;
    exp_62_ram[3185] = 0;
    exp_62_ram[3186] = 0;
    exp_62_ram[3187] = 65;
    exp_62_ram[3188] = 64;
    exp_62_ram[3189] = 0;
    exp_62_ram[3190] = 248;
    exp_62_ram[3191] = 248;
    exp_62_ram[3192] = 245;
    exp_62_ram[3193] = 0;
    exp_62_ram[3194] = 250;
    exp_62_ram[3195] = 252;
    exp_62_ram[3196] = 251;
    exp_62_ram[3197] = 0;
    exp_62_ram[3198] = 251;
    exp_62_ram[3199] = 0;
    exp_62_ram[3200] = 0;
    exp_62_ram[3201] = 167;
    exp_62_ram[3202] = 252;
    exp_62_ram[3203] = 252;
    exp_62_ram[3204] = 0;
    exp_62_ram[3205] = 24;
    exp_62_ram[3206] = 2;
    exp_62_ram[3207] = 252;
    exp_62_ram[3208] = 252;
    exp_62_ram[3209] = 0;
    exp_62_ram[3210] = 0;
    exp_62_ram[3211] = 248;
    exp_62_ram[3212] = 0;
    exp_62_ram[3213] = 8;
    exp_62_ram[3214] = 248;
    exp_62_ram[3215] = 0;
    exp_62_ram[3216] = 0;
    exp_62_ram[3217] = 248;
    exp_62_ram[3218] = 0;
    exp_62_ram[3219] = 6;
    exp_62_ram[3220] = 251;
    exp_62_ram[3221] = 0;
    exp_62_ram[3222] = 250;
    exp_62_ram[3223] = 251;
    exp_62_ram[3224] = 0;
    exp_62_ram[3225] = 252;
    exp_62_ram[3226] = 0;
    exp_62_ram[3227] = 250;
    exp_62_ram[3228] = 252;
    exp_62_ram[3229] = 0;
    exp_62_ram[3230] = 252;
    exp_62_ram[3231] = 0;
    exp_62_ram[3232] = 252;
    exp_62_ram[3233] = 252;
    exp_62_ram[3234] = 0;
    exp_62_ram[3235] = 0;
    exp_62_ram[3236] = 248;
    exp_62_ram[3237] = 248;
    exp_62_ram[3238] = 65;
    exp_62_ram[3239] = 0;
    exp_62_ram[3240] = 0;
    exp_62_ram[3241] = 65;
    exp_62_ram[3242] = 64;
    exp_62_ram[3243] = 0;
    exp_62_ram[3244] = 248;
    exp_62_ram[3245] = 248;
    exp_62_ram[3246] = 243;
    exp_62_ram[3247] = 0;
    exp_62_ram[3248] = 251;
    exp_62_ram[3249] = 137;
    exp_62_ram[3250] = 250;
    exp_62_ram[3251] = 248;
    exp_62_ram[3252] = 0;
    exp_62_ram[3253] = 24;
    exp_62_ram[3254] = 0;
    exp_62_ram[3255] = 87;
    exp_62_ram[3256] = 0;
    exp_62_ram[3257] = 0;
    exp_62_ram[3258] = 248;
    exp_62_ram[3259] = 250;
    exp_62_ram[3260] = 249;
    exp_62_ram[3261] = 0;
    exp_62_ram[3262] = 250;
    exp_62_ram[3263] = 251;
    exp_62_ram[3264] = 249;
    exp_62_ram[3265] = 0;
    exp_62_ram[3266] = 250;
    exp_62_ram[3267] = 251;
    exp_62_ram[3268] = 0;
    exp_62_ram[3269] = 2;
    exp_62_ram[3270] = 250;
    exp_62_ram[3271] = 252;
    exp_62_ram[3272] = 249;
    exp_62_ram[3273] = 0;
    exp_62_ram[3274] = 252;
    exp_62_ram[3275] = 250;
    exp_62_ram[3276] = 248;
    exp_62_ram[3277] = 65;
    exp_62_ram[3278] = 248;
    exp_62_ram[3279] = 248;
    exp_62_ram[3280] = 0;
    exp_62_ram[3281] = 225;
    exp_62_ram[3282] = 0;
    exp_62_ram[3283] = 80;
    exp_62_ram[3284] = 0;
    exp_62_ram[3285] = 0;
    exp_62_ram[3286] = 248;
    exp_62_ram[3287] = 250;
    exp_62_ram[3288] = 249;
    exp_62_ram[3289] = 250;
    exp_62_ram[3290] = 250;
    exp_62_ram[3291] = 248;
    exp_62_ram[3292] = 65;
    exp_62_ram[3293] = 248;
    exp_62_ram[3294] = 248;
    exp_62_ram[3295] = 3;
    exp_62_ram[3296] = 0;
    exp_62_ram[3297] = 77;
    exp_62_ram[3298] = 0;
    exp_62_ram[3299] = 0;
    exp_62_ram[3300] = 248;
    exp_62_ram[3301] = 250;
    exp_62_ram[3302] = 249;
    exp_62_ram[3303] = 250;
    exp_62_ram[3304] = 250;
    exp_62_ram[3305] = 248;
    exp_62_ram[3306] = 65;
    exp_62_ram[3307] = 248;
    exp_62_ram[3308] = 248;
    exp_62_ram[3309] = 250;
    exp_62_ram[3310] = 248;
    exp_62_ram[3311] = 250;
    exp_62_ram[3312] = 250;
    exp_62_ram[3313] = 250;
    exp_62_ram[3314] = 251;
    exp_62_ram[3315] = 251;
    exp_62_ram[3316] = 251;
    exp_62_ram[3317] = 251;
    exp_62_ram[3318] = 252;
    exp_62_ram[3319] = 252;
    exp_62_ram[3320] = 1;
    exp_62_ram[3321] = 0;
    exp_62_ram[3322] = 1;
    exp_62_ram[3323] = 1;
    exp_62_ram[3324] = 0;
    exp_62_ram[3325] = 0;
    exp_62_ram[3326] = 0;
    exp_62_ram[3327] = 0;
    exp_62_ram[3328] = 2;
    exp_62_ram[3329] = 248;
    exp_62_ram[3330] = 7;
    exp_62_ram[3331] = 7;
    exp_62_ram[3332] = 7;
    exp_62_ram[3333] = 7;
    exp_62_ram[3334] = 6;
    exp_62_ram[3335] = 6;
    exp_62_ram[3336] = 6;
    exp_62_ram[3337] = 6;
    exp_62_ram[3338] = 5;
    exp_62_ram[3339] = 5;
    exp_62_ram[3340] = 8;
    exp_62_ram[3341] = 0;
    exp_62_ram[3342] = 246;
    exp_62_ram[3343] = 8;
    exp_62_ram[3344] = 8;
    exp_62_ram[3345] = 8;
    exp_62_ram[3346] = 9;
    exp_62_ram[3347] = 9;
    exp_62_ram[3348] = 10;
    exp_62_ram[3349] = 248;
    exp_62_ram[3350] = 0;
    exp_62_ram[3351] = 0;
    exp_62_ram[3352] = 252;
    exp_62_ram[3353] = 253;
    exp_62_ram[3354] = 249;
    exp_62_ram[3355] = 0;
    exp_62_ram[3356] = 0;
    exp_62_ram[3357] = 252;
    exp_62_ram[3358] = 252;
    exp_62_ram[3359] = 253;
    exp_62_ram[3360] = 253;
    exp_62_ram[3361] = 220;
    exp_62_ram[3362] = 0;
    exp_62_ram[3363] = 0;
    exp_62_ram[3364] = 0;
    exp_62_ram[3365] = 225;
    exp_62_ram[3366] = 0;
    exp_62_ram[3367] = 252;
    exp_62_ram[3368] = 252;
    exp_62_ram[3369] = 0;
    exp_62_ram[3370] = 40;
    exp_62_ram[3371] = 0;
    exp_62_ram[3372] = 65;
    exp_62_ram[3373] = 0;
    exp_62_ram[3374] = 253;
    exp_62_ram[3375] = 253;
    exp_62_ram[3376] = 0;
    exp_62_ram[3377] = 0;
    exp_62_ram[3378] = 1;
    exp_62_ram[3379] = 0;
    exp_62_ram[3380] = 0;
    exp_62_ram[3381] = 0;
    exp_62_ram[3382] = 0;
    exp_62_ram[3383] = 0;
    exp_62_ram[3384] = 253;
    exp_62_ram[3385] = 253;
    exp_62_ram[3386] = 0;
    exp_62_ram[3387] = 0;
    exp_62_ram[3388] = 0;
    exp_62_ram[3389] = 0;
    exp_62_ram[3390] = 0;
    exp_62_ram[3391] = 0;
    exp_62_ram[3392] = 252;
    exp_62_ram[3393] = 252;
    exp_62_ram[3394] = 0;
    exp_62_ram[3395] = 42;
    exp_62_ram[3396] = 246;
    exp_62_ram[3397] = 252;
    exp_62_ram[3398] = 252;
    exp_62_ram[3399] = 0;
    exp_62_ram[3400] = 188;
    exp_62_ram[3401] = 246;
    exp_62_ram[3402] = 246;
    exp_62_ram[3403] = 246;
    exp_62_ram[3404] = 246;
    exp_62_ram[3405] = 247;
    exp_62_ram[3406] = 247;
    exp_62_ram[3407] = 247;
    exp_62_ram[3408] = 247;
    exp_62_ram[3409] = 248;
    exp_62_ram[3410] = 0;
    exp_62_ram[3411] = 1;
    exp_62_ram[3412] = 1;
    exp_62_ram[3413] = 0;
    exp_62_ram[3414] = 0;
    exp_62_ram[3415] = 0;
    exp_62_ram[3416] = 0;
    exp_62_ram[3417] = 0;
    exp_62_ram[3418] = 2;
    exp_62_ram[3419] = 253;
    exp_62_ram[3420] = 253;
    exp_62_ram[3421] = 205;
    exp_62_ram[3422] = 0;
    exp_62_ram[3423] = 0;
    exp_62_ram[3424] = 42;
    exp_62_ram[3425] = 2;
    exp_62_ram[3426] = 0;
    exp_62_ram[3427] = 42;
    exp_62_ram[3428] = 0;
    exp_62_ram[3429] = 9;
    exp_62_ram[3430] = 9;
    exp_62_ram[3431] = 9;
    exp_62_ram[3432] = 9;
    exp_62_ram[3433] = 8;
    exp_62_ram[3434] = 10;
    exp_62_ram[3435] = 0;
    exp_62_ram[3436] = 253;
    exp_62_ram[3437] = 2;
    exp_62_ram[3438] = 2;
    exp_62_ram[3439] = 3;
    exp_62_ram[3440] = 252;
    exp_62_ram[3441] = 254;
    exp_62_ram[3442] = 253;
    exp_62_ram[3443] = 216;
    exp_62_ram[3444] = 0;
    exp_62_ram[3445] = 254;
    exp_62_ram[3446] = 254;
    exp_62_ram[3447] = 253;
    exp_62_ram[3448] = 0;
    exp_62_ram[3449] = 2;
    exp_62_ram[3450] = 254;
    exp_62_ram[3451] = 0;
    exp_62_ram[3452] = 0;
    exp_62_ram[3453] = 0;
    exp_62_ram[3454] = 0;
    exp_62_ram[3455] = 254;
    exp_62_ram[3456] = 254;
    exp_62_ram[3457] = 254;
    exp_62_ram[3458] = 0;
    exp_62_ram[3459] = 253;
    exp_62_ram[3460] = 254;
    exp_62_ram[3461] = 251;
    exp_62_ram[3462] = 0;
    exp_62_ram[3463] = 254;
    exp_62_ram[3464] = 0;
    exp_62_ram[3465] = 2;
    exp_62_ram[3466] = 2;
    exp_62_ram[3467] = 3;
    exp_62_ram[3468] = 0;
    exp_62_ram[3469] = 255;
    exp_62_ram[3470] = 0;
    exp_62_ram[3471] = 0;
    exp_62_ram[3472] = 1;
    exp_62_ram[3473] = 0;
    exp_62_ram[3474] = 9;
    exp_62_ram[3475] = 0;
    exp_62_ram[3476] = 246;
    exp_62_ram[3477] = 0;
    exp_62_ram[3478] = 0;
    exp_62_ram[3479] = 0;
    exp_62_ram[3480] = 0;
    exp_62_ram[3481] = 1;
    exp_62_ram[3482] = 0;
    exp_62_ram[3483] = 253;
    exp_62_ram[3484] = 2;
    exp_62_ram[3485] = 2;
    exp_62_ram[3486] = 3;
    exp_62_ram[3487] = 3;
    exp_62_ram[3488] = 3;
    exp_62_ram[3489] = 252;
    exp_62_ram[3490] = 197;
    exp_62_ram[3491] = 254;
    exp_62_ram[3492] = 254;
    exp_62_ram[3493] = 0;
    exp_62_ram[3494] = 196;
    exp_62_ram[3495] = 0;
    exp_62_ram[3496] = 0;
    exp_62_ram[3497] = 254;
    exp_62_ram[3498] = 254;
    exp_62_ram[3499] = 64;
    exp_62_ram[3500] = 0;
    exp_62_ram[3501] = 1;
    exp_62_ram[3502] = 64;
    exp_62_ram[3503] = 65;
    exp_62_ram[3504] = 0;
    exp_62_ram[3505] = 253;
    exp_62_ram[3506] = 0;
    exp_62_ram[3507] = 0;
    exp_62_ram[3508] = 0;
    exp_62_ram[3509] = 0;
    exp_62_ram[3510] = 252;
    exp_62_ram[3511] = 0;
    exp_62_ram[3512] = 0;
    exp_62_ram[3513] = 0;
    exp_62_ram[3514] = 0;
    exp_62_ram[3515] = 0;
    exp_62_ram[3516] = 250;
    exp_62_ram[3517] = 0;
    exp_62_ram[3518] = 0;
    exp_62_ram[3519] = 2;
    exp_62_ram[3520] = 2;
    exp_62_ram[3521] = 2;
    exp_62_ram[3522] = 2;
    exp_62_ram[3523] = 3;
    exp_62_ram[3524] = 0;
    exp_62_ram[3525] = 255;
    exp_62_ram[3526] = 0;
    exp_62_ram[3527] = 0;
    exp_62_ram[3528] = 1;
    exp_62_ram[3529] = 0;
    exp_62_ram[3530] = 142;
    exp_62_ram[3531] = 246;
    exp_62_ram[3532] = 0;
    exp_62_ram[3533] = 0;
    exp_62_ram[3534] = 0;
    exp_62_ram[3535] = 1;
    exp_62_ram[3536] = 0;
    exp_62_ram[3537] = 254;
    exp_62_ram[3538] = 0;
    exp_62_ram[3539] = 0;
    exp_62_ram[3540] = 2;
    exp_62_ram[3541] = 0;
    exp_62_ram[3542] = 143;
    exp_62_ram[3543] = 243;
    exp_62_ram[3544] = 0;
    exp_62_ram[3545] = 254;
    exp_62_ram[3546] = 254;
    exp_62_ram[3547] = 11;
    exp_62_ram[3548] = 254;
    exp_62_ram[3549] = 0;
    exp_62_ram[3550] = 145;
    exp_62_ram[3551] = 241;
    exp_62_ram[3552] = 3;
    exp_62_ram[3553] = 254;
    exp_62_ram[3554] = 0;
    exp_62_ram[3555] = 254;
    exp_62_ram[3556] = 0;
    exp_62_ram[3557] = 9;
    exp_62_ram[3558] = 0;
    exp_62_ram[3559] = 254;
    exp_62_ram[3560] = 190;
    exp_62_ram[3561] = 0;
    exp_62_ram[3562] = 9;
    exp_62_ram[3563] = 0;
    exp_62_ram[3564] = 2;
    exp_62_ram[3565] = 0;
    exp_62_ram[3566] = 235;
    exp_62_ram[3567] = 254;
    exp_62_ram[3568] = 7;
    exp_62_ram[3569] = 252;
    exp_62_ram[3570] = 3;
    exp_62_ram[3571] = 254;
    exp_62_ram[3572] = 64;
    exp_62_ram[3573] = 254;
    exp_62_ram[3574] = 0;
    exp_62_ram[3575] = 9;
    exp_62_ram[3576] = 0;
    exp_62_ram[3577] = 254;
    exp_62_ram[3578] = 185;
    exp_62_ram[3579] = 0;
    exp_62_ram[3580] = 9;
    exp_62_ram[3581] = 0;
    exp_62_ram[3582] = 2;
    exp_62_ram[3583] = 0;
    exp_62_ram[3584] = 230;
    exp_62_ram[3585] = 254;
    exp_62_ram[3586] = 0;
    exp_62_ram[3587] = 252;
    exp_62_ram[3588] = 254;
    exp_62_ram[3589] = 0;
    exp_62_ram[3590] = 254;
    exp_62_ram[3591] = 254;
    exp_62_ram[3592] = 0;
    exp_62_ram[3593] = 244;
    exp_62_ram[3594] = 0;
    exp_62_ram[3595] = 9;
    exp_62_ram[3596] = 0;
    exp_62_ram[3597] = 0;
    exp_62_ram[3598] = 180;
    exp_62_ram[3599] = 0;
    exp_62_ram[3600] = 1;
    exp_62_ram[3601] = 1;
    exp_62_ram[3602] = 2;
    exp_62_ram[3603] = 0;
    exp_62_ram[3604] = 249;
    exp_62_ram[3605] = 6;
    exp_62_ram[3606] = 6;
    exp_62_ram[3607] = 7;
    exp_62_ram[3608] = 7;
    exp_62_ram[3609] = 5;
    exp_62_ram[3610] = 5;
    exp_62_ram[3611] = 5;
    exp_62_ram[3612] = 5;
    exp_62_ram[3613] = 5;
    exp_62_ram[3614] = 5;
    exp_62_ram[3615] = 5;
    exp_62_ram[3616] = 5;
    exp_62_ram[3617] = 7;
    exp_62_ram[3618] = 0;
    exp_62_ram[3619] = 250;
    exp_62_ram[3620] = 0;
    exp_62_ram[3621] = 0;
    exp_62_ram[3622] = 250;
    exp_62_ram[3623] = 250;
    exp_62_ram[3624] = 164;
    exp_62_ram[3625] = 252;
    exp_62_ram[3626] = 252;
    exp_62_ram[3627] = 252;
    exp_62_ram[3628] = 6;
    exp_62_ram[3629] = 251;
    exp_62_ram[3630] = 18;
    exp_62_ram[3631] = 103;
    exp_62_ram[3632] = 2;
    exp_62_ram[3633] = 250;
    exp_62_ram[3634] = 251;
    exp_62_ram[3635] = 18;
    exp_62_ram[3636] = 103;
    exp_62_ram[3637] = 2;
    exp_62_ram[3638] = 250;
    exp_62_ram[3639] = 251;
    exp_62_ram[3640] = 18;
    exp_62_ram[3641] = 103;
    exp_62_ram[3642] = 2;
    exp_62_ram[3643] = 250;
    exp_62_ram[3644] = 251;
    exp_62_ram[3645] = 18;
    exp_62_ram[3646] = 103;
    exp_62_ram[3647] = 2;
    exp_62_ram[3648] = 250;
    exp_62_ram[3649] = 252;
    exp_62_ram[3650] = 0;
    exp_62_ram[3651] = 252;
    exp_62_ram[3652] = 157;
    exp_62_ram[3653] = 0;
    exp_62_ram[3654] = 0;
    exp_62_ram[3655] = 252;
    exp_62_ram[3656] = 252;
    exp_62_ram[3657] = 64;
    exp_62_ram[3658] = 0;
    exp_62_ram[3659] = 1;
    exp_62_ram[3660] = 64;
    exp_62_ram[3661] = 65;
    exp_62_ram[3662] = 0;
    exp_62_ram[3663] = 0;
    exp_62_ram[3664] = 9;
    exp_62_ram[3665] = 250;
    exp_62_ram[3666] = 250;
    exp_62_ram[3667] = 250;
    exp_62_ram[3668] = 250;
    exp_62_ram[3669] = 0;
    exp_62_ram[3670] = 0;
    exp_62_ram[3671] = 244;
    exp_62_ram[3672] = 0;
    exp_62_ram[3673] = 0;
    exp_62_ram[3674] = 0;
    exp_62_ram[3675] = 0;
    exp_62_ram[3676] = 0;
    exp_62_ram[3677] = 244;
    exp_62_ram[3678] = 252;
    exp_62_ram[3679] = 0;
    exp_62_ram[3680] = 145;
    exp_62_ram[3681] = 209;
    exp_62_ram[3682] = 149;
    exp_62_ram[3683] = 252;
    exp_62_ram[3684] = 252;
    exp_62_ram[3685] = 252;
    exp_62_ram[3686] = 18;
    exp_62_ram[3687] = 251;
    exp_62_ram[3688] = 251;
    exp_62_ram[3689] = 18;
    exp_62_ram[3690] = 103;
    exp_62_ram[3691] = 2;
    exp_62_ram[3692] = 0;
    exp_62_ram[3693] = 2;
    exp_62_ram[3694] = 0;
    exp_62_ram[3695] = 18;
    exp_62_ram[3696] = 103;
    exp_62_ram[3697] = 2;
    exp_62_ram[3698] = 2;
    exp_62_ram[3699] = 0;
    exp_62_ram[3700] = 1;
    exp_62_ram[3701] = 0;
    exp_62_ram[3702] = 251;
    exp_62_ram[3703] = 251;
    exp_62_ram[3704] = 251;
    exp_62_ram[3705] = 251;
    exp_62_ram[3706] = 18;
    exp_62_ram[3707] = 103;
    exp_62_ram[3708] = 2;
    exp_62_ram[3709] = 0;
    exp_62_ram[3710] = 2;
    exp_62_ram[3711] = 0;
    exp_62_ram[3712] = 18;
    exp_62_ram[3713] = 103;
    exp_62_ram[3714] = 2;
    exp_62_ram[3715] = 2;
    exp_62_ram[3716] = 0;
    exp_62_ram[3717] = 1;
    exp_62_ram[3718] = 0;
    exp_62_ram[3719] = 251;
    exp_62_ram[3720] = 251;
    exp_62_ram[3721] = 251;
    exp_62_ram[3722] = 251;
    exp_62_ram[3723] = 18;
    exp_62_ram[3724] = 103;
    exp_62_ram[3725] = 2;
    exp_62_ram[3726] = 0;
    exp_62_ram[3727] = 2;
    exp_62_ram[3728] = 0;
    exp_62_ram[3729] = 18;
    exp_62_ram[3730] = 103;
    exp_62_ram[3731] = 2;
    exp_62_ram[3732] = 2;
    exp_62_ram[3733] = 0;
    exp_62_ram[3734] = 1;
    exp_62_ram[3735] = 0;
    exp_62_ram[3736] = 251;
    exp_62_ram[3737] = 251;
    exp_62_ram[3738] = 251;
    exp_62_ram[3739] = 251;
    exp_62_ram[3740] = 18;
    exp_62_ram[3741] = 103;
    exp_62_ram[3742] = 2;
    exp_62_ram[3743] = 0;
    exp_62_ram[3744] = 2;
    exp_62_ram[3745] = 0;
    exp_62_ram[3746] = 18;
    exp_62_ram[3747] = 103;
    exp_62_ram[3748] = 2;
    exp_62_ram[3749] = 2;
    exp_62_ram[3750] = 0;
    exp_62_ram[3751] = 1;
    exp_62_ram[3752] = 0;
    exp_62_ram[3753] = 251;
    exp_62_ram[3754] = 251;
    exp_62_ram[3755] = 252;
    exp_62_ram[3756] = 0;
    exp_62_ram[3757] = 252;
    exp_62_ram[3758] = 130;
    exp_62_ram[3759] = 0;
    exp_62_ram[3760] = 0;
    exp_62_ram[3761] = 252;
    exp_62_ram[3762] = 252;
    exp_62_ram[3763] = 64;
    exp_62_ram[3764] = 0;
    exp_62_ram[3765] = 1;
    exp_62_ram[3766] = 64;
    exp_62_ram[3767] = 65;
    exp_62_ram[3768] = 0;
    exp_62_ram[3769] = 0;
    exp_62_ram[3770] = 9;
    exp_62_ram[3771] = 250;
    exp_62_ram[3772] = 250;
    exp_62_ram[3773] = 250;
    exp_62_ram[3774] = 250;
    exp_62_ram[3775] = 0;
    exp_62_ram[3776] = 0;
    exp_62_ram[3777] = 232;
    exp_62_ram[3778] = 0;
    exp_62_ram[3779] = 0;
    exp_62_ram[3780] = 0;
    exp_62_ram[3781] = 0;
    exp_62_ram[3782] = 0;
    exp_62_ram[3783] = 232;
    exp_62_ram[3784] = 252;
    exp_62_ram[3785] = 0;
    exp_62_ram[3786] = 148;
    exp_62_ram[3787] = 182;
    exp_62_ram[3788] = 251;
    exp_62_ram[3789] = 252;
    exp_62_ram[3790] = 252;
    exp_62_ram[3791] = 252;
    exp_62_ram[3792] = 6;
    exp_62_ram[3793] = 251;
    exp_62_ram[3794] = 18;
    exp_62_ram[3795] = 103;
    exp_62_ram[3796] = 2;
    exp_62_ram[3797] = 250;
    exp_62_ram[3798] = 251;
    exp_62_ram[3799] = 18;
    exp_62_ram[3800] = 103;
    exp_62_ram[3801] = 2;
    exp_62_ram[3802] = 250;
    exp_62_ram[3803] = 251;
    exp_62_ram[3804] = 18;
    exp_62_ram[3805] = 103;
    exp_62_ram[3806] = 2;
    exp_62_ram[3807] = 250;
    exp_62_ram[3808] = 251;
    exp_62_ram[3809] = 18;
    exp_62_ram[3810] = 103;
    exp_62_ram[3811] = 2;
    exp_62_ram[3812] = 250;
    exp_62_ram[3813] = 252;
    exp_62_ram[3814] = 0;
    exp_62_ram[3815] = 252;
    exp_62_ram[3816] = 244;
    exp_62_ram[3817] = 0;
    exp_62_ram[3818] = 0;
    exp_62_ram[3819] = 252;
    exp_62_ram[3820] = 252;
    exp_62_ram[3821] = 64;
    exp_62_ram[3822] = 0;
    exp_62_ram[3823] = 1;
    exp_62_ram[3824] = 64;
    exp_62_ram[3825] = 65;
    exp_62_ram[3826] = 0;
    exp_62_ram[3827] = 0;
    exp_62_ram[3828] = 9;
    exp_62_ram[3829] = 248;
    exp_62_ram[3830] = 248;
    exp_62_ram[3831] = 249;
    exp_62_ram[3832] = 249;
    exp_62_ram[3833] = 0;
    exp_62_ram[3834] = 0;
    exp_62_ram[3835] = 244;
    exp_62_ram[3836] = 0;
    exp_62_ram[3837] = 0;
    exp_62_ram[3838] = 0;
    exp_62_ram[3839] = 0;
    exp_62_ram[3840] = 0;
    exp_62_ram[3841] = 244;
    exp_62_ram[3842] = 252;
    exp_62_ram[3843] = 0;
    exp_62_ram[3844] = 151;
    exp_62_ram[3845] = 168;
    exp_62_ram[3846] = 236;
    exp_62_ram[3847] = 252;
    exp_62_ram[3848] = 252;
    exp_62_ram[3849] = 252;
    exp_62_ram[3850] = 13;
    exp_62_ram[3851] = 251;
    exp_62_ram[3852] = 251;
    exp_62_ram[3853] = 18;
    exp_62_ram[3854] = 103;
    exp_62_ram[3855] = 0;
    exp_62_ram[3856] = 0;
    exp_62_ram[3857] = 0;
    exp_62_ram[3858] = 196;
    exp_62_ram[3859] = 0;
    exp_62_ram[3860] = 0;
    exp_62_ram[3861] = 250;
    exp_62_ram[3862] = 250;
    exp_62_ram[3863] = 251;
    exp_62_ram[3864] = 251;
    exp_62_ram[3865] = 18;
    exp_62_ram[3866] = 103;
    exp_62_ram[3867] = 0;
    exp_62_ram[3868] = 0;
    exp_62_ram[3869] = 0;
    exp_62_ram[3870] = 193;
    exp_62_ram[3871] = 0;
    exp_62_ram[3872] = 0;
    exp_62_ram[3873] = 250;
    exp_62_ram[3874] = 250;
    exp_62_ram[3875] = 251;
    exp_62_ram[3876] = 251;
    exp_62_ram[3877] = 18;
    exp_62_ram[3878] = 103;
    exp_62_ram[3879] = 0;
    exp_62_ram[3880] = 0;
    exp_62_ram[3881] = 0;
    exp_62_ram[3882] = 190;
    exp_62_ram[3883] = 0;
    exp_62_ram[3884] = 0;
    exp_62_ram[3885] = 250;
    exp_62_ram[3886] = 250;
    exp_62_ram[3887] = 251;
    exp_62_ram[3888] = 251;
    exp_62_ram[3889] = 18;
    exp_62_ram[3890] = 103;
    exp_62_ram[3891] = 0;
    exp_62_ram[3892] = 0;
    exp_62_ram[3893] = 0;
    exp_62_ram[3894] = 187;
    exp_62_ram[3895] = 0;
    exp_62_ram[3896] = 0;
    exp_62_ram[3897] = 250;
    exp_62_ram[3898] = 250;
    exp_62_ram[3899] = 252;
    exp_62_ram[3900] = 0;
    exp_62_ram[3901] = 252;
    exp_62_ram[3902] = 222;
    exp_62_ram[3903] = 0;
    exp_62_ram[3904] = 0;
    exp_62_ram[3905] = 252;
    exp_62_ram[3906] = 252;
    exp_62_ram[3907] = 64;
    exp_62_ram[3908] = 0;
    exp_62_ram[3909] = 1;
    exp_62_ram[3910] = 64;
    exp_62_ram[3911] = 65;
    exp_62_ram[3912] = 0;
    exp_62_ram[3913] = 0;
    exp_62_ram[3914] = 9;
    exp_62_ram[3915] = 0;
    exp_62_ram[3916] = 0;
    exp_62_ram[3917] = 0;
    exp_62_ram[3918] = 0;
    exp_62_ram[3919] = 238;
    exp_62_ram[3920] = 0;
    exp_62_ram[3921] = 0;
    exp_62_ram[3922] = 0;
    exp_62_ram[3923] = 0;
    exp_62_ram[3924] = 0;
    exp_62_ram[3925] = 236;
    exp_62_ram[3926] = 252;
    exp_62_ram[3927] = 0;
    exp_62_ram[3928] = 153;
    exp_62_ram[3929] = 147;
    exp_62_ram[3930] = 0;
    exp_62_ram[3931] = 6;
    exp_62_ram[3932] = 6;
    exp_62_ram[3933] = 6;
    exp_62_ram[3934] = 6;
    exp_62_ram[3935] = 5;
    exp_62_ram[3936] = 5;
    exp_62_ram[3937] = 5;
    exp_62_ram[3938] = 5;
    exp_62_ram[3939] = 4;
    exp_62_ram[3940] = 4;
    exp_62_ram[3941] = 4;
    exp_62_ram[3942] = 4;
    exp_62_ram[3943] = 7;
    exp_62_ram[3944] = 0;
    exp_62_ram[3945] = 250;
    exp_62_ram[3946] = 4;
    exp_62_ram[3947] = 4;
    exp_62_ram[3948] = 5;
    exp_62_ram[3949] = 5;
    exp_62_ram[3950] = 5;
    exp_62_ram[3951] = 5;
    exp_62_ram[3952] = 6;
    exp_62_ram[3953] = 0;
    exp_62_ram[3954] = 156;
    exp_62_ram[3955] = 140;
    exp_62_ram[3956] = 134;
    exp_62_ram[3957] = 0;
    exp_62_ram[3958] = 137;
    exp_62_ram[3959] = 252;
    exp_62_ram[3960] = 0;
    exp_62_ram[3961] = 156;
    exp_62_ram[3962] = 139;
    exp_62_ram[3963] = 132;
    exp_62_ram[3964] = 0;
    exp_62_ram[3965] = 255;
    exp_62_ram[3966] = 252;
    exp_62_ram[3967] = 0;
    exp_62_ram[3968] = 157;
    exp_62_ram[3969] = 137;
    exp_62_ram[3970] = 130;
    exp_62_ram[3971] = 0;
    exp_62_ram[3972] = 250;
    exp_62_ram[3973] = 0;
    exp_62_ram[3974] = 157;
    exp_62_ram[3975] = 135;
    exp_62_ram[3976] = 129;
    exp_62_ram[3977] = 0;
    exp_62_ram[3978] = 250;
    exp_62_ram[3979] = 0;
    exp_62_ram[3980] = 158;
    exp_62_ram[3981] = 134;
    exp_62_ram[3982] = 255;
    exp_62_ram[3983] = 0;
    exp_62_ram[3984] = 250;
    exp_62_ram[3985] = 3;
    exp_62_ram[3986] = 250;
    exp_62_ram[3987] = 0;
    exp_62_ram[3988] = 252;
    exp_62_ram[3989] = 251;
    exp_62_ram[3990] = 0;
    exp_62_ram[3991] = 150;
    exp_62_ram[3992] = 0;
    exp_62_ram[3993] = 0;
    exp_62_ram[3994] = 250;
    exp_62_ram[3995] = 250;
    exp_62_ram[3996] = 250;
    exp_62_ram[3997] = 250;
    exp_62_ram[3998] = 0;
    exp_62_ram[3999] = 0;
    exp_62_ram[4000] = 211;
    exp_62_ram[4001] = 198;
    exp_62_ram[4002] = 252;
    exp_62_ram[4003] = 252;
    exp_62_ram[4004] = 252;
    exp_62_ram[4005] = 13;
    exp_62_ram[4006] = 0;
    exp_62_ram[4007] = 196;
    exp_62_ram[4008] = 0;
    exp_62_ram[4009] = 0;
    exp_62_ram[4010] = 253;
    exp_62_ram[4011] = 253;
    exp_62_ram[4012] = 0;
    exp_62_ram[4013] = 0;
    exp_62_ram[4014] = 203;
    exp_62_ram[4015] = 0;
    exp_62_ram[4016] = 0;
    exp_62_ram[4017] = 0;
    exp_62_ram[4018] = 9;
    exp_62_ram[4019] = 0;
    exp_62_ram[4020] = 237;
    exp_62_ram[4021] = 0;
    exp_62_ram[4022] = 0;
    exp_62_ram[4023] = 0;
    exp_62_ram[4024] = 0;
    exp_62_ram[4025] = 0;
    exp_62_ram[4026] = 0;
    exp_62_ram[4027] = 221;
    exp_62_ram[4028] = 0;
    exp_62_ram[4029] = 250;
    exp_62_ram[4030] = 0;
    exp_62_ram[4031] = 9;
    exp_62_ram[4032] = 0;
    exp_62_ram[4033] = 0;
    exp_62_ram[4034] = 253;
    exp_62_ram[4035] = 253;
    exp_62_ram[4036] = 1;
    exp_62_ram[4037] = 0;
    exp_62_ram[4038] = 0;
    exp_62_ram[4039] = 1;
    exp_62_ram[4040] = 0;
    exp_62_ram[4041] = 0;
    exp_62_ram[4042] = 252;
    exp_62_ram[4043] = 252;
    exp_62_ram[4044] = 0;
    exp_62_ram[4045] = 185;
    exp_62_ram[4046] = 0;
    exp_62_ram[4047] = 0;
    exp_62_ram[4048] = 250;
    exp_62_ram[4049] = 250;
    exp_62_ram[4050] = 250;
    exp_62_ram[4051] = 0;
    exp_62_ram[4052] = 149;
    exp_62_ram[4053] = 0;
    exp_62_ram[4054] = 0;
    exp_62_ram[4055] = 208;
    exp_62_ram[4056] = 253;
    exp_62_ram[4057] = 0;
    exp_62_ram[4058] = 252;
    exp_62_ram[4059] = 253;
    exp_62_ram[4060] = 6;
    exp_62_ram[4061] = 242;
    exp_62_ram[4062] = 0;
    exp_62_ram[4063] = 0;
    exp_62_ram[4064] = 5;
    exp_62_ram[4065] = 5;
    exp_62_ram[4066] = 5;
    exp_62_ram[4067] = 5;
    exp_62_ram[4068] = 4;
    exp_62_ram[4069] = 4;
    exp_62_ram[4070] = 6;
    exp_62_ram[4071] = 0;
    exp_62_ram[4072] = 254;
    exp_62_ram[4073] = 0;
    exp_62_ram[4074] = 0;
    exp_62_ram[4075] = 2;
    exp_62_ram[4076] = 0;
    exp_62_ram[4077] = 159;
    exp_62_ram[4078] = 238;
    exp_62_ram[4079] = 0;
    exp_62_ram[4080] = 160;
    exp_62_ram[4081] = 237;
    exp_62_ram[4082] = 0;
    exp_62_ram[4083] = 161;
    exp_62_ram[4084] = 236;
    exp_62_ram[4085] = 0;
    exp_62_ram[4086] = 162;
    exp_62_ram[4087] = 235;
    exp_62_ram[4088] = 0;
    exp_62_ram[4089] = 164;
    exp_62_ram[4090] = 235;
    exp_62_ram[4091] = 189;
    exp_62_ram[4092] = 0;
    exp_62_ram[4093] = 254;
    exp_62_ram[4094] = 254;
    exp_62_ram[4095] = 6;
    exp_62_ram[4096] = 4;
    exp_62_ram[4097] = 6;
    exp_62_ram[4098] = 250;
    exp_62_ram[4099] = 6;
    exp_62_ram[4100] = 2;
    exp_62_ram[4101] = 6;
    exp_62_ram[4102] = 248;
    exp_62_ram[4103] = 6;
    exp_62_ram[4104] = 0;
    exp_62_ram[4105] = 6;
    exp_62_ram[4106] = 0;
    exp_62_ram[4107] = 2;
    exp_62_ram[4108] = 238;
    exp_62_ram[4109] = 1;
    exp_62_ram[4110] = 240;
    exp_62_ram[4111] = 1;
    exp_62_ram[4112] = 129;
    exp_62_ram[4113] = 0;
    exp_62_ram[4114] = 213;
    exp_62_ram[4115] = 0;
    exp_62_ram[4116] = 246;
    exp_62_ram[4117] = 0;
    exp_62_ram[4118] = 0;
    exp_62_ram[4119] = 2;
    exp_62_ram[4120] = 255;
    exp_62_ram[4121] = 2;
    exp_62_ram[4122] = 0;
    exp_62_ram[4123] = 0;
    exp_62_ram[4124] = 0;
    exp_62_ram[4125] = 64;
    exp_62_ram[4126] = 1;
    exp_62_ram[4127] = 0;
    exp_62_ram[4128] = 254;
    exp_62_ram[4129] = 255;
    exp_62_ram[4130] = 0;
    exp_62_ram[4131] = 254;
    exp_62_ram[4132] = 2;
    exp_62_ram[4133] = 128;
    exp_62_ram[4134] = 128;
    exp_62_ram[4135] = 128;
    exp_62_ram[4136] = 0;
    exp_62_ram[4137] = 0;
    exp_62_ram[4138] = 0;
    exp_62_ram[4139] = 0;
    exp_62_ram[4140] = 0;
    exp_62_ram[4141] = 0;
    exp_62_ram[4142] = 0;
    exp_62_ram[4143] = 0;
    exp_62_ram[4144] = 0;
    exp_62_ram[4145] = 0;
    exp_62_ram[4146] = 0;
    exp_62_ram[4147] = 0;
    exp_62_ram[4148] = 0;
    exp_62_ram[4149] = 0;
    exp_62_ram[4150] = 0;
    exp_62_ram[4151] = 0;
    exp_62_ram[4152] = 0;
    exp_62_ram[4153] = 0;
    exp_62_ram[4154] = 0;
    exp_62_ram[4155] = 0;
    exp_62_ram[4156] = 0;
    exp_62_ram[4157] = 0;
    exp_62_ram[4158] = 0;
    exp_62_ram[4159] = 0;
    exp_62_ram[4160] = 0;
    exp_62_ram[4161] = 0;
    exp_62_ram[4162] = 0;
    exp_62_ram[4163] = 0;
    exp_62_ram[4164] = 0;
    exp_62_ram[4165] = 0;
    exp_62_ram[4166] = 0;
    exp_62_ram[4167] = 0;
    exp_62_ram[4168] = 0;
    exp_62_ram[4169] = 0;
    exp_62_ram[4170] = 0;
    exp_62_ram[4171] = 0;
    exp_62_ram[4172] = 0;
    exp_62_ram[4173] = 0;
    exp_62_ram[4174] = 0;
    exp_62_ram[4175] = 0;
    exp_62_ram[4176] = 0;
    exp_62_ram[4177] = 0;
    exp_62_ram[4178] = 0;
    exp_62_ram[4179] = 0;
    exp_62_ram[4180] = 0;
    exp_62_ram[4181] = 0;
    exp_62_ram[4182] = 0;
    exp_62_ram[4183] = 0;
    exp_62_ram[4184] = 0;
    exp_62_ram[4185] = 0;
    exp_62_ram[4186] = 0;
    exp_62_ram[4187] = 0;
    exp_62_ram[4188] = 0;
    exp_62_ram[4189] = 0;
    exp_62_ram[4190] = 0;
    exp_62_ram[4191] = 0;
    exp_62_ram[4192] = 0;
    exp_62_ram[4193] = 0;
    exp_62_ram[4194] = 0;
    exp_62_ram[4195] = 0;
    exp_62_ram[4196] = 0;
    exp_62_ram[4197] = 0;
    exp_62_ram[4198] = 0;
    exp_62_ram[4199] = 0;
    exp_62_ram[4200] = 0;
    exp_62_ram[4201] = 0;
    exp_62_ram[4202] = 0;
    exp_62_ram[4203] = 0;
    exp_62_ram[4204] = 0;
    exp_62_ram[4205] = 0;
    exp_62_ram[4206] = 0;
    exp_62_ram[4207] = 0;
    exp_62_ram[4208] = 0;
    exp_62_ram[4209] = 0;
    exp_62_ram[4210] = 0;
    exp_62_ram[4211] = 0;
    exp_62_ram[4212] = 0;
    exp_62_ram[4213] = 0;
    exp_62_ram[4214] = 0;
    exp_62_ram[4215] = 0;
    exp_62_ram[4216] = 0;
    exp_62_ram[4217] = 0;
    exp_62_ram[4218] = 0;
    exp_62_ram[4219] = 0;
    exp_62_ram[4220] = 0;
    exp_62_ram[4221] = 0;
    exp_62_ram[4222] = 0;
    exp_62_ram[4223] = 0;
    exp_62_ram[4224] = 0;
    exp_62_ram[4225] = 0;
    exp_62_ram[4226] = 0;
    exp_62_ram[4227] = 0;
    exp_62_ram[4228] = 0;
    exp_62_ram[4229] = 0;
    exp_62_ram[4230] = 0;
    exp_62_ram[4231] = 0;
    exp_62_ram[4232] = 0;
    exp_62_ram[4233] = 0;
    exp_62_ram[4234] = 0;
    exp_62_ram[4235] = 0;
    exp_62_ram[4236] = 0;
    exp_62_ram[4237] = 0;
    exp_62_ram[4238] = 0;
    exp_62_ram[4239] = 0;
    exp_62_ram[4240] = 0;
    exp_62_ram[4241] = 0;
    exp_62_ram[4242] = 0;
    exp_62_ram[4243] = 0;
    exp_62_ram[4244] = 0;
    exp_62_ram[4245] = 0;
    exp_62_ram[4246] = 0;
    exp_62_ram[4247] = 0;
    exp_62_ram[4248] = 0;
    exp_62_ram[4249] = 0;
    exp_62_ram[4250] = 0;
    exp_62_ram[4251] = 0;
    exp_62_ram[4252] = 0;
    exp_62_ram[4253] = 0;
    exp_62_ram[4254] = 0;
    exp_62_ram[4255] = 0;
    exp_62_ram[4256] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_60) begin
      exp_62_ram[exp_56] <= exp_58;
    end
  end
  assign exp_62 = exp_62_ram[exp_57];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_88) begin
        exp_62_ram[exp_84] <= exp_86;
    end
  end
  assign exp_90 = exp_62_ram[exp_85];
  assign exp_61 = exp_129;
  assign exp_129 = 1;
  assign exp_57 = exp_128;
  assign exp_128 = exp_18[31:2];
  assign exp_18 = exp_9;
  assign exp_60 = exp_124;
  assign exp_124 = exp_122 & exp_123;
  assign exp_122 = exp_22 & exp_23;
  assign exp_123 = exp_24[3:3];
  assign exp_24 = exp_13;
  assign exp_13 = exp_404;
  assign exp_404 = exp_685;

  reg [3:0] exp_685_reg;
  always@(*) begin
    case (exp_537)
      0:exp_685_reg <= exp_672;
      1:exp_685_reg <= exp_677;
      2:exp_685_reg <= exp_678;
      3:exp_685_reg <= exp_679;
      4:exp_685_reg <= exp_680;
      5:exp_685_reg <= exp_681;
      6:exp_685_reg <= exp_682;
      7:exp_685_reg <= exp_683;
      default:exp_685_reg <= exp_684;
    endcase
  end
  assign exp_685 = exp_685_reg;
  assign exp_684 = 0;
  assign exp_672 = exp_668 << exp_671;
  assign exp_668 = 1;
  assign exp_671 = exp_670 + exp_669;
  assign exp_670 = 0;
  assign exp_669 = exp_605[1:0];
  assign exp_677 = exp_673 << exp_676;
  assign exp_673 = 3;
  assign exp_676 = exp_675 + exp_674;
  assign exp_675 = 0;
  assign exp_674 = exp_605[1:1];
  assign exp_678 = 15;
  assign exp_679 = 0;
  assign exp_680 = 0;
  assign exp_681 = 0;
  assign exp_682 = 0;
  assign exp_683 = 0;
  assign exp_56 = exp_120;
  assign exp_120 = exp_18[31:2];
  assign exp_58 = exp_121;
  assign exp_121 = exp_19[31:24];
  assign exp_19 = exp_10;
  assign exp_10 = exp_399;
  assign exp_399 = exp_667;

  reg [31:0] exp_667_reg;
  always@(*) begin
    case (exp_537)
      0:exp_667_reg <= exp_654;
      1:exp_667_reg <= exp_658;
      2:exp_667_reg <= exp_660;
      3:exp_667_reg <= exp_661;
      4:exp_667_reg <= exp_662;
      5:exp_667_reg <= exp_663;
      6:exp_667_reg <= exp_664;
      7:exp_667_reg <= exp_665;
      default:exp_667_reg <= exp_666;
    endcase
  end
  assign exp_667 = exp_667_reg;
  assign exp_666 = 0;

  reg [31:0] exp_654_reg;
  always@(*) begin
    case (exp_608)
      0:exp_654_reg <= exp_640;
      1:exp_654_reg <= exp_648;
      2:exp_654_reg <= exp_650;
      3:exp_654_reg <= exp_652;
      default:exp_654_reg <= exp_653;
    endcase
  end
  assign exp_654 = exp_654_reg;
  assign exp_653 = 0;
  assign exp_640 = exp_639;
  assign exp_639 = exp_638 + exp_637;
  assign exp_638 = 0;
  assign exp_637 = exp_527[7:0];

      reg [31:0] exp_527_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_527_reg <= exp_470;
        end
      end
      assign exp_527 = exp_527_reg;
      assign exp_648 = exp_640 << exp_647;
  assign exp_647 = 8;
  assign exp_650 = exp_640 << exp_649;
  assign exp_649 = 16;
  assign exp_652 = exp_640 << exp_651;
  assign exp_651 = 24;

  reg [31:0] exp_658_reg;
  always@(*) begin
    case (exp_611)
      0:exp_658_reg <= exp_644;
      1:exp_658_reg <= exp_656;
      default:exp_658_reg <= exp_657;
    endcase
  end
  assign exp_658 = exp_658_reg;
  assign exp_611 = exp_610 + exp_609;
  assign exp_610 = 0;
  assign exp_609 = exp_605[1:1];
  assign exp_657 = 0;
  assign exp_644 = exp_643;
  assign exp_643 = exp_642 + exp_641;
  assign exp_642 = 0;
  assign exp_641 = exp_527[15:0];
  assign exp_656 = exp_644 << exp_655;
  assign exp_655 = 16;
  assign exp_660 = exp_659 + exp_646;
  assign exp_659 = 0;
  assign exp_646 = exp_645 + exp_527;
  assign exp_645 = 0;
  assign exp_661 = 0;
  assign exp_662 = 0;
  assign exp_663 = 0;
  assign exp_664 = 0;
  assign exp_665 = 0;

  //Create RAM
  reg [7:0] exp_55_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_55_ram[0] = 0;
    exp_55_ram[1] = 0;
    exp_55_ram[2] = 0;
    exp_55_ram[3] = 0;
    exp_55_ram[4] = 0;
    exp_55_ram[5] = 0;
    exp_55_ram[6] = 0;
    exp_55_ram[7] = 0;
    exp_55_ram[8] = 0;
    exp_55_ram[9] = 0;
    exp_55_ram[10] = 0;
    exp_55_ram[11] = 0;
    exp_55_ram[12] = 0;
    exp_55_ram[13] = 0;
    exp_55_ram[14] = 0;
    exp_55_ram[15] = 0;
    exp_55_ram[16] = 0;
    exp_55_ram[17] = 0;
    exp_55_ram[18] = 0;
    exp_55_ram[19] = 0;
    exp_55_ram[20] = 0;
    exp_55_ram[21] = 0;
    exp_55_ram[22] = 0;
    exp_55_ram[23] = 0;
    exp_55_ram[24] = 0;
    exp_55_ram[25] = 0;
    exp_55_ram[26] = 0;
    exp_55_ram[27] = 0;
    exp_55_ram[28] = 0;
    exp_55_ram[29] = 0;
    exp_55_ram[30] = 0;
    exp_55_ram[31] = 0;
    exp_55_ram[32] = 1;
    exp_55_ram[33] = 208;
    exp_55_ram[34] = 0;
    exp_55_ram[35] = 5;
    exp_55_ram[36] = 5;
    exp_55_ram[37] = 6;
    exp_55_ram[38] = 6;
    exp_55_ram[39] = 8;
    exp_55_ram[40] = 6;
    exp_55_ram[41] = 0;
    exp_55_ram[42] = 6;
    exp_55_ram[43] = 197;
    exp_55_ram[44] = 1;
    exp_55_ram[45] = 230;
    exp_55_ram[46] = 240;
    exp_55_ram[47] = 199;
    exp_55_ram[48] = 55;
    exp_55_ram[49] = 230;
    exp_55_ram[50] = 166;
    exp_55_ram[51] = 6;
    exp_55_ram[52] = 0;
    exp_55_ram[53] = 230;
    exp_55_ram[54] = 229;
    exp_55_ram[55] = 229;
    exp_55_ram[56] = 215;
    exp_55_ram[57] = 232;
    exp_55_ram[58] = 214;
    exp_55_ram[59] = 183;
    exp_55_ram[60] = 216;
    exp_55_ram[61] = 8;
    exp_55_ram[62] = 21;
    exp_55_ram[63] = 8;
    exp_55_ram[64] = 6;
    exp_55_ram[65] = 3;
    exp_55_ram[66] = 21;
    exp_55_ram[67] = 6;
    exp_55_ram[68] = 214;
    exp_55_ram[69] = 7;
    exp_55_ram[70] = 247;
    exp_55_ram[71] = 183;
    exp_55_ram[72] = 7;
    exp_55_ram[73] = 246;
    exp_55_ram[74] = 7;
    exp_55_ram[75] = 183;
    exp_55_ram[76] = 230;
    exp_55_ram[77] = 7;
    exp_55_ram[78] = 183;
    exp_55_ram[79] = 23;
    exp_55_ram[80] = 3;
    exp_55_ram[81] = 3;
    exp_55_ram[82] = 23;
    exp_55_ram[83] = 7;
    exp_55_ram[84] = 103;
    exp_55_ram[85] = 246;
    exp_55_ram[86] = 7;
    exp_55_ram[87] = 211;
    exp_55_ram[88] = 104;
    exp_55_ram[89] = 247;
    exp_55_ram[90] = 3;
    exp_55_ram[91] = 211;
    exp_55_ram[92] = 231;
    exp_55_ram[93] = 5;
    exp_55_ram[94] = 197;
    exp_55_ram[95] = 0;
    exp_55_ram[96] = 64;
    exp_55_ram[97] = 0;
    exp_55_ram[98] = 0;
    exp_55_ram[99] = 166;
    exp_55_ram[100] = 128;
    exp_55_ram[101] = 31;
    exp_55_ram[102] = 6;
    exp_55_ram[103] = 16;
    exp_55_ram[104] = 199;
    exp_55_ram[105] = 1;
    exp_55_ram[106] = 232;
    exp_55_ram[107] = 240;
    exp_55_ram[108] = 7;
    exp_55_ram[109] = 128;
    exp_55_ram[110] = 168;
    exp_55_ram[111] = 230;
    exp_55_ram[112] = 6;
    exp_55_ram[113] = 0;
    exp_55_ram[114] = 167;
    exp_55_ram[115] = 230;
    exp_55_ram[116] = 230;
    exp_55_ram[117] = 7;
    exp_55_ram[118] = 16;
    exp_55_ram[119] = 8;
    exp_55_ram[120] = 8;
    exp_55_ram[121] = 6;
    exp_55_ram[122] = 3;
    exp_55_ram[123] = 23;
    exp_55_ram[124] = 23;
    exp_55_ram[125] = 6;
    exp_55_ram[126] = 230;
    exp_55_ram[127] = 246;
    exp_55_ram[128] = 7;
    exp_55_ram[129] = 199;
    exp_55_ram[130] = 7;
    exp_55_ram[131] = 247;
    exp_55_ram[132] = 7;
    exp_55_ram[133] = 199;
    exp_55_ram[134] = 231;
    exp_55_ram[135] = 7;
    exp_55_ram[136] = 199;
    exp_55_ram[137] = 23;
    exp_55_ram[138] = 3;
    exp_55_ram[139] = 3;
    exp_55_ram[140] = 23;
    exp_55_ram[141] = 7;
    exp_55_ram[142] = 103;
    exp_55_ram[143] = 230;
    exp_55_ram[144] = 7;
    exp_55_ram[145] = 211;
    exp_55_ram[146] = 104;
    exp_55_ram[147] = 247;
    exp_55_ram[148] = 3;
    exp_55_ram[149] = 211;
    exp_55_ram[150] = 231;
    exp_55_ram[151] = 5;
    exp_55_ram[152] = 197;
    exp_55_ram[153] = 0;
    exp_55_ram[154] = 0;
    exp_55_ram[155] = 0;
    exp_55_ram[156] = 232;
    exp_55_ram[157] = 128;
    exp_55_ram[158] = 31;
    exp_55_ram[159] = 216;
    exp_55_ram[160] = 231;
    exp_55_ram[161] = 216;
    exp_55_ram[162] = 215;
    exp_55_ram[163] = 232;
    exp_55_ram[164] = 8;
    exp_55_ram[165] = 247;
    exp_55_ram[166] = 21;
    exp_55_ram[167] = 8;
    exp_55_ram[168] = 7;
    exp_55_ram[169] = 6;
    exp_55_ram[170] = 21;
    exp_55_ram[171] = 7;
    exp_55_ram[172] = 183;
    exp_55_ram[173] = 167;
    exp_55_ram[174] = 5;
    exp_55_ram[175] = 215;
    exp_55_ram[176] = 7;
    exp_55_ram[177] = 245;
    exp_55_ram[178] = 7;
    exp_55_ram[179] = 215;
    exp_55_ram[180] = 229;
    exp_55_ram[181] = 7;
    exp_55_ram[182] = 215;
    exp_55_ram[183] = 22;
    exp_55_ram[184] = 6;
    exp_55_ram[185] = 6;
    exp_55_ram[186] = 22;
    exp_55_ram[187] = 7;
    exp_55_ram[188] = 215;
    exp_55_ram[189] = 199;
    exp_55_ram[190] = 6;
    exp_55_ram[191] = 167;
    exp_55_ram[192] = 7;
    exp_55_ram[193] = 246;
    exp_55_ram[194] = 7;
    exp_55_ram[195] = 167;
    exp_55_ram[196] = 230;
    exp_55_ram[197] = 7;
    exp_55_ram[198] = 5;
    exp_55_ram[199] = 167;
    exp_55_ram[200] = 229;
    exp_55_ram[201] = 159;
    exp_55_ram[202] = 213;
    exp_55_ram[203] = 1;
    exp_55_ram[204] = 230;
    exp_55_ram[205] = 240;
    exp_55_ram[206] = 215;
    exp_55_ram[207] = 53;
    exp_55_ram[208] = 0;
    exp_55_ram[209] = 182;
    exp_55_ram[210] = 7;
    exp_55_ram[211] = 167;
    exp_55_ram[212] = 7;
    exp_55_ram[213] = 0;
    exp_55_ram[214] = 183;
    exp_55_ram[215] = 229;
    exp_55_ram[216] = 229;
    exp_55_ram[217] = 16;
    exp_55_ram[218] = 246;
    exp_55_ram[219] = 200;
    exp_55_ram[220] = 21;
    exp_55_ram[221] = 31;
    exp_55_ram[222] = 0;
    exp_55_ram[223] = 0;
    exp_55_ram[224] = 230;
    exp_55_ram[225] = 128;
    exp_55_ram[226] = 159;
    exp_55_ram[227] = 230;
    exp_55_ram[228] = 182;
    exp_55_ram[229] = 216;
    exp_55_ram[230] = 231;
    exp_55_ram[231] = 8;
    exp_55_ram[232] = 222;
    exp_55_ram[233] = 183;
    exp_55_ram[234] = 232;
    exp_55_ram[235] = 182;
    exp_55_ram[236] = 247;
    exp_55_ram[237] = 8;
    exp_55_ram[238] = 7;
    exp_55_ram[239] = 6;
    exp_55_ram[240] = 222;
    exp_55_ram[241] = 6;
    exp_55_ram[242] = 230;
    exp_55_ram[243] = 199;
    exp_55_ram[244] = 14;
    exp_55_ram[245] = 231;
    exp_55_ram[246] = 7;
    exp_55_ram[247] = 254;
    exp_55_ram[248] = 7;
    exp_55_ram[249] = 231;
    exp_55_ram[250] = 238;
    exp_55_ram[251] = 7;
    exp_55_ram[252] = 231;
    exp_55_ram[253] = 215;
    exp_55_ram[254] = 215;
    exp_55_ram[255] = 6;
    exp_55_ram[256] = 231;
    exp_55_ram[257] = 6;
    exp_55_ram[258] = 7;
    exp_55_ram[259] = 246;
    exp_55_ram[260] = 7;
    exp_55_ram[261] = 199;
    exp_55_ram[262] = 7;
    exp_55_ram[263] = 247;
    exp_55_ram[264] = 7;
    exp_55_ram[265] = 199;
    exp_55_ram[266] = 231;
    exp_55_ram[267] = 7;
    exp_55_ram[268] = 5;
    exp_55_ram[269] = 1;
    exp_55_ram[270] = 197;
    exp_55_ram[271] = 254;
    exp_55_ram[272] = 213;
    exp_55_ram[273] = 5;
    exp_55_ram[274] = 211;
    exp_55_ram[275] = 3;
    exp_55_ram[276] = 199;
    exp_55_ram[277] = 216;
    exp_55_ram[278] = 214;
    exp_55_ram[279] = 14;
    exp_55_ram[280] = 104;
    exp_55_ram[281] = 216;
    exp_55_ram[282] = 7;
    exp_55_ram[283] = 102;
    exp_55_ram[284] = 215;
    exp_55_ram[285] = 214;
    exp_55_ram[286] = 7;
    exp_55_ram[287] = 198;
    exp_55_ram[288] = 199;
    exp_55_ram[289] = 199;
    exp_55_ram[290] = 1;
    exp_55_ram[291] = 247;
    exp_55_ram[292] = 247;
    exp_55_ram[293] = 7;
    exp_55_ram[294] = 254;
    exp_55_ram[295] = 184;
    exp_55_ram[296] = 199;
    exp_55_ram[297] = 0;
    exp_55_ram[298] = 232;
    exp_55_ram[299] = 245;
    exp_55_ram[300] = 223;
    exp_55_ram[301] = 0;
    exp_55_ram[302] = 0;
    exp_55_ram[303] = 159;
    exp_55_ram[304] = 16;
    exp_55_ram[305] = 247;
    exp_55_ram[306] = 69;
    exp_55_ram[307] = 183;
    exp_55_ram[308] = 5;
    exp_55_ram[309] = 5;
    exp_55_ram[310] = 248;
    exp_55_ram[311] = 245;
    exp_55_ram[312] = 240;
    exp_55_ram[313] = 70;
    exp_55_ram[314] = 215;
    exp_55_ram[315] = 6;
    exp_55_ram[316] = 245;
    exp_55_ram[317] = 246;
    exp_55_ram[318] = 216;
    exp_55_ram[319] = 248;
    exp_55_ram[320] = 14;
    exp_55_ram[321] = 32;
    exp_55_ram[322] = 0;
    exp_55_ram[323] = 213;
    exp_55_ram[324] = 199;
    exp_55_ram[325] = 14;
    exp_55_ram[326] = 8;
    exp_55_ram[327] = 248;
    exp_55_ram[328] = 23;
    exp_55_ram[329] = 5;
    exp_55_ram[330] = 199;
    exp_55_ram[331] = 6;
    exp_55_ram[332] = 7;
    exp_55_ram[333] = 213;
    exp_55_ram[334] = 5;
    exp_55_ram[335] = 5;
    exp_55_ram[336] = 240;
    exp_55_ram[337] = 0;
    exp_55_ram[338] = 240;
    exp_55_ram[339] = 6;
    exp_55_ram[340] = 6;
    exp_55_ram[341] = 0;
    exp_55_ram[342] = 184;
    exp_55_ram[343] = 5;
    exp_55_ram[344] = 0;
    exp_55_ram[345] = 23;
    exp_55_ram[346] = 232;
    exp_55_ram[347] = 110;
    exp_55_ram[348] = 195;
    exp_55_ram[349] = 0;
    exp_55_ram[350] = 0;
    exp_55_ram[351] = 16;
    exp_55_ram[352] = 0;
    exp_55_ram[353] = 7;
    exp_55_ram[354] = 95;
    exp_55_ram[355] = 232;
    exp_55_ram[356] = 95;
    exp_55_ram[357] = 5;
    exp_55_ram[358] = 5;
    exp_55_ram[359] = 0;
    exp_55_ram[360] = 159;
    exp_55_ram[361] = 1;
    exp_55_ram[362] = 129;
    exp_55_ram[363] = 17;
    exp_55_ram[364] = 5;
    exp_55_ram[365] = 5;
    exp_55_ram[366] = 64;
    exp_55_ram[367] = 224;
    exp_55_ram[368] = 160;
    exp_55_ram[369] = 167;
    exp_55_ram[370] = 167;
    exp_55_ram[371] = 176;
    exp_55_ram[372] = 167;
    exp_55_ram[373] = 85;
    exp_55_ram[374] = 244;
    exp_55_ram[375] = 164;
    exp_55_ram[376] = 193;
    exp_55_ram[377] = 4;
    exp_55_ram[378] = 199;
    exp_55_ram[379] = 129;
    exp_55_ram[380] = 71;
    exp_55_ram[381] = 199;
    exp_55_ram[382] = 247;
    exp_55_ram[383] = 6;
    exp_55_ram[384] = 1;
    exp_55_ram[385] = 0;
    exp_55_ram[386] = 85;
    exp_55_ram[387] = 244;
    exp_55_ram[388] = 0;
    exp_55_ram[389] = 223;
    exp_55_ram[390] = 0;
    exp_55_ram[391] = 0;
    exp_55_ram[392] = 31;
    exp_55_ram[393] = 1;
    exp_55_ram[394] = 17;
    exp_55_ram[395] = 129;
    exp_55_ram[396] = 145;
    exp_55_ram[397] = 33;
    exp_55_ram[398] = 49;
    exp_55_ram[399] = 65;
    exp_55_ram[400] = 181;
    exp_55_ram[401] = 7;
    exp_55_ram[402] = 5;
    exp_55_ram[403] = 5;
    exp_55_ram[404] = 5;
    exp_55_ram[405] = 5;
    exp_55_ram[406] = 5;
    exp_55_ram[407] = 0;
    exp_55_ram[408] = 5;
    exp_55_ram[409] = 224;
    exp_55_ram[410] = 58;
    exp_55_ram[411] = 48;
    exp_55_ram[412] = 71;
    exp_55_ram[413] = 176;
    exp_55_ram[414] = 4;
    exp_55_ram[415] = 55;
    exp_55_ram[416] = 160;
    exp_55_ram[417] = 55;
    exp_55_ram[418] = 176;
    exp_55_ram[419] = 89;
    exp_55_ram[420] = 52;
    exp_55_ram[421] = 148;
    exp_55_ram[422] = 233;
    exp_55_ram[423] = 180;
    exp_55_ram[424] = 228;
    exp_55_ram[425] = 193;
    exp_55_ram[426] = 129;
    exp_55_ram[427] = 196;
    exp_55_ram[428] = 74;
    exp_55_ram[429] = 197;
    exp_55_ram[430] = 186;
    exp_55_ram[431] = 65;
    exp_55_ram[432] = 1;
    exp_55_ram[433] = 193;
    exp_55_ram[434] = 129;
    exp_55_ram[435] = 7;
    exp_55_ram[436] = 7;
    exp_55_ram[437] = 1;
    exp_55_ram[438] = 0;
    exp_55_ram[439] = 0;
    exp_55_ram[440] = 5;
    exp_55_ram[441] = 31;
    exp_55_ram[442] = 89;
    exp_55_ram[443] = 180;
    exp_55_ram[444] = 0;
    exp_55_ram[445] = 31;
    exp_55_ram[446] = 96;
    exp_55_ram[447] = 71;
    exp_55_ram[448] = 137;
    exp_55_ram[449] = 4;
    exp_55_ram[450] = 9;
    exp_55_ram[451] = 128;
    exp_55_ram[452] = 181;
    exp_55_ram[453] = 128;
    exp_55_ram[454] = 160;
    exp_55_ram[455] = 9;
    exp_55_ram[456] = 4;
    exp_55_ram[457] = 54;
    exp_55_ram[458] = 64;
    exp_55_ram[459] = 164;
    exp_55_ram[460] = 5;
    exp_55_ram[461] = 128;
    exp_55_ram[462] = 4;
    exp_55_ram[463] = 9;
    exp_55_ram[464] = 55;
    exp_55_ram[465] = 112;
    exp_55_ram[466] = 55;
    exp_55_ram[467] = 137;
    exp_55_ram[468] = 233;
    exp_55_ram[469] = 128;
    exp_55_ram[470] = 57;
    exp_55_ram[471] = 36;
    exp_55_ram[472] = 185;
    exp_55_ram[473] = 228;
    exp_55_ram[474] = 128;
    exp_55_ram[475] = 247;
    exp_55_ram[476] = 229;
    exp_55_ram[477] = 119;
    exp_55_ram[478] = 7;
    exp_55_ram[479] = 247;
    exp_55_ram[480] = 64;
    exp_55_ram[481] = 215;
    exp_55_ram[482] = 71;
    exp_55_ram[483] = 247;
    exp_55_ram[484] = 245;
    exp_55_ram[485] = 7;
    exp_55_ram[486] = 128;
    exp_55_ram[487] = 229;
    exp_55_ram[488] = 7;
    exp_55_ram[489] = 128;
    exp_55_ram[490] = 247;
    exp_55_ram[491] = 240;
    exp_55_ram[492] = 229;
    exp_55_ram[493] = 58;
    exp_55_ram[494] = 55;
    exp_55_ram[495] = 213;
    exp_55_ram[496] = 245;
    exp_55_ram[497] = 53;
    exp_55_ram[498] = 223;
    exp_55_ram[499] = 137;
    exp_55_ram[500] = 180;
    exp_55_ram[501] = 0;
    exp_55_ram[502] = 31;
    exp_55_ram[503] = 0;
    exp_55_ram[504] = 0;
    exp_55_ram[505] = 0;
    exp_55_ram[506] = 223;
    exp_55_ram[507] = 6;
    exp_55_ram[508] = 0;
    exp_55_ram[509] = 199;
    exp_55_ram[510] = 240;
    exp_55_ram[511] = 6;
    exp_55_ram[512] = 0;
    exp_55_ram[513] = 165;
    exp_55_ram[514] = 7;
    exp_55_ram[515] = 0;
    exp_55_ram[516] = 197;
    exp_55_ram[517] = 197;
    exp_55_ram[518] = 245;
    exp_55_ram[519] = 181;
    exp_55_ram[520] = 159;
    exp_55_ram[521] = 6;
    exp_55_ram[522] = 0;
    exp_55_ram[523] = 199;
    exp_55_ram[524] = 240;
    exp_55_ram[525] = 6;
    exp_55_ram[526] = 0;
    exp_55_ram[527] = 181;
    exp_55_ram[528] = 7;
    exp_55_ram[529] = 0;
    exp_55_ram[530] = 197;
    exp_55_ram[531] = 197;
    exp_55_ram[532] = 245;
    exp_55_ram[533] = 165;
    exp_55_ram[534] = 159;
    exp_55_ram[535] = 1;
    exp_55_ram[536] = 245;
    exp_55_ram[537] = 240;
    exp_55_ram[538] = 167;
    exp_55_ram[539] = 55;
    exp_55_ram[540] = 0;
    exp_55_ram[541] = 0;
    exp_55_ram[542] = 246;
    exp_55_ram[543] = 245;
    exp_55_ram[544] = 7;
    exp_55_ram[545] = 167;
    exp_55_ram[546] = 5;
    exp_55_ram[547] = 166;
    exp_55_ram[548] = 0;
    exp_55_ram[549] = 0;
    exp_55_ram[550] = 0;
    exp_55_ram[551] = 229;
    exp_55_ram[552] = 128;
    exp_55_ram[553] = 223;
    exp_55_ram[554] = 110;
    exp_55_ram[555] = 84;
    exp_55_ram[556] = 101;
    exp_55_ram[557] = 117;
    exp_55_ram[558] = 83;
    exp_55_ram[559] = 0;
    exp_55_ram[560] = 110;
    exp_55_ram[561] = 77;
    exp_55_ram[562] = 112;
    exp_55_ram[563] = 121;
    exp_55_ram[564] = 74;
    exp_55_ram[565] = 117;
    exp_55_ram[566] = 112;
    exp_55_ram[567] = 78;
    exp_55_ram[568] = 101;
    exp_55_ram[569] = 0;
    exp_55_ram[570] = 108;
    exp_55_ram[571] = 87;
    exp_55_ram[572] = 100;
    exp_55_ram[573] = 0;
    exp_55_ram[574] = 110;
    exp_55_ram[575] = 103;
    exp_55_ram[576] = 105;
    exp_55_ram[577] = 32;
    exp_55_ram[578] = 101;
    exp_55_ram[579] = 101;
    exp_55_ram[580] = 46;
    exp_55_ram[581] = 0;
    exp_55_ram[582] = 10;
    exp_55_ram[583] = 32;
    exp_55_ram[584] = 98;
    exp_55_ram[585] = 105;
    exp_55_ram[586] = 103;
    exp_55_ram[587] = 109;
    exp_55_ram[588] = 105;
    exp_55_ram[589] = 101;
    exp_55_ram[590] = 110;
    exp_55_ram[591] = 115;
    exp_55_ram[592] = 110;
    exp_55_ram[593] = 0;
    exp_55_ram[594] = 32;
    exp_55_ram[595] = 98;
    exp_55_ram[596] = 105;
    exp_55_ram[597] = 103;
    exp_55_ram[598] = 109;
    exp_55_ram[599] = 105;
    exp_55_ram[600] = 101;
    exp_55_ram[601] = 110;
    exp_55_ram[602] = 115;
    exp_55_ram[603] = 110;
    exp_55_ram[604] = 0;
    exp_55_ram[605] = 32;
    exp_55_ram[606] = 98;
    exp_55_ram[607] = 105;
    exp_55_ram[608] = 103;
    exp_55_ram[609] = 100;
    exp_55_ram[610] = 100;
    exp_55_ram[611] = 105;
    exp_55_ram[612] = 32;
    exp_55_ram[613] = 111;
    exp_55_ram[614] = 0;
    exp_55_ram[615] = 32;
    exp_55_ram[616] = 98;
    exp_55_ram[617] = 105;
    exp_55_ram[618] = 103;
    exp_55_ram[619] = 100;
    exp_55_ram[620] = 100;
    exp_55_ram[621] = 105;
    exp_55_ram[622] = 32;
    exp_55_ram[623] = 111;
    exp_55_ram[624] = 0;
    exp_55_ram[625] = 97;
    exp_55_ram[626] = 0;
    exp_55_ram[627] = 110;
    exp_55_ram[628] = 10;
    exp_55_ram[629] = 121;
    exp_55_ram[630] = 0;
    exp_55_ram[631] = 117;
    exp_55_ram[632] = 0;
    exp_55_ram[633] = 110;
    exp_55_ram[634] = 58;
    exp_55_ram[635] = 0;
    exp_55_ram[636] = 104;
    exp_55_ram[637] = 45;
    exp_55_ram[638] = 101;
    exp_55_ram[639] = 0;
    exp_55_ram[640] = 41;
    exp_55_ram[641] = 108;
    exp_55_ram[642] = 87;
    exp_55_ram[643] = 100;
    exp_55_ram[644] = 0;
    exp_55_ram[645] = 32;
    exp_55_ram[646] = 103;
    exp_55_ram[647] = 82;
    exp_55_ram[648] = 114;
    exp_55_ram[649] = 0;
    exp_55_ram[650] = 32;
    exp_55_ram[651] = 116;
    exp_55_ram[652] = 108;
    exp_55_ram[653] = 108;
    exp_55_ram[654] = 116;
    exp_55_ram[655] = 10;
    exp_55_ram[656] = 32;
    exp_55_ram[657] = 108;
    exp_55_ram[658] = 111;
    exp_55_ram[659] = 0;
    exp_55_ram[660] = 2;
    exp_55_ram[661] = 3;
    exp_55_ram[662] = 4;
    exp_55_ram[663] = 4;
    exp_55_ram[664] = 5;
    exp_55_ram[665] = 5;
    exp_55_ram[666] = 5;
    exp_55_ram[667] = 5;
    exp_55_ram[668] = 6;
    exp_55_ram[669] = 6;
    exp_55_ram[670] = 6;
    exp_55_ram[671] = 6;
    exp_55_ram[672] = 6;
    exp_55_ram[673] = 6;
    exp_55_ram[674] = 6;
    exp_55_ram[675] = 6;
    exp_55_ram[676] = 7;
    exp_55_ram[677] = 7;
    exp_55_ram[678] = 7;
    exp_55_ram[679] = 7;
    exp_55_ram[680] = 7;
    exp_55_ram[681] = 7;
    exp_55_ram[682] = 7;
    exp_55_ram[683] = 7;
    exp_55_ram[684] = 7;
    exp_55_ram[685] = 7;
    exp_55_ram[686] = 7;
    exp_55_ram[687] = 7;
    exp_55_ram[688] = 7;
    exp_55_ram[689] = 7;
    exp_55_ram[690] = 7;
    exp_55_ram[691] = 7;
    exp_55_ram[692] = 8;
    exp_55_ram[693] = 8;
    exp_55_ram[694] = 8;
    exp_55_ram[695] = 8;
    exp_55_ram[696] = 8;
    exp_55_ram[697] = 8;
    exp_55_ram[698] = 8;
    exp_55_ram[699] = 8;
    exp_55_ram[700] = 8;
    exp_55_ram[701] = 8;
    exp_55_ram[702] = 8;
    exp_55_ram[703] = 8;
    exp_55_ram[704] = 8;
    exp_55_ram[705] = 8;
    exp_55_ram[706] = 8;
    exp_55_ram[707] = 8;
    exp_55_ram[708] = 8;
    exp_55_ram[709] = 8;
    exp_55_ram[710] = 8;
    exp_55_ram[711] = 8;
    exp_55_ram[712] = 8;
    exp_55_ram[713] = 8;
    exp_55_ram[714] = 8;
    exp_55_ram[715] = 8;
    exp_55_ram[716] = 8;
    exp_55_ram[717] = 8;
    exp_55_ram[718] = 8;
    exp_55_ram[719] = 8;
    exp_55_ram[720] = 8;
    exp_55_ram[721] = 8;
    exp_55_ram[722] = 8;
    exp_55_ram[723] = 8;
    exp_55_ram[724] = 1;
    exp_55_ram[725] = 129;
    exp_55_ram[726] = 1;
    exp_55_ram[727] = 164;
    exp_55_ram[728] = 196;
    exp_55_ram[729] = 244;
    exp_55_ram[730] = 196;
    exp_55_ram[731] = 7;
    exp_55_ram[732] = 7;
    exp_55_ram[733] = 193;
    exp_55_ram[734] = 1;
    exp_55_ram[735] = 0;
    exp_55_ram[736] = 1;
    exp_55_ram[737] = 129;
    exp_55_ram[738] = 1;
    exp_55_ram[739] = 164;
    exp_55_ram[740] = 180;
    exp_55_ram[741] = 132;
    exp_55_ram[742] = 244;
    exp_55_ram[743] = 196;
    exp_55_ram[744] = 196;
    exp_55_ram[745] = 231;
    exp_55_ram[746] = 196;
    exp_55_ram[747] = 7;
    exp_55_ram[748] = 193;
    exp_55_ram[749] = 1;
    exp_55_ram[750] = 0;
    exp_55_ram[751] = 1;
    exp_55_ram[752] = 17;
    exp_55_ram[753] = 129;
    exp_55_ram[754] = 1;
    exp_55_ram[755] = 0;
    exp_55_ram[756] = 71;
    exp_55_ram[757] = 7;
    exp_55_ram[758] = 159;
    exp_55_ram[759] = 5;
    exp_55_ram[760] = 7;
    exp_55_ram[761] = 193;
    exp_55_ram[762] = 129;
    exp_55_ram[763] = 1;
    exp_55_ram[764] = 0;
    exp_55_ram[765] = 1;
    exp_55_ram[766] = 17;
    exp_55_ram[767] = 129;
    exp_55_ram[768] = 1;
    exp_55_ram[769] = 164;
    exp_55_ram[770] = 180;
    exp_55_ram[771] = 4;
    exp_55_ram[772] = 128;
    exp_55_ram[773] = 196;
    exp_55_ram[774] = 23;
    exp_55_ram[775] = 228;
    exp_55_ram[776] = 196;
    exp_55_ram[777] = 247;
    exp_55_ram[778] = 7;
    exp_55_ram[779] = 132;
    exp_55_ram[780] = 7;
    exp_55_ram[781] = 223;
    exp_55_ram[782] = 196;
    exp_55_ram[783] = 196;
    exp_55_ram[784] = 247;
    exp_55_ram[785] = 7;
    exp_55_ram[786] = 7;
    exp_55_ram[787] = 196;
    exp_55_ram[788] = 7;
    exp_55_ram[789] = 193;
    exp_55_ram[790] = 129;
    exp_55_ram[791] = 1;
    exp_55_ram[792] = 0;
    exp_55_ram[793] = 1;
    exp_55_ram[794] = 17;
    exp_55_ram[795] = 129;
    exp_55_ram[796] = 1;
    exp_55_ram[797] = 164;
    exp_55_ram[798] = 0;
    exp_55_ram[799] = 135;
    exp_55_ram[800] = 7;
    exp_55_ram[801] = 196;
    exp_55_ram[802] = 223;
    exp_55_ram[803] = 0;
    exp_55_ram[804] = 135;
    exp_55_ram[805] = 7;
    exp_55_ram[806] = 160;
    exp_55_ram[807] = 95;
    exp_55_ram[808] = 0;
    exp_55_ram[809] = 7;
    exp_55_ram[810] = 193;
    exp_55_ram[811] = 129;
    exp_55_ram[812] = 1;
    exp_55_ram[813] = 0;
    exp_55_ram[814] = 1;
    exp_55_ram[815] = 129;
    exp_55_ram[816] = 1;
    exp_55_ram[817] = 5;
    exp_55_ram[818] = 180;
    exp_55_ram[819] = 196;
    exp_55_ram[820] = 212;
    exp_55_ram[821] = 244;
    exp_55_ram[822] = 0;
    exp_55_ram[823] = 193;
    exp_55_ram[824] = 1;
    exp_55_ram[825] = 0;
    exp_55_ram[826] = 1;
    exp_55_ram[827] = 17;
    exp_55_ram[828] = 129;
    exp_55_ram[829] = 1;
    exp_55_ram[830] = 5;
    exp_55_ram[831] = 180;
    exp_55_ram[832] = 196;
    exp_55_ram[833] = 212;
    exp_55_ram[834] = 244;
    exp_55_ram[835] = 244;
    exp_55_ram[836] = 7;
    exp_55_ram[837] = 244;
    exp_55_ram[838] = 7;
    exp_55_ram[839] = 192;
    exp_55_ram[840] = 0;
    exp_55_ram[841] = 193;
    exp_55_ram[842] = 129;
    exp_55_ram[843] = 1;
    exp_55_ram[844] = 0;
    exp_55_ram[845] = 1;
    exp_55_ram[846] = 129;
    exp_55_ram[847] = 1;
    exp_55_ram[848] = 164;
    exp_55_ram[849] = 180;
    exp_55_ram[850] = 196;
    exp_55_ram[851] = 244;
    exp_55_ram[852] = 0;
    exp_55_ram[853] = 196;
    exp_55_ram[854] = 23;
    exp_55_ram[855] = 244;
    exp_55_ram[856] = 196;
    exp_55_ram[857] = 7;
    exp_55_ram[858] = 7;
    exp_55_ram[859] = 132;
    exp_55_ram[860] = 247;
    exp_55_ram[861] = 228;
    exp_55_ram[862] = 7;
    exp_55_ram[863] = 196;
    exp_55_ram[864] = 196;
    exp_55_ram[865] = 247;
    exp_55_ram[866] = 7;
    exp_55_ram[867] = 193;
    exp_55_ram[868] = 1;
    exp_55_ram[869] = 0;
    exp_55_ram[870] = 1;
    exp_55_ram[871] = 129;
    exp_55_ram[872] = 1;
    exp_55_ram[873] = 5;
    exp_55_ram[874] = 244;
    exp_55_ram[875] = 244;
    exp_55_ram[876] = 240;
    exp_55_ram[877] = 231;
    exp_55_ram[878] = 244;
    exp_55_ram[879] = 144;
    exp_55_ram[880] = 231;
    exp_55_ram[881] = 16;
    exp_55_ram[882] = 128;
    exp_55_ram[883] = 0;
    exp_55_ram[884] = 23;
    exp_55_ram[885] = 247;
    exp_55_ram[886] = 7;
    exp_55_ram[887] = 193;
    exp_55_ram[888] = 1;
    exp_55_ram[889] = 0;
    exp_55_ram[890] = 1;
    exp_55_ram[891] = 17;
    exp_55_ram[892] = 129;
    exp_55_ram[893] = 1;
    exp_55_ram[894] = 164;
    exp_55_ram[895] = 4;
    exp_55_ram[896] = 0;
    exp_55_ram[897] = 196;
    exp_55_ram[898] = 7;
    exp_55_ram[899] = 39;
    exp_55_ram[900] = 231;
    exp_55_ram[901] = 23;
    exp_55_ram[902] = 7;
    exp_55_ram[903] = 196;
    exp_55_ram[904] = 7;
    exp_55_ram[905] = 23;
    exp_55_ram[906] = 196;
    exp_55_ram[907] = 215;
    exp_55_ram[908] = 7;
    exp_55_ram[909] = 246;
    exp_55_ram[910] = 7;
    exp_55_ram[911] = 244;
    exp_55_ram[912] = 196;
    exp_55_ram[913] = 7;
    exp_55_ram[914] = 7;
    exp_55_ram[915] = 7;
    exp_55_ram[916] = 159;
    exp_55_ram[917] = 5;
    exp_55_ram[918] = 7;
    exp_55_ram[919] = 196;
    exp_55_ram[920] = 7;
    exp_55_ram[921] = 193;
    exp_55_ram[922] = 129;
    exp_55_ram[923] = 1;
    exp_55_ram[924] = 0;
    exp_55_ram[925] = 1;
    exp_55_ram[926] = 17;
    exp_55_ram[927] = 129;
    exp_55_ram[928] = 1;
    exp_55_ram[929] = 164;
    exp_55_ram[930] = 180;
    exp_55_ram[931] = 196;
    exp_55_ram[932] = 212;
    exp_55_ram[933] = 228;
    exp_55_ram[934] = 244;
    exp_55_ram[935] = 4;
    exp_55_ram[936] = 20;
    exp_55_ram[937] = 68;
    exp_55_ram[938] = 244;
    exp_55_ram[939] = 4;
    exp_55_ram[940] = 39;
    exp_55_ram[941] = 7;
    exp_55_ram[942] = 4;
    exp_55_ram[943] = 23;
    exp_55_ram[944] = 7;
    exp_55_ram[945] = 132;
    exp_55_ram[946] = 244;
    exp_55_ram[947] = 64;
    exp_55_ram[948] = 68;
    exp_55_ram[949] = 23;
    exp_55_ram[950] = 228;
    exp_55_ram[951] = 196;
    exp_55_ram[952] = 4;
    exp_55_ram[953] = 7;
    exp_55_ram[954] = 132;
    exp_55_ram[955] = 0;
    exp_55_ram[956] = 7;
    exp_55_ram[957] = 196;
    exp_55_ram[958] = 23;
    exp_55_ram[959] = 244;
    exp_55_ram[960] = 196;
    exp_55_ram[961] = 68;
    exp_55_ram[962] = 247;
    exp_55_ram[963] = 0;
    exp_55_ram[964] = 132;
    exp_55_ram[965] = 247;
    exp_55_ram[966] = 244;
    exp_55_ram[967] = 196;
    exp_55_ram[968] = 132;
    exp_55_ram[969] = 247;
    exp_55_ram[970] = 7;
    exp_55_ram[971] = 68;
    exp_55_ram[972] = 23;
    exp_55_ram[973] = 228;
    exp_55_ram[974] = 196;
    exp_55_ram[975] = 4;
    exp_55_ram[976] = 7;
    exp_55_ram[977] = 132;
    exp_55_ram[978] = 7;
    exp_55_ram[979] = 132;
    exp_55_ram[980] = 7;
    exp_55_ram[981] = 4;
    exp_55_ram[982] = 39;
    exp_55_ram[983] = 7;
    exp_55_ram[984] = 128;
    exp_55_ram[985] = 68;
    exp_55_ram[986] = 23;
    exp_55_ram[987] = 228;
    exp_55_ram[988] = 196;
    exp_55_ram[989] = 4;
    exp_55_ram[990] = 7;
    exp_55_ram[991] = 132;
    exp_55_ram[992] = 0;
    exp_55_ram[993] = 7;
    exp_55_ram[994] = 68;
    exp_55_ram[995] = 132;
    exp_55_ram[996] = 247;
    exp_55_ram[997] = 68;
    exp_55_ram[998] = 231;
    exp_55_ram[999] = 68;
    exp_55_ram[1000] = 7;
    exp_55_ram[1001] = 193;
    exp_55_ram[1002] = 129;
    exp_55_ram[1003] = 1;
    exp_55_ram[1004] = 0;
    exp_55_ram[1005] = 1;
    exp_55_ram[1006] = 17;
    exp_55_ram[1007] = 129;
    exp_55_ram[1008] = 1;
    exp_55_ram[1009] = 164;
    exp_55_ram[1010] = 180;
    exp_55_ram[1011] = 196;
    exp_55_ram[1012] = 212;
    exp_55_ram[1013] = 228;
    exp_55_ram[1014] = 244;
    exp_55_ram[1015] = 8;
    exp_55_ram[1016] = 20;
    exp_55_ram[1017] = 244;
    exp_55_ram[1018] = 132;
    exp_55_ram[1019] = 39;
    exp_55_ram[1020] = 7;
    exp_55_ram[1021] = 68;
    exp_55_ram[1022] = 7;
    exp_55_ram[1023] = 132;
    exp_55_ram[1024] = 23;
    exp_55_ram[1025] = 7;
    exp_55_ram[1026] = 116;
    exp_55_ram[1027] = 7;
    exp_55_ram[1028] = 132;
    exp_55_ram[1029] = 199;
    exp_55_ram[1030] = 7;
    exp_55_ram[1031] = 68;
    exp_55_ram[1032] = 247;
    exp_55_ram[1033] = 244;
    exp_55_ram[1034] = 0;
    exp_55_ram[1035] = 132;
    exp_55_ram[1036] = 23;
    exp_55_ram[1037] = 228;
    exp_55_ram[1038] = 196;
    exp_55_ram[1039] = 247;
    exp_55_ram[1040] = 0;
    exp_55_ram[1041] = 231;
    exp_55_ram[1042] = 132;
    exp_55_ram[1043] = 4;
    exp_55_ram[1044] = 247;
    exp_55_ram[1045] = 132;
    exp_55_ram[1046] = 240;
    exp_55_ram[1047] = 231;
    exp_55_ram[1048] = 0;
    exp_55_ram[1049] = 132;
    exp_55_ram[1050] = 23;
    exp_55_ram[1051] = 228;
    exp_55_ram[1052] = 196;
    exp_55_ram[1053] = 247;
    exp_55_ram[1054] = 0;
    exp_55_ram[1055] = 231;
    exp_55_ram[1056] = 132;
    exp_55_ram[1057] = 23;
    exp_55_ram[1058] = 7;
    exp_55_ram[1059] = 132;
    exp_55_ram[1060] = 68;
    exp_55_ram[1061] = 247;
    exp_55_ram[1062] = 132;
    exp_55_ram[1063] = 240;
    exp_55_ram[1064] = 231;
    exp_55_ram[1065] = 132;
    exp_55_ram[1066] = 7;
    exp_55_ram[1067] = 7;
    exp_55_ram[1068] = 132;
    exp_55_ram[1069] = 7;
    exp_55_ram[1070] = 7;
    exp_55_ram[1071] = 132;
    exp_55_ram[1072] = 7;
    exp_55_ram[1073] = 132;
    exp_55_ram[1074] = 4;
    exp_55_ram[1075] = 247;
    exp_55_ram[1076] = 132;
    exp_55_ram[1077] = 68;
    exp_55_ram[1078] = 247;
    exp_55_ram[1079] = 132;
    exp_55_ram[1080] = 247;
    exp_55_ram[1081] = 244;
    exp_55_ram[1082] = 132;
    exp_55_ram[1083] = 7;
    exp_55_ram[1084] = 4;
    exp_55_ram[1085] = 0;
    exp_55_ram[1086] = 247;
    exp_55_ram[1087] = 132;
    exp_55_ram[1088] = 247;
    exp_55_ram[1089] = 244;
    exp_55_ram[1090] = 4;
    exp_55_ram[1091] = 0;
    exp_55_ram[1092] = 247;
    exp_55_ram[1093] = 132;
    exp_55_ram[1094] = 7;
    exp_55_ram[1095] = 7;
    exp_55_ram[1096] = 132;
    exp_55_ram[1097] = 240;
    exp_55_ram[1098] = 231;
    exp_55_ram[1099] = 132;
    exp_55_ram[1100] = 23;
    exp_55_ram[1101] = 228;
    exp_55_ram[1102] = 196;
    exp_55_ram[1103] = 247;
    exp_55_ram[1104] = 128;
    exp_55_ram[1105] = 231;
    exp_55_ram[1106] = 192;
    exp_55_ram[1107] = 4;
    exp_55_ram[1108] = 0;
    exp_55_ram[1109] = 247;
    exp_55_ram[1110] = 132;
    exp_55_ram[1111] = 7;
    exp_55_ram[1112] = 7;
    exp_55_ram[1113] = 132;
    exp_55_ram[1114] = 240;
    exp_55_ram[1115] = 231;
    exp_55_ram[1116] = 132;
    exp_55_ram[1117] = 23;
    exp_55_ram[1118] = 228;
    exp_55_ram[1119] = 196;
    exp_55_ram[1120] = 247;
    exp_55_ram[1121] = 128;
    exp_55_ram[1122] = 231;
    exp_55_ram[1123] = 128;
    exp_55_ram[1124] = 4;
    exp_55_ram[1125] = 32;
    exp_55_ram[1126] = 247;
    exp_55_ram[1127] = 132;
    exp_55_ram[1128] = 240;
    exp_55_ram[1129] = 231;
    exp_55_ram[1130] = 132;
    exp_55_ram[1131] = 23;
    exp_55_ram[1132] = 228;
    exp_55_ram[1133] = 196;
    exp_55_ram[1134] = 247;
    exp_55_ram[1135] = 32;
    exp_55_ram[1136] = 231;
    exp_55_ram[1137] = 132;
    exp_55_ram[1138] = 240;
    exp_55_ram[1139] = 231;
    exp_55_ram[1140] = 132;
    exp_55_ram[1141] = 23;
    exp_55_ram[1142] = 228;
    exp_55_ram[1143] = 196;
    exp_55_ram[1144] = 247;
    exp_55_ram[1145] = 0;
    exp_55_ram[1146] = 231;
    exp_55_ram[1147] = 132;
    exp_55_ram[1148] = 240;
    exp_55_ram[1149] = 231;
    exp_55_ram[1150] = 116;
    exp_55_ram[1151] = 7;
    exp_55_ram[1152] = 132;
    exp_55_ram[1153] = 23;
    exp_55_ram[1154] = 228;
    exp_55_ram[1155] = 196;
    exp_55_ram[1156] = 247;
    exp_55_ram[1157] = 208;
    exp_55_ram[1158] = 231;
    exp_55_ram[1159] = 128;
    exp_55_ram[1160] = 132;
    exp_55_ram[1161] = 71;
    exp_55_ram[1162] = 7;
    exp_55_ram[1163] = 132;
    exp_55_ram[1164] = 23;
    exp_55_ram[1165] = 228;
    exp_55_ram[1166] = 196;
    exp_55_ram[1167] = 247;
    exp_55_ram[1168] = 176;
    exp_55_ram[1169] = 231;
    exp_55_ram[1170] = 192;
    exp_55_ram[1171] = 132;
    exp_55_ram[1172] = 135;
    exp_55_ram[1173] = 7;
    exp_55_ram[1174] = 132;
    exp_55_ram[1175] = 23;
    exp_55_ram[1176] = 228;
    exp_55_ram[1177] = 196;
    exp_55_ram[1178] = 247;
    exp_55_ram[1179] = 0;
    exp_55_ram[1180] = 231;
    exp_55_ram[1181] = 132;
    exp_55_ram[1182] = 68;
    exp_55_ram[1183] = 132;
    exp_55_ram[1184] = 196;
    exp_55_ram[1185] = 4;
    exp_55_ram[1186] = 68;
    exp_55_ram[1187] = 132;
    exp_55_ram[1188] = 196;
    exp_55_ram[1189] = 31;
    exp_55_ram[1190] = 5;
    exp_55_ram[1191] = 7;
    exp_55_ram[1192] = 193;
    exp_55_ram[1193] = 129;
    exp_55_ram[1194] = 1;
    exp_55_ram[1195] = 0;
    exp_55_ram[1196] = 1;
    exp_55_ram[1197] = 17;
    exp_55_ram[1198] = 129;
    exp_55_ram[1199] = 1;
    exp_55_ram[1200] = 164;
    exp_55_ram[1201] = 180;
    exp_55_ram[1202] = 196;
    exp_55_ram[1203] = 212;
    exp_55_ram[1204] = 228;
    exp_55_ram[1205] = 4;
    exp_55_ram[1206] = 20;
    exp_55_ram[1207] = 244;
    exp_55_ram[1208] = 4;
    exp_55_ram[1209] = 196;
    exp_55_ram[1210] = 7;
    exp_55_ram[1211] = 68;
    exp_55_ram[1212] = 247;
    exp_55_ram[1213] = 244;
    exp_55_ram[1214] = 68;
    exp_55_ram[1215] = 7;
    exp_55_ram[1216] = 7;
    exp_55_ram[1217] = 196;
    exp_55_ram[1218] = 7;
    exp_55_ram[1219] = 196;
    exp_55_ram[1220] = 68;
    exp_55_ram[1221] = 247;
    exp_55_ram[1222] = 244;
    exp_55_ram[1223] = 180;
    exp_55_ram[1224] = 144;
    exp_55_ram[1225] = 231;
    exp_55_ram[1226] = 180;
    exp_55_ram[1227] = 7;
    exp_55_ram[1228] = 247;
    exp_55_ram[1229] = 0;
    exp_55_ram[1230] = 68;
    exp_55_ram[1231] = 7;
    exp_55_ram[1232] = 7;
    exp_55_ram[1233] = 16;
    exp_55_ram[1234] = 128;
    exp_55_ram[1235] = 16;
    exp_55_ram[1236] = 180;
    exp_55_ram[1237] = 231;
    exp_55_ram[1238] = 247;
    exp_55_ram[1239] = 103;
    exp_55_ram[1240] = 247;
    exp_55_ram[1241] = 196;
    exp_55_ram[1242] = 23;
    exp_55_ram[1243] = 212;
    exp_55_ram[1244] = 4;
    exp_55_ram[1245] = 230;
    exp_55_ram[1246] = 247;
    exp_55_ram[1247] = 196;
    exp_55_ram[1248] = 68;
    exp_55_ram[1249] = 247;
    exp_55_ram[1250] = 244;
    exp_55_ram[1251] = 196;
    exp_55_ram[1252] = 7;
    exp_55_ram[1253] = 196;
    exp_55_ram[1254] = 240;
    exp_55_ram[1255] = 231;
    exp_55_ram[1256] = 180;
    exp_55_ram[1257] = 132;
    exp_55_ram[1258] = 68;
    exp_55_ram[1259] = 241;
    exp_55_ram[1260] = 4;
    exp_55_ram[1261] = 241;
    exp_55_ram[1262] = 4;
    exp_55_ram[1263] = 241;
    exp_55_ram[1264] = 68;
    exp_55_ram[1265] = 6;
    exp_55_ram[1266] = 196;
    exp_55_ram[1267] = 4;
    exp_55_ram[1268] = 68;
    exp_55_ram[1269] = 132;
    exp_55_ram[1270] = 196;
    exp_55_ram[1271] = 159;
    exp_55_ram[1272] = 5;
    exp_55_ram[1273] = 7;
    exp_55_ram[1274] = 193;
    exp_55_ram[1275] = 129;
    exp_55_ram[1276] = 1;
    exp_55_ram[1277] = 0;
    exp_55_ram[1278] = 1;
    exp_55_ram[1279] = 17;
    exp_55_ram[1280] = 129;
    exp_55_ram[1281] = 1;
    exp_55_ram[1282] = 164;
    exp_55_ram[1283] = 180;
    exp_55_ram[1284] = 196;
    exp_55_ram[1285] = 212;
    exp_55_ram[1286] = 228;
    exp_55_ram[1287] = 4;
    exp_55_ram[1288] = 132;
    exp_55_ram[1289] = 7;
    exp_55_ram[1290] = 0;
    exp_55_ram[1291] = 135;
    exp_55_ram[1292] = 244;
    exp_55_ram[1293] = 208;
    exp_55_ram[1294] = 4;
    exp_55_ram[1295] = 7;
    exp_55_ram[1296] = 80;
    exp_55_ram[1297] = 247;
    exp_55_ram[1298] = 4;
    exp_55_ram[1299] = 7;
    exp_55_ram[1300] = 196;
    exp_55_ram[1301] = 23;
    exp_55_ram[1302] = 228;
    exp_55_ram[1303] = 196;
    exp_55_ram[1304] = 68;
    exp_55_ram[1305] = 7;
    exp_55_ram[1306] = 132;
    exp_55_ram[1307] = 7;
    exp_55_ram[1308] = 4;
    exp_55_ram[1309] = 23;
    exp_55_ram[1310] = 244;
    exp_55_ram[1311] = 80;
    exp_55_ram[1312] = 4;
    exp_55_ram[1313] = 23;
    exp_55_ram[1314] = 244;
    exp_55_ram[1315] = 4;
    exp_55_ram[1316] = 4;
    exp_55_ram[1317] = 7;
    exp_55_ram[1318] = 7;
    exp_55_ram[1319] = 0;
    exp_55_ram[1320] = 247;
    exp_55_ram[1321] = 39;
    exp_55_ram[1322] = 0;
    exp_55_ram[1323] = 7;
    exp_55_ram[1324] = 247;
    exp_55_ram[1325] = 7;
    exp_55_ram[1326] = 7;
    exp_55_ram[1327] = 196;
    exp_55_ram[1328] = 23;
    exp_55_ram[1329] = 244;
    exp_55_ram[1330] = 4;
    exp_55_ram[1331] = 23;
    exp_55_ram[1332] = 244;
    exp_55_ram[1333] = 16;
    exp_55_ram[1334] = 244;
    exp_55_ram[1335] = 192;
    exp_55_ram[1336] = 196;
    exp_55_ram[1337] = 39;
    exp_55_ram[1338] = 244;
    exp_55_ram[1339] = 4;
    exp_55_ram[1340] = 23;
    exp_55_ram[1341] = 244;
    exp_55_ram[1342] = 16;
    exp_55_ram[1343] = 244;
    exp_55_ram[1344] = 128;
    exp_55_ram[1345] = 196;
    exp_55_ram[1346] = 71;
    exp_55_ram[1347] = 244;
    exp_55_ram[1348] = 4;
    exp_55_ram[1349] = 23;
    exp_55_ram[1350] = 244;
    exp_55_ram[1351] = 16;
    exp_55_ram[1352] = 244;
    exp_55_ram[1353] = 64;
    exp_55_ram[1354] = 196;
    exp_55_ram[1355] = 135;
    exp_55_ram[1356] = 244;
    exp_55_ram[1357] = 4;
    exp_55_ram[1358] = 23;
    exp_55_ram[1359] = 244;
    exp_55_ram[1360] = 16;
    exp_55_ram[1361] = 244;
    exp_55_ram[1362] = 0;
    exp_55_ram[1363] = 196;
    exp_55_ram[1364] = 7;
    exp_55_ram[1365] = 244;
    exp_55_ram[1366] = 4;
    exp_55_ram[1367] = 23;
    exp_55_ram[1368] = 244;
    exp_55_ram[1369] = 16;
    exp_55_ram[1370] = 244;
    exp_55_ram[1371] = 192;
    exp_55_ram[1372] = 4;
    exp_55_ram[1373] = 0;
    exp_55_ram[1374] = 4;
    exp_55_ram[1375] = 7;
    exp_55_ram[1376] = 4;
    exp_55_ram[1377] = 4;
    exp_55_ram[1378] = 7;
    exp_55_ram[1379] = 7;
    exp_55_ram[1380] = 159;
    exp_55_ram[1381] = 5;
    exp_55_ram[1382] = 7;
    exp_55_ram[1383] = 4;
    exp_55_ram[1384] = 7;
    exp_55_ram[1385] = 95;
    exp_55_ram[1386] = 164;
    exp_55_ram[1387] = 0;
    exp_55_ram[1388] = 4;
    exp_55_ram[1389] = 7;
    exp_55_ram[1390] = 160;
    exp_55_ram[1391] = 247;
    exp_55_ram[1392] = 196;
    exp_55_ram[1393] = 71;
    exp_55_ram[1394] = 228;
    exp_55_ram[1395] = 7;
    exp_55_ram[1396] = 244;
    exp_55_ram[1397] = 132;
    exp_55_ram[1398] = 7;
    exp_55_ram[1399] = 196;
    exp_55_ram[1400] = 39;
    exp_55_ram[1401] = 244;
    exp_55_ram[1402] = 132;
    exp_55_ram[1403] = 240;
    exp_55_ram[1404] = 244;
    exp_55_ram[1405] = 192;
    exp_55_ram[1406] = 132;
    exp_55_ram[1407] = 244;
    exp_55_ram[1408] = 4;
    exp_55_ram[1409] = 23;
    exp_55_ram[1410] = 244;
    exp_55_ram[1411] = 4;
    exp_55_ram[1412] = 4;
    exp_55_ram[1413] = 7;
    exp_55_ram[1414] = 224;
    exp_55_ram[1415] = 247;
    exp_55_ram[1416] = 196;
    exp_55_ram[1417] = 7;
    exp_55_ram[1418] = 244;
    exp_55_ram[1419] = 4;
    exp_55_ram[1420] = 23;
    exp_55_ram[1421] = 244;
    exp_55_ram[1422] = 4;
    exp_55_ram[1423] = 7;
    exp_55_ram[1424] = 7;
    exp_55_ram[1425] = 79;
    exp_55_ram[1426] = 5;
    exp_55_ram[1427] = 7;
    exp_55_ram[1428] = 4;
    exp_55_ram[1429] = 7;
    exp_55_ram[1430] = 15;
    exp_55_ram[1431] = 164;
    exp_55_ram[1432] = 64;
    exp_55_ram[1433] = 4;
    exp_55_ram[1434] = 7;
    exp_55_ram[1435] = 160;
    exp_55_ram[1436] = 247;
    exp_55_ram[1437] = 196;
    exp_55_ram[1438] = 71;
    exp_55_ram[1439] = 228;
    exp_55_ram[1440] = 7;
    exp_55_ram[1441] = 244;
    exp_55_ram[1442] = 68;
    exp_55_ram[1443] = 7;
    exp_55_ram[1444] = 0;
    exp_55_ram[1445] = 244;
    exp_55_ram[1446] = 4;
    exp_55_ram[1447] = 23;
    exp_55_ram[1448] = 244;
    exp_55_ram[1449] = 4;
    exp_55_ram[1450] = 7;
    exp_55_ram[1451] = 135;
    exp_55_ram[1452] = 32;
    exp_55_ram[1453] = 247;
    exp_55_ram[1454] = 39;
    exp_55_ram[1455] = 0;
    exp_55_ram[1456] = 71;
    exp_55_ram[1457] = 247;
    exp_55_ram[1458] = 7;
    exp_55_ram[1459] = 7;
    exp_55_ram[1460] = 196;
    exp_55_ram[1461] = 7;
    exp_55_ram[1462] = 244;
    exp_55_ram[1463] = 4;
    exp_55_ram[1464] = 23;
    exp_55_ram[1465] = 244;
    exp_55_ram[1466] = 4;
    exp_55_ram[1467] = 7;
    exp_55_ram[1468] = 192;
    exp_55_ram[1469] = 247;
    exp_55_ram[1470] = 196;
    exp_55_ram[1471] = 7;
    exp_55_ram[1472] = 244;
    exp_55_ram[1473] = 4;
    exp_55_ram[1474] = 23;
    exp_55_ram[1475] = 244;
    exp_55_ram[1476] = 64;
    exp_55_ram[1477] = 196;
    exp_55_ram[1478] = 7;
    exp_55_ram[1479] = 244;
    exp_55_ram[1480] = 4;
    exp_55_ram[1481] = 23;
    exp_55_ram[1482] = 244;
    exp_55_ram[1483] = 4;
    exp_55_ram[1484] = 7;
    exp_55_ram[1485] = 128;
    exp_55_ram[1486] = 247;
    exp_55_ram[1487] = 196;
    exp_55_ram[1488] = 7;
    exp_55_ram[1489] = 244;
    exp_55_ram[1490] = 4;
    exp_55_ram[1491] = 23;
    exp_55_ram[1492] = 244;
    exp_55_ram[1493] = 128;
    exp_55_ram[1494] = 196;
    exp_55_ram[1495] = 7;
    exp_55_ram[1496] = 244;
    exp_55_ram[1497] = 4;
    exp_55_ram[1498] = 23;
    exp_55_ram[1499] = 244;
    exp_55_ram[1500] = 0;
    exp_55_ram[1501] = 196;
    exp_55_ram[1502] = 7;
    exp_55_ram[1503] = 244;
    exp_55_ram[1504] = 4;
    exp_55_ram[1505] = 23;
    exp_55_ram[1506] = 244;
    exp_55_ram[1507] = 64;
    exp_55_ram[1508] = 196;
    exp_55_ram[1509] = 7;
    exp_55_ram[1510] = 244;
    exp_55_ram[1511] = 4;
    exp_55_ram[1512] = 23;
    exp_55_ram[1513] = 244;
    exp_55_ram[1514] = 128;
    exp_55_ram[1515] = 0;
    exp_55_ram[1516] = 0;
    exp_55_ram[1517] = 0;
    exp_55_ram[1518] = 128;
    exp_55_ram[1519] = 0;
    exp_55_ram[1520] = 4;
    exp_55_ram[1521] = 7;
    exp_55_ram[1522] = 183;
    exp_55_ram[1523] = 48;
    exp_55_ram[1524] = 247;
    exp_55_ram[1525] = 39;
    exp_55_ram[1526] = 0;
    exp_55_ram[1527] = 7;
    exp_55_ram[1528] = 247;
    exp_55_ram[1529] = 7;
    exp_55_ram[1530] = 7;
    exp_55_ram[1531] = 4;
    exp_55_ram[1532] = 7;
    exp_55_ram[1533] = 128;
    exp_55_ram[1534] = 247;
    exp_55_ram[1535] = 4;
    exp_55_ram[1536] = 7;
    exp_55_ram[1537] = 128;
    exp_55_ram[1538] = 247;
    exp_55_ram[1539] = 0;
    exp_55_ram[1540] = 244;
    exp_55_ram[1541] = 0;
    exp_55_ram[1542] = 4;
    exp_55_ram[1543] = 7;
    exp_55_ram[1544] = 240;
    exp_55_ram[1545] = 247;
    exp_55_ram[1546] = 128;
    exp_55_ram[1547] = 244;
    exp_55_ram[1548] = 64;
    exp_55_ram[1549] = 4;
    exp_55_ram[1550] = 7;
    exp_55_ram[1551] = 32;
    exp_55_ram[1552] = 247;
    exp_55_ram[1553] = 32;
    exp_55_ram[1554] = 244;
    exp_55_ram[1555] = 128;
    exp_55_ram[1556] = 160;
    exp_55_ram[1557] = 244;
    exp_55_ram[1558] = 196;
    exp_55_ram[1559] = 247;
    exp_55_ram[1560] = 244;
    exp_55_ram[1561] = 4;
    exp_55_ram[1562] = 7;
    exp_55_ram[1563] = 128;
    exp_55_ram[1564] = 247;
    exp_55_ram[1565] = 196;
    exp_55_ram[1566] = 7;
    exp_55_ram[1567] = 244;
    exp_55_ram[1568] = 4;
    exp_55_ram[1569] = 7;
    exp_55_ram[1570] = 144;
    exp_55_ram[1571] = 247;
    exp_55_ram[1572] = 4;
    exp_55_ram[1573] = 7;
    exp_55_ram[1574] = 64;
    exp_55_ram[1575] = 247;
    exp_55_ram[1576] = 196;
    exp_55_ram[1577] = 55;
    exp_55_ram[1578] = 244;
    exp_55_ram[1579] = 196;
    exp_55_ram[1580] = 7;
    exp_55_ram[1581] = 7;
    exp_55_ram[1582] = 196;
    exp_55_ram[1583] = 231;
    exp_55_ram[1584] = 244;
    exp_55_ram[1585] = 4;
    exp_55_ram[1586] = 7;
    exp_55_ram[1587] = 144;
    exp_55_ram[1588] = 247;
    exp_55_ram[1589] = 4;
    exp_55_ram[1590] = 7;
    exp_55_ram[1591] = 64;
    exp_55_ram[1592] = 247;
    exp_55_ram[1593] = 196;
    exp_55_ram[1594] = 7;
    exp_55_ram[1595] = 7;
    exp_55_ram[1596] = 196;
    exp_55_ram[1597] = 7;
    exp_55_ram[1598] = 7;
    exp_55_ram[1599] = 196;
    exp_55_ram[1600] = 71;
    exp_55_ram[1601] = 228;
    exp_55_ram[1602] = 7;
    exp_55_ram[1603] = 244;
    exp_55_ram[1604] = 132;
    exp_55_ram[1605] = 247;
    exp_55_ram[1606] = 132;
    exp_55_ram[1607] = 247;
    exp_55_ram[1608] = 231;
    exp_55_ram[1609] = 7;
    exp_55_ram[1610] = 132;
    exp_55_ram[1611] = 247;
    exp_55_ram[1612] = 247;
    exp_55_ram[1613] = 196;
    exp_55_ram[1614] = 241;
    exp_55_ram[1615] = 132;
    exp_55_ram[1616] = 241;
    exp_55_ram[1617] = 68;
    exp_55_ram[1618] = 132;
    exp_55_ram[1619] = 7;
    exp_55_ram[1620] = 6;
    exp_55_ram[1621] = 68;
    exp_55_ram[1622] = 196;
    exp_55_ram[1623] = 132;
    exp_55_ram[1624] = 196;
    exp_55_ram[1625] = 223;
    exp_55_ram[1626] = 164;
    exp_55_ram[1627] = 192;
    exp_55_ram[1628] = 196;
    exp_55_ram[1629] = 7;
    exp_55_ram[1630] = 7;
    exp_55_ram[1631] = 196;
    exp_55_ram[1632] = 71;
    exp_55_ram[1633] = 228;
    exp_55_ram[1634] = 7;
    exp_55_ram[1635] = 247;
    exp_55_ram[1636] = 192;
    exp_55_ram[1637] = 196;
    exp_55_ram[1638] = 7;
    exp_55_ram[1639] = 7;
    exp_55_ram[1640] = 196;
    exp_55_ram[1641] = 71;
    exp_55_ram[1642] = 228;
    exp_55_ram[1643] = 7;
    exp_55_ram[1644] = 7;
    exp_55_ram[1645] = 7;
    exp_55_ram[1646] = 64;
    exp_55_ram[1647] = 196;
    exp_55_ram[1648] = 71;
    exp_55_ram[1649] = 228;
    exp_55_ram[1650] = 7;
    exp_55_ram[1651] = 244;
    exp_55_ram[1652] = 196;
    exp_55_ram[1653] = 247;
    exp_55_ram[1654] = 196;
    exp_55_ram[1655] = 247;
    exp_55_ram[1656] = 231;
    exp_55_ram[1657] = 7;
    exp_55_ram[1658] = 196;
    exp_55_ram[1659] = 247;
    exp_55_ram[1660] = 247;
    exp_55_ram[1661] = 196;
    exp_55_ram[1662] = 241;
    exp_55_ram[1663] = 132;
    exp_55_ram[1664] = 241;
    exp_55_ram[1665] = 68;
    exp_55_ram[1666] = 132;
    exp_55_ram[1667] = 7;
    exp_55_ram[1668] = 6;
    exp_55_ram[1669] = 68;
    exp_55_ram[1670] = 196;
    exp_55_ram[1671] = 132;
    exp_55_ram[1672] = 196;
    exp_55_ram[1673] = 223;
    exp_55_ram[1674] = 164;
    exp_55_ram[1675] = 192;
    exp_55_ram[1676] = 196;
    exp_55_ram[1677] = 7;
    exp_55_ram[1678] = 7;
    exp_55_ram[1679] = 196;
    exp_55_ram[1680] = 7;
    exp_55_ram[1681] = 7;
    exp_55_ram[1682] = 196;
    exp_55_ram[1683] = 71;
    exp_55_ram[1684] = 228;
    exp_55_ram[1685] = 7;
    exp_55_ram[1686] = 196;
    exp_55_ram[1687] = 241;
    exp_55_ram[1688] = 132;
    exp_55_ram[1689] = 241;
    exp_55_ram[1690] = 68;
    exp_55_ram[1691] = 132;
    exp_55_ram[1692] = 0;
    exp_55_ram[1693] = 68;
    exp_55_ram[1694] = 196;
    exp_55_ram[1695] = 132;
    exp_55_ram[1696] = 196;
    exp_55_ram[1697] = 223;
    exp_55_ram[1698] = 164;
    exp_55_ram[1699] = 192;
    exp_55_ram[1700] = 196;
    exp_55_ram[1701] = 7;
    exp_55_ram[1702] = 7;
    exp_55_ram[1703] = 196;
    exp_55_ram[1704] = 71;
    exp_55_ram[1705] = 228;
    exp_55_ram[1706] = 7;
    exp_55_ram[1707] = 247;
    exp_55_ram[1708] = 192;
    exp_55_ram[1709] = 196;
    exp_55_ram[1710] = 7;
    exp_55_ram[1711] = 7;
    exp_55_ram[1712] = 196;
    exp_55_ram[1713] = 71;
    exp_55_ram[1714] = 228;
    exp_55_ram[1715] = 7;
    exp_55_ram[1716] = 7;
    exp_55_ram[1717] = 7;
    exp_55_ram[1718] = 64;
    exp_55_ram[1719] = 196;
    exp_55_ram[1720] = 71;
    exp_55_ram[1721] = 228;
    exp_55_ram[1722] = 7;
    exp_55_ram[1723] = 244;
    exp_55_ram[1724] = 196;
    exp_55_ram[1725] = 241;
    exp_55_ram[1726] = 132;
    exp_55_ram[1727] = 241;
    exp_55_ram[1728] = 68;
    exp_55_ram[1729] = 132;
    exp_55_ram[1730] = 0;
    exp_55_ram[1731] = 4;
    exp_55_ram[1732] = 68;
    exp_55_ram[1733] = 196;
    exp_55_ram[1734] = 132;
    exp_55_ram[1735] = 196;
    exp_55_ram[1736] = 15;
    exp_55_ram[1737] = 164;
    exp_55_ram[1738] = 4;
    exp_55_ram[1739] = 23;
    exp_55_ram[1740] = 244;
    exp_55_ram[1741] = 192;
    exp_55_ram[1742] = 16;
    exp_55_ram[1743] = 244;
    exp_55_ram[1744] = 196;
    exp_55_ram[1745] = 39;
    exp_55_ram[1746] = 7;
    exp_55_ram[1747] = 128;
    exp_55_ram[1748] = 196;
    exp_55_ram[1749] = 23;
    exp_55_ram[1750] = 228;
    exp_55_ram[1751] = 196;
    exp_55_ram[1752] = 68;
    exp_55_ram[1753] = 7;
    exp_55_ram[1754] = 132;
    exp_55_ram[1755] = 0;
    exp_55_ram[1756] = 7;
    exp_55_ram[1757] = 68;
    exp_55_ram[1758] = 23;
    exp_55_ram[1759] = 228;
    exp_55_ram[1760] = 132;
    exp_55_ram[1761] = 231;
    exp_55_ram[1762] = 196;
    exp_55_ram[1763] = 71;
    exp_55_ram[1764] = 228;
    exp_55_ram[1765] = 7;
    exp_55_ram[1766] = 247;
    exp_55_ram[1767] = 196;
    exp_55_ram[1768] = 23;
    exp_55_ram[1769] = 228;
    exp_55_ram[1770] = 196;
    exp_55_ram[1771] = 68;
    exp_55_ram[1772] = 7;
    exp_55_ram[1773] = 132;
    exp_55_ram[1774] = 7;
    exp_55_ram[1775] = 196;
    exp_55_ram[1776] = 39;
    exp_55_ram[1777] = 7;
    exp_55_ram[1778] = 128;
    exp_55_ram[1779] = 196;
    exp_55_ram[1780] = 23;
    exp_55_ram[1781] = 228;
    exp_55_ram[1782] = 196;
    exp_55_ram[1783] = 68;
    exp_55_ram[1784] = 7;
    exp_55_ram[1785] = 132;
    exp_55_ram[1786] = 0;
    exp_55_ram[1787] = 7;
    exp_55_ram[1788] = 68;
    exp_55_ram[1789] = 23;
    exp_55_ram[1790] = 228;
    exp_55_ram[1791] = 132;
    exp_55_ram[1792] = 231;
    exp_55_ram[1793] = 4;
    exp_55_ram[1794] = 23;
    exp_55_ram[1795] = 244;
    exp_55_ram[1796] = 0;
    exp_55_ram[1797] = 196;
    exp_55_ram[1798] = 71;
    exp_55_ram[1799] = 228;
    exp_55_ram[1800] = 7;
    exp_55_ram[1801] = 244;
    exp_55_ram[1802] = 68;
    exp_55_ram[1803] = 7;
    exp_55_ram[1804] = 68;
    exp_55_ram[1805] = 128;
    exp_55_ram[1806] = 240;
    exp_55_ram[1807] = 7;
    exp_55_ram[1808] = 4;
    exp_55_ram[1809] = 15;
    exp_55_ram[1810] = 164;
    exp_55_ram[1811] = 196;
    exp_55_ram[1812] = 7;
    exp_55_ram[1813] = 7;
    exp_55_ram[1814] = 196;
    exp_55_ram[1815] = 68;
    exp_55_ram[1816] = 247;
    exp_55_ram[1817] = 7;
    exp_55_ram[1818] = 244;
    exp_55_ram[1819] = 196;
    exp_55_ram[1820] = 39;
    exp_55_ram[1821] = 7;
    exp_55_ram[1822] = 128;
    exp_55_ram[1823] = 196;
    exp_55_ram[1824] = 23;
    exp_55_ram[1825] = 228;
    exp_55_ram[1826] = 196;
    exp_55_ram[1827] = 68;
    exp_55_ram[1828] = 7;
    exp_55_ram[1829] = 132;
    exp_55_ram[1830] = 0;
    exp_55_ram[1831] = 7;
    exp_55_ram[1832] = 196;
    exp_55_ram[1833] = 23;
    exp_55_ram[1834] = 228;
    exp_55_ram[1835] = 132;
    exp_55_ram[1836] = 231;
    exp_55_ram[1837] = 64;
    exp_55_ram[1838] = 4;
    exp_55_ram[1839] = 23;
    exp_55_ram[1840] = 228;
    exp_55_ram[1841] = 7;
    exp_55_ram[1842] = 196;
    exp_55_ram[1843] = 23;
    exp_55_ram[1844] = 228;
    exp_55_ram[1845] = 196;
    exp_55_ram[1846] = 68;
    exp_55_ram[1847] = 7;
    exp_55_ram[1848] = 132;
    exp_55_ram[1849] = 7;
    exp_55_ram[1850] = 4;
    exp_55_ram[1851] = 7;
    exp_55_ram[1852] = 7;
    exp_55_ram[1853] = 196;
    exp_55_ram[1854] = 7;
    exp_55_ram[1855] = 7;
    exp_55_ram[1856] = 68;
    exp_55_ram[1857] = 247;
    exp_55_ram[1858] = 228;
    exp_55_ram[1859] = 7;
    exp_55_ram[1860] = 196;
    exp_55_ram[1861] = 39;
    exp_55_ram[1862] = 7;
    exp_55_ram[1863] = 128;
    exp_55_ram[1864] = 196;
    exp_55_ram[1865] = 23;
    exp_55_ram[1866] = 228;
    exp_55_ram[1867] = 196;
    exp_55_ram[1868] = 68;
    exp_55_ram[1869] = 7;
    exp_55_ram[1870] = 132;
    exp_55_ram[1871] = 0;
    exp_55_ram[1872] = 7;
    exp_55_ram[1873] = 196;
    exp_55_ram[1874] = 23;
    exp_55_ram[1875] = 228;
    exp_55_ram[1876] = 132;
    exp_55_ram[1877] = 231;
    exp_55_ram[1878] = 4;
    exp_55_ram[1879] = 23;
    exp_55_ram[1880] = 244;
    exp_55_ram[1881] = 192;
    exp_55_ram[1882] = 128;
    exp_55_ram[1883] = 244;
    exp_55_ram[1884] = 196;
    exp_55_ram[1885] = 23;
    exp_55_ram[1886] = 244;
    exp_55_ram[1887] = 196;
    exp_55_ram[1888] = 71;
    exp_55_ram[1889] = 228;
    exp_55_ram[1890] = 7;
    exp_55_ram[1891] = 7;
    exp_55_ram[1892] = 196;
    exp_55_ram[1893] = 241;
    exp_55_ram[1894] = 132;
    exp_55_ram[1895] = 241;
    exp_55_ram[1896] = 68;
    exp_55_ram[1897] = 0;
    exp_55_ram[1898] = 0;
    exp_55_ram[1899] = 68;
    exp_55_ram[1900] = 196;
    exp_55_ram[1901] = 132;
    exp_55_ram[1902] = 196;
    exp_55_ram[1903] = 79;
    exp_55_ram[1904] = 164;
    exp_55_ram[1905] = 4;
    exp_55_ram[1906] = 23;
    exp_55_ram[1907] = 244;
    exp_55_ram[1908] = 0;
    exp_55_ram[1909] = 196;
    exp_55_ram[1910] = 23;
    exp_55_ram[1911] = 228;
    exp_55_ram[1912] = 196;
    exp_55_ram[1913] = 68;
    exp_55_ram[1914] = 7;
    exp_55_ram[1915] = 132;
    exp_55_ram[1916] = 80;
    exp_55_ram[1917] = 7;
    exp_55_ram[1918] = 4;
    exp_55_ram[1919] = 23;
    exp_55_ram[1920] = 244;
    exp_55_ram[1921] = 192;
    exp_55_ram[1922] = 4;
    exp_55_ram[1923] = 7;
    exp_55_ram[1924] = 196;
    exp_55_ram[1925] = 23;
    exp_55_ram[1926] = 228;
    exp_55_ram[1927] = 196;
    exp_55_ram[1928] = 68;
    exp_55_ram[1929] = 7;
    exp_55_ram[1930] = 132;
    exp_55_ram[1931] = 7;
    exp_55_ram[1932] = 4;
    exp_55_ram[1933] = 23;
    exp_55_ram[1934] = 244;
    exp_55_ram[1935] = 0;
    exp_55_ram[1936] = 4;
    exp_55_ram[1937] = 7;
    exp_55_ram[1938] = 7;
    exp_55_ram[1939] = 196;
    exp_55_ram[1940] = 68;
    exp_55_ram[1941] = 247;
    exp_55_ram[1942] = 68;
    exp_55_ram[1943] = 247;
    exp_55_ram[1944] = 128;
    exp_55_ram[1945] = 196;
    exp_55_ram[1946] = 196;
    exp_55_ram[1947] = 68;
    exp_55_ram[1948] = 7;
    exp_55_ram[1949] = 132;
    exp_55_ram[1950] = 0;
    exp_55_ram[1951] = 7;
    exp_55_ram[1952] = 196;
    exp_55_ram[1953] = 7;
    exp_55_ram[1954] = 193;
    exp_55_ram[1955] = 129;
    exp_55_ram[1956] = 1;
    exp_55_ram[1957] = 0;
    exp_55_ram[1958] = 1;
    exp_55_ram[1959] = 17;
    exp_55_ram[1960] = 129;
    exp_55_ram[1961] = 1;
    exp_55_ram[1962] = 164;
    exp_55_ram[1963] = 180;
    exp_55_ram[1964] = 196;
    exp_55_ram[1965] = 212;
    exp_55_ram[1966] = 228;
    exp_55_ram[1967] = 244;
    exp_55_ram[1968] = 4;
    exp_55_ram[1969] = 20;
    exp_55_ram[1970] = 4;
    exp_55_ram[1971] = 244;
    exp_55_ram[1972] = 132;
    exp_55_ram[1973] = 71;
    exp_55_ram[1974] = 244;
    exp_55_ram[1975] = 132;
    exp_55_ram[1976] = 68;
    exp_55_ram[1977] = 196;
    exp_55_ram[1978] = 240;
    exp_55_ram[1979] = 7;
    exp_55_ram[1980] = 0;
    exp_55_ram[1981] = 135;
    exp_55_ram[1982] = 15;
    exp_55_ram[1983] = 164;
    exp_55_ram[1984] = 196;
    exp_55_ram[1985] = 7;
    exp_55_ram[1986] = 193;
    exp_55_ram[1987] = 129;
    exp_55_ram[1988] = 1;
    exp_55_ram[1989] = 0;
    exp_55_ram[1990] = 1;
    exp_55_ram[1991] = 17;
    exp_55_ram[1992] = 129;
    exp_55_ram[1993] = 1;
    exp_55_ram[1994] = 5;
    exp_55_ram[1995] = 244;
    exp_55_ram[1996] = 244;
    exp_55_ram[1997] = 0;
    exp_55_ram[1998] = 135;
    exp_55_ram[1999] = 7;
    exp_55_ram[2000] = 7;
    exp_55_ram[2001] = 223;
    exp_55_ram[2002] = 0;
    exp_55_ram[2003] = 193;
    exp_55_ram[2004] = 129;
    exp_55_ram[2005] = 1;
    exp_55_ram[2006] = 0;
    exp_55_ram[2007] = 1;
    exp_55_ram[2008] = 17;
    exp_55_ram[2009] = 129;
    exp_55_ram[2010] = 145;
    exp_55_ram[2011] = 1;
    exp_55_ram[2012] = 5;
    exp_55_ram[2013] = 68;
    exp_55_ram[2014] = 244;
    exp_55_ram[2015] = 144;
    exp_55_ram[2016] = 244;
    exp_55_ram[2017] = 240;
    exp_55_ram[2018] = 244;
    exp_55_ram[2019] = 16;
    exp_55_ram[2020] = 244;
    exp_55_ram[2021] = 4;
    exp_55_ram[2022] = 4;
    exp_55_ram[2023] = 4;
    exp_55_ram[2024] = 68;
    exp_55_ram[2025] = 132;
    exp_55_ram[2026] = 196;
    exp_55_ram[2027] = 4;
    exp_55_ram[2028] = 68;
    exp_55_ram[2029] = 132;
    exp_55_ram[2030] = 196;
    exp_55_ram[2031] = 4;
    exp_55_ram[2032] = 68;
    exp_55_ram[2033] = 100;
    exp_55_ram[2034] = 20;
    exp_55_ram[2035] = 4;
    exp_55_ram[2036] = 164;
    exp_55_ram[2037] = 180;
    exp_55_ram[2038] = 196;
    exp_55_ram[2039] = 212;
    exp_55_ram[2040] = 228;
    exp_55_ram[2041] = 244;
    exp_55_ram[2042] = 4;
    exp_55_ram[2043] = 7;
    exp_55_ram[2044] = 64;
    exp_55_ram[2045] = 164;
    exp_55_ram[2046] = 180;
    exp_55_ram[2047] = 68;
    exp_55_ram[2048] = 132;
    exp_55_ram[2049] = 196;
    exp_55_ram[2050] = 7;
    exp_55_ram[2051] = 0;
    exp_55_ram[2052] = 4;
    exp_55_ram[2053] = 196;
    exp_55_ram[2054] = 247;
    exp_55_ram[2055] = 244;
    exp_55_ram[2056] = 68;
    exp_55_ram[2057] = 132;
    exp_55_ram[2058] = 196;
    exp_55_ram[2059] = 4;
    exp_55_ram[2060] = 68;
    exp_55_ram[2061] = 132;
    exp_55_ram[2062] = 196;
    exp_55_ram[2063] = 4;
    exp_55_ram[2064] = 68;
    exp_55_ram[2065] = 100;
    exp_55_ram[2066] = 20;
    exp_55_ram[2067] = 4;
    exp_55_ram[2068] = 164;
    exp_55_ram[2069] = 180;
    exp_55_ram[2070] = 196;
    exp_55_ram[2071] = 212;
    exp_55_ram[2072] = 228;
    exp_55_ram[2073] = 244;
    exp_55_ram[2074] = 4;
    exp_55_ram[2075] = 7;
    exp_55_ram[2076] = 64;
    exp_55_ram[2077] = 164;
    exp_55_ram[2078] = 180;
    exp_55_ram[2079] = 68;
    exp_55_ram[2080] = 244;
    exp_55_ram[2081] = 32;
    exp_55_ram[2082] = 244;
    exp_55_ram[2083] = 240;
    exp_55_ram[2084] = 244;
    exp_55_ram[2085] = 16;
    exp_55_ram[2086] = 244;
    exp_55_ram[2087] = 4;
    exp_55_ram[2088] = 4;
    exp_55_ram[2089] = 4;
    exp_55_ram[2090] = 4;
    exp_55_ram[2091] = 68;
    exp_55_ram[2092] = 132;
    exp_55_ram[2093] = 196;
    exp_55_ram[2094] = 4;
    exp_55_ram[2095] = 68;
    exp_55_ram[2096] = 132;
    exp_55_ram[2097] = 196;
    exp_55_ram[2098] = 4;
    exp_55_ram[2099] = 100;
    exp_55_ram[2100] = 20;
    exp_55_ram[2101] = 4;
    exp_55_ram[2102] = 164;
    exp_55_ram[2103] = 180;
    exp_55_ram[2104] = 196;
    exp_55_ram[2105] = 212;
    exp_55_ram[2106] = 228;
    exp_55_ram[2107] = 244;
    exp_55_ram[2108] = 4;
    exp_55_ram[2109] = 7;
    exp_55_ram[2110] = 192;
    exp_55_ram[2111] = 164;
    exp_55_ram[2112] = 180;
    exp_55_ram[2113] = 4;
    exp_55_ram[2114] = 4;
    exp_55_ram[2115] = 68;
    exp_55_ram[2116] = 7;
    exp_55_ram[2117] = 144;
    exp_55_ram[2118] = 196;
    exp_55_ram[2119] = 132;
    exp_55_ram[2120] = 247;
    exp_55_ram[2121] = 244;
    exp_55_ram[2122] = 4;
    exp_55_ram[2123] = 68;
    exp_55_ram[2124] = 132;
    exp_55_ram[2125] = 196;
    exp_55_ram[2126] = 4;
    exp_55_ram[2127] = 68;
    exp_55_ram[2128] = 132;
    exp_55_ram[2129] = 196;
    exp_55_ram[2130] = 4;
    exp_55_ram[2131] = 100;
    exp_55_ram[2132] = 20;
    exp_55_ram[2133] = 4;
    exp_55_ram[2134] = 164;
    exp_55_ram[2135] = 180;
    exp_55_ram[2136] = 196;
    exp_55_ram[2137] = 212;
    exp_55_ram[2138] = 228;
    exp_55_ram[2139] = 244;
    exp_55_ram[2140] = 4;
    exp_55_ram[2141] = 7;
    exp_55_ram[2142] = 192;
    exp_55_ram[2143] = 164;
    exp_55_ram[2144] = 180;
    exp_55_ram[2145] = 4;
    exp_55_ram[2146] = 68;
    exp_55_ram[2147] = 132;
    exp_55_ram[2148] = 196;
    exp_55_ram[2149] = 4;
    exp_55_ram[2150] = 68;
    exp_55_ram[2151] = 132;
    exp_55_ram[2152] = 196;
    exp_55_ram[2153] = 4;
    exp_55_ram[2154] = 100;
    exp_55_ram[2155] = 20;
    exp_55_ram[2156] = 4;
    exp_55_ram[2157] = 164;
    exp_55_ram[2158] = 180;
    exp_55_ram[2159] = 196;
    exp_55_ram[2160] = 212;
    exp_55_ram[2161] = 228;
    exp_55_ram[2162] = 244;
    exp_55_ram[2163] = 4;
    exp_55_ram[2164] = 7;
    exp_55_ram[2165] = 0;
    exp_55_ram[2166] = 164;
    exp_55_ram[2167] = 180;
    exp_55_ram[2168] = 68;
    exp_55_ram[2169] = 196;
    exp_55_ram[2170] = 231;
    exp_55_ram[2171] = 68;
    exp_55_ram[2172] = 196;
    exp_55_ram[2173] = 247;
    exp_55_ram[2174] = 4;
    exp_55_ram[2175] = 132;
    exp_55_ram[2176] = 231;
    exp_55_ram[2177] = 196;
    exp_55_ram[2178] = 196;
    exp_55_ram[2179] = 231;
    exp_55_ram[2180] = 196;
    exp_55_ram[2181] = 196;
    exp_55_ram[2182] = 247;
    exp_55_ram[2183] = 132;
    exp_55_ram[2184] = 132;
    exp_55_ram[2185] = 231;
    exp_55_ram[2186] = 16;
    exp_55_ram[2187] = 128;
    exp_55_ram[2188] = 0;
    exp_55_ram[2189] = 7;
    exp_55_ram[2190] = 193;
    exp_55_ram[2191] = 129;
    exp_55_ram[2192] = 65;
    exp_55_ram[2193] = 1;
    exp_55_ram[2194] = 0;
    exp_55_ram[2195] = 1;
    exp_55_ram[2196] = 17;
    exp_55_ram[2197] = 129;
    exp_55_ram[2198] = 1;
    exp_55_ram[2199] = 164;
    exp_55_ram[2200] = 180;
    exp_55_ram[2201] = 196;
    exp_55_ram[2202] = 132;
    exp_55_ram[2203] = 196;
    exp_55_ram[2204] = 7;
    exp_55_ram[2205] = 144;
    exp_55_ram[2206] = 196;
    exp_55_ram[2207] = 4;
    exp_55_ram[2208] = 68;
    exp_55_ram[2209] = 132;
    exp_55_ram[2210] = 196;
    exp_55_ram[2211] = 4;
    exp_55_ram[2212] = 68;
    exp_55_ram[2213] = 132;
    exp_55_ram[2214] = 196;
    exp_55_ram[2215] = 100;
    exp_55_ram[2216] = 20;
    exp_55_ram[2217] = 4;
    exp_55_ram[2218] = 164;
    exp_55_ram[2219] = 180;
    exp_55_ram[2220] = 196;
    exp_55_ram[2221] = 212;
    exp_55_ram[2222] = 228;
    exp_55_ram[2223] = 244;
    exp_55_ram[2224] = 4;
    exp_55_ram[2225] = 7;
    exp_55_ram[2226] = 95;
    exp_55_ram[2227] = 5;
    exp_55_ram[2228] = 7;
    exp_55_ram[2229] = 193;
    exp_55_ram[2230] = 129;
    exp_55_ram[2231] = 1;
    exp_55_ram[2232] = 0;
    exp_55_ram[2233] = 1;
    exp_55_ram[2234] = 129;
    exp_55_ram[2235] = 1;
    exp_55_ram[2236] = 0;
    exp_55_ram[2237] = 212;
    exp_55_ram[2238] = 0;
    exp_55_ram[2239] = 70;
    exp_55_ram[2240] = 212;
    exp_55_ram[2241] = 132;
    exp_55_ram[2242] = 6;
    exp_55_ram[2243] = 212;
    exp_55_ram[2244] = 4;
    exp_55_ram[2245] = 4;
    exp_55_ram[2246] = 6;
    exp_55_ram[2247] = 212;
    exp_55_ram[2248] = 4;
    exp_55_ram[2249] = 196;
    exp_55_ram[2250] = 6;
    exp_55_ram[2251] = 6;
    exp_55_ram[2252] = 0;
    exp_55_ram[2253] = 4;
    exp_55_ram[2254] = 230;
    exp_55_ram[2255] = 212;
    exp_55_ram[2256] = 68;
    exp_55_ram[2257] = 246;
    exp_55_ram[2258] = 244;
    exp_55_ram[2259] = 4;
    exp_55_ram[2260] = 68;
    exp_55_ram[2261] = 7;
    exp_55_ram[2262] = 7;
    exp_55_ram[2263] = 193;
    exp_55_ram[2264] = 1;
    exp_55_ram[2265] = 0;
    exp_55_ram[2266] = 1;
    exp_55_ram[2267] = 17;
    exp_55_ram[2268] = 129;
    exp_55_ram[2269] = 1;
    exp_55_ram[2270] = 164;
    exp_55_ram[2271] = 180;
    exp_55_ram[2272] = 196;
    exp_55_ram[2273] = 212;
    exp_55_ram[2274] = 132;
    exp_55_ram[2275] = 196;
    exp_55_ram[2276] = 4;
    exp_55_ram[2277] = 68;
    exp_55_ram[2278] = 167;
    exp_55_ram[2279] = 6;
    exp_55_ram[2280] = 7;
    exp_55_ram[2281] = 183;
    exp_55_ram[2282] = 6;
    exp_55_ram[2283] = 7;
    exp_55_ram[2284] = 6;
    exp_55_ram[2285] = 6;
    exp_55_ram[2286] = 7;
    exp_55_ram[2287] = 7;
    exp_55_ram[2288] = 79;
    exp_55_ram[2289] = 5;
    exp_55_ram[2290] = 5;
    exp_55_ram[2291] = 7;
    exp_55_ram[2292] = 7;
    exp_55_ram[2293] = 193;
    exp_55_ram[2294] = 129;
    exp_55_ram[2295] = 1;
    exp_55_ram[2296] = 0;
    exp_55_ram[2297] = 1;
    exp_55_ram[2298] = 129;
    exp_55_ram[2299] = 1;
    exp_55_ram[2300] = 164;
    exp_55_ram[2301] = 196;
    exp_55_ram[2302] = 55;
    exp_55_ram[2303] = 7;
    exp_55_ram[2304] = 196;
    exp_55_ram[2305] = 64;
    exp_55_ram[2306] = 247;
    exp_55_ram[2307] = 7;
    exp_55_ram[2308] = 196;
    exp_55_ram[2309] = 0;
    exp_55_ram[2310] = 247;
    exp_55_ram[2311] = 7;
    exp_55_ram[2312] = 16;
    exp_55_ram[2313] = 128;
    exp_55_ram[2314] = 0;
    exp_55_ram[2315] = 7;
    exp_55_ram[2316] = 193;
    exp_55_ram[2317] = 1;
    exp_55_ram[2318] = 0;
    exp_55_ram[2319] = 1;
    exp_55_ram[2320] = 17;
    exp_55_ram[2321] = 129;
    exp_55_ram[2322] = 1;
    exp_55_ram[2323] = 164;
    exp_55_ram[2324] = 196;
    exp_55_ram[2325] = 31;
    exp_55_ram[2326] = 5;
    exp_55_ram[2327] = 7;
    exp_55_ram[2328] = 224;
    exp_55_ram[2329] = 128;
    exp_55_ram[2330] = 208;
    exp_55_ram[2331] = 7;
    exp_55_ram[2332] = 193;
    exp_55_ram[2333] = 129;
    exp_55_ram[2334] = 1;
    exp_55_ram[2335] = 0;
    exp_55_ram[2336] = 1;
    exp_55_ram[2337] = 17;
    exp_55_ram[2338] = 129;
    exp_55_ram[2339] = 1;
    exp_55_ram[2340] = 164;
    exp_55_ram[2341] = 180;
    exp_55_ram[2342] = 132;
    exp_55_ram[2343] = 48;
    exp_55_ram[2344] = 247;
    exp_55_ram[2345] = 132;
    exp_55_ram[2346] = 128;
    exp_55_ram[2347] = 247;
    exp_55_ram[2348] = 132;
    exp_55_ram[2349] = 80;
    exp_55_ram[2350] = 247;
    exp_55_ram[2351] = 132;
    exp_55_ram[2352] = 160;
    exp_55_ram[2353] = 247;
    exp_55_ram[2354] = 224;
    exp_55_ram[2355] = 64;
    exp_55_ram[2356] = 132;
    exp_55_ram[2357] = 16;
    exp_55_ram[2358] = 247;
    exp_55_ram[2359] = 196;
    exp_55_ram[2360] = 95;
    exp_55_ram[2361] = 5;
    exp_55_ram[2362] = 7;
    exp_55_ram[2363] = 208;
    exp_55_ram[2364] = 0;
    exp_55_ram[2365] = 192;
    exp_55_ram[2366] = 128;
    exp_55_ram[2367] = 240;
    exp_55_ram[2368] = 7;
    exp_55_ram[2369] = 193;
    exp_55_ram[2370] = 129;
    exp_55_ram[2371] = 1;
    exp_55_ram[2372] = 0;
    exp_55_ram[2373] = 1;
    exp_55_ram[2374] = 17;
    exp_55_ram[2375] = 129;
    exp_55_ram[2376] = 145;
    exp_55_ram[2377] = 33;
    exp_55_ram[2378] = 49;
    exp_55_ram[2379] = 65;
    exp_55_ram[2380] = 81;
    exp_55_ram[2381] = 97;
    exp_55_ram[2382] = 113;
    exp_55_ram[2383] = 129;
    exp_55_ram[2384] = 145;
    exp_55_ram[2385] = 161;
    exp_55_ram[2386] = 177;
    exp_55_ram[2387] = 1;
    exp_55_ram[2388] = 5;
    exp_55_ram[2389] = 0;
    exp_55_ram[2390] = 0;
    exp_55_ram[2391] = 244;
    exp_55_ram[2392] = 4;
    exp_55_ram[2393] = 32;
    exp_55_ram[2394] = 244;
    exp_55_ram[2395] = 68;
    exp_55_ram[2396] = 244;
    exp_55_ram[2397] = 196;
    exp_55_ram[2398] = 199;
    exp_55_ram[2399] = 68;
    exp_55_ram[2400] = 247;
    exp_55_ram[2401] = 68;
    exp_55_ram[2402] = 95;
    exp_55_ram[2403] = 5;
    exp_55_ram[2404] = 1;
    exp_55_ram[2405] = 7;
    exp_55_ram[2406] = 247;
    exp_55_ram[2407] = 244;
    exp_55_ram[2408] = 4;
    exp_55_ram[2409] = 132;
    exp_55_ram[2410] = 196;
    exp_55_ram[2411] = 132;
    exp_55_ram[2412] = 196;
    exp_55_ram[2413] = 8;
    exp_55_ram[2414] = 182;
    exp_55_ram[2415] = 7;
    exp_55_ram[2416] = 197;
    exp_55_ram[2417] = 8;
    exp_55_ram[2418] = 166;
    exp_55_ram[2419] = 245;
    exp_55_ram[2420] = 6;
    exp_55_ram[2421] = 228;
    exp_55_ram[2422] = 244;
    exp_55_ram[2423] = 68;
    exp_55_ram[2424] = 23;
    exp_55_ram[2425] = 244;
    exp_55_ram[2426] = 223;
    exp_55_ram[2427] = 0;
    exp_55_ram[2428] = 4;
    exp_55_ram[2429] = 4;
    exp_55_ram[2430] = 7;
    exp_55_ram[2431] = 4;
    exp_55_ram[2432] = 231;
    exp_55_ram[2433] = 4;
    exp_55_ram[2434] = 68;
    exp_55_ram[2435] = 95;
    exp_55_ram[2436] = 5;
    exp_55_ram[2437] = 1;
    exp_55_ram[2438] = 7;
    exp_55_ram[2439] = 247;
    exp_55_ram[2440] = 7;
    exp_55_ram[2441] = 0;
    exp_55_ram[2442] = 132;
    exp_55_ram[2443] = 196;
    exp_55_ram[2444] = 166;
    exp_55_ram[2445] = 7;
    exp_55_ram[2446] = 197;
    exp_55_ram[2447] = 182;
    exp_55_ram[2448] = 245;
    exp_55_ram[2449] = 6;
    exp_55_ram[2450] = 228;
    exp_55_ram[2451] = 244;
    exp_55_ram[2452] = 4;
    exp_55_ram[2453] = 23;
    exp_55_ram[2454] = 244;
    exp_55_ram[2455] = 159;
    exp_55_ram[2456] = 0;
    exp_55_ram[2457] = 196;
    exp_55_ram[2458] = 247;
    exp_55_ram[2459] = 1;
    exp_55_ram[2460] = 7;
    exp_55_ram[2461] = 247;
    exp_55_ram[2462] = 7;
    exp_55_ram[2463] = 247;
    exp_55_ram[2464] = 7;
    exp_55_ram[2465] = 132;
    exp_55_ram[2466] = 196;
    exp_55_ram[2467] = 134;
    exp_55_ram[2468] = 7;
    exp_55_ram[2469] = 197;
    exp_55_ram[2470] = 150;
    exp_55_ram[2471] = 245;
    exp_55_ram[2472] = 6;
    exp_55_ram[2473] = 228;
    exp_55_ram[2474] = 244;
    exp_55_ram[2475] = 132;
    exp_55_ram[2476] = 0;
    exp_55_ram[2477] = 7;
    exp_55_ram[2478] = 247;
    exp_55_ram[2479] = 7;
    exp_55_ram[2480] = 247;
    exp_55_ram[2481] = 7;
    exp_55_ram[2482] = 132;
    exp_55_ram[2483] = 196;
    exp_55_ram[2484] = 102;
    exp_55_ram[2485] = 7;
    exp_55_ram[2486] = 197;
    exp_55_ram[2487] = 118;
    exp_55_ram[2488] = 245;
    exp_55_ram[2489] = 6;
    exp_55_ram[2490] = 228;
    exp_55_ram[2491] = 244;
    exp_55_ram[2492] = 68;
    exp_55_ram[2493] = 7;
    exp_55_ram[2494] = 71;
    exp_55_ram[2495] = 231;
    exp_55_ram[2496] = 39;
    exp_55_ram[2497] = 7;
    exp_55_ram[2498] = 247;
    exp_55_ram[2499] = 7;
    exp_55_ram[2500] = 132;
    exp_55_ram[2501] = 196;
    exp_55_ram[2502] = 70;
    exp_55_ram[2503] = 7;
    exp_55_ram[2504] = 197;
    exp_55_ram[2505] = 86;
    exp_55_ram[2506] = 245;
    exp_55_ram[2507] = 6;
    exp_55_ram[2508] = 228;
    exp_55_ram[2509] = 244;
    exp_55_ram[2510] = 4;
    exp_55_ram[2511] = 7;
    exp_55_ram[2512] = 247;
    exp_55_ram[2513] = 7;
    exp_55_ram[2514] = 132;
    exp_55_ram[2515] = 196;
    exp_55_ram[2516] = 38;
    exp_55_ram[2517] = 7;
    exp_55_ram[2518] = 197;
    exp_55_ram[2519] = 54;
    exp_55_ram[2520] = 245;
    exp_55_ram[2521] = 6;
    exp_55_ram[2522] = 228;
    exp_55_ram[2523] = 244;
    exp_55_ram[2524] = 132;
    exp_55_ram[2525] = 196;
    exp_55_ram[2526] = 7;
    exp_55_ram[2527] = 7;
    exp_55_ram[2528] = 193;
    exp_55_ram[2529] = 129;
    exp_55_ram[2530] = 65;
    exp_55_ram[2531] = 1;
    exp_55_ram[2532] = 193;
    exp_55_ram[2533] = 129;
    exp_55_ram[2534] = 65;
    exp_55_ram[2535] = 1;
    exp_55_ram[2536] = 193;
    exp_55_ram[2537] = 129;
    exp_55_ram[2538] = 65;
    exp_55_ram[2539] = 1;
    exp_55_ram[2540] = 193;
    exp_55_ram[2541] = 1;
    exp_55_ram[2542] = 0;
    exp_55_ram[2543] = 1;
    exp_55_ram[2544] = 17;
    exp_55_ram[2545] = 129;
    exp_55_ram[2546] = 145;
    exp_55_ram[2547] = 33;
    exp_55_ram[2548] = 49;
    exp_55_ram[2549] = 1;
    exp_55_ram[2550] = 164;
    exp_55_ram[2551] = 196;
    exp_55_ram[2552] = 7;
    exp_55_ram[2553] = 71;
    exp_55_ram[2554] = 135;
    exp_55_ram[2555] = 199;
    exp_55_ram[2556] = 7;
    exp_55_ram[2557] = 71;
    exp_55_ram[2558] = 135;
    exp_55_ram[2559] = 199;
    exp_55_ram[2560] = 7;
    exp_55_ram[2561] = 100;
    exp_55_ram[2562] = 20;
    exp_55_ram[2563] = 4;
    exp_55_ram[2564] = 164;
    exp_55_ram[2565] = 180;
    exp_55_ram[2566] = 196;
    exp_55_ram[2567] = 212;
    exp_55_ram[2568] = 228;
    exp_55_ram[2569] = 244;
    exp_55_ram[2570] = 196;
    exp_55_ram[2571] = 4;
    exp_55_ram[2572] = 68;
    exp_55_ram[2573] = 132;
    exp_55_ram[2574] = 196;
    exp_55_ram[2575] = 4;
    exp_55_ram[2576] = 68;
    exp_55_ram[2577] = 132;
    exp_55_ram[2578] = 196;
    exp_55_ram[2579] = 100;
    exp_55_ram[2580] = 20;
    exp_55_ram[2581] = 4;
    exp_55_ram[2582] = 164;
    exp_55_ram[2583] = 180;
    exp_55_ram[2584] = 196;
    exp_55_ram[2585] = 212;
    exp_55_ram[2586] = 228;
    exp_55_ram[2587] = 244;
    exp_55_ram[2588] = 4;
    exp_55_ram[2589] = 7;
    exp_55_ram[2590] = 223;
    exp_55_ram[2591] = 164;
    exp_55_ram[2592] = 180;
    exp_55_ram[2593] = 196;
    exp_55_ram[2594] = 240;
    exp_55_ram[2595] = 4;
    exp_55_ram[2596] = 68;
    exp_55_ram[2597] = 255;
    exp_55_ram[2598] = 5;
    exp_55_ram[2599] = 240;
    exp_55_ram[2600] = 166;
    exp_55_ram[2601] = 7;
    exp_55_ram[2602] = 200;
    exp_55_ram[2603] = 182;
    exp_55_ram[2604] = 248;
    exp_55_ram[2605] = 6;
    exp_55_ram[2606] = 228;
    exp_55_ram[2607] = 244;
    exp_55_ram[2608] = 192;
    exp_55_ram[2609] = 196;
    exp_55_ram[2610] = 7;
    exp_55_ram[2611] = 196;
    exp_55_ram[2612] = 4;
    exp_55_ram[2613] = 68;
    exp_55_ram[2614] = 132;
    exp_55_ram[2615] = 196;
    exp_55_ram[2616] = 4;
    exp_55_ram[2617] = 68;
    exp_55_ram[2618] = 132;
    exp_55_ram[2619] = 196;
    exp_55_ram[2620] = 100;
    exp_55_ram[2621] = 20;
    exp_55_ram[2622] = 4;
    exp_55_ram[2623] = 164;
    exp_55_ram[2624] = 180;
    exp_55_ram[2625] = 196;
    exp_55_ram[2626] = 212;
    exp_55_ram[2627] = 228;
    exp_55_ram[2628] = 244;
    exp_55_ram[2629] = 4;
    exp_55_ram[2630] = 7;
    exp_55_ram[2631] = 15;
    exp_55_ram[2632] = 5;
    exp_55_ram[2633] = 7;
    exp_55_ram[2634] = 0;
    exp_55_ram[2635] = 6;
    exp_55_ram[2636] = 0;
    exp_55_ram[2637] = 192;
    exp_55_ram[2638] = 0;
    exp_55_ram[2639] = 0;
    exp_55_ram[2640] = 4;
    exp_55_ram[2641] = 68;
    exp_55_ram[2642] = 197;
    exp_55_ram[2643] = 7;
    exp_55_ram[2644] = 5;
    exp_55_ram[2645] = 213;
    exp_55_ram[2646] = 7;
    exp_55_ram[2647] = 6;
    exp_55_ram[2648] = 228;
    exp_55_ram[2649] = 244;
    exp_55_ram[2650] = 64;
    exp_55_ram[2651] = 4;
    exp_55_ram[2652] = 68;
    exp_55_ram[2653] = 228;
    exp_55_ram[2654] = 244;
    exp_55_ram[2655] = 0;
    exp_55_ram[2656] = 7;
    exp_55_ram[2657] = 7;
    exp_55_ram[2658] = 247;
    exp_55_ram[2659] = 7;
    exp_55_ram[2660] = 132;
    exp_55_ram[2661] = 196;
    exp_55_ram[2662] = 38;
    exp_55_ram[2663] = 7;
    exp_55_ram[2664] = 182;
    exp_55_ram[2665] = 54;
    exp_55_ram[2666] = 183;
    exp_55_ram[2667] = 6;
    exp_55_ram[2668] = 228;
    exp_55_ram[2669] = 244;
    exp_55_ram[2670] = 196;
    exp_55_ram[2671] = 4;
    exp_55_ram[2672] = 132;
    exp_55_ram[2673] = 196;
    exp_55_ram[2674] = 7;
    exp_55_ram[2675] = 0;
    exp_55_ram[2676] = 4;
    exp_55_ram[2677] = 68;
    exp_55_ram[2678] = 132;
    exp_55_ram[2679] = 196;
    exp_55_ram[2680] = 4;
    exp_55_ram[2681] = 68;
    exp_55_ram[2682] = 132;
    exp_55_ram[2683] = 196;
    exp_55_ram[2684] = 4;
    exp_55_ram[2685] = 100;
    exp_55_ram[2686] = 20;
    exp_55_ram[2687] = 4;
    exp_55_ram[2688] = 164;
    exp_55_ram[2689] = 180;
    exp_55_ram[2690] = 196;
    exp_55_ram[2691] = 212;
    exp_55_ram[2692] = 228;
    exp_55_ram[2693] = 244;
    exp_55_ram[2694] = 196;
    exp_55_ram[2695] = 240;
    exp_55_ram[2696] = 196;
    exp_55_ram[2697] = 16;
    exp_55_ram[2698] = 231;
    exp_55_ram[2699] = 128;
    exp_55_ram[2700] = 196;
    exp_55_ram[2701] = 7;
    exp_55_ram[2702] = 196;
    exp_55_ram[2703] = 4;
    exp_55_ram[2704] = 68;
    exp_55_ram[2705] = 132;
    exp_55_ram[2706] = 196;
    exp_55_ram[2707] = 4;
    exp_55_ram[2708] = 68;
    exp_55_ram[2709] = 132;
    exp_55_ram[2710] = 196;
    exp_55_ram[2711] = 100;
    exp_55_ram[2712] = 20;
    exp_55_ram[2713] = 4;
    exp_55_ram[2714] = 164;
    exp_55_ram[2715] = 180;
    exp_55_ram[2716] = 196;
    exp_55_ram[2717] = 212;
    exp_55_ram[2718] = 228;
    exp_55_ram[2719] = 244;
    exp_55_ram[2720] = 4;
    exp_55_ram[2721] = 7;
    exp_55_ram[2722] = 79;
    exp_55_ram[2723] = 5;
    exp_55_ram[2724] = 196;
    exp_55_ram[2725] = 231;
    exp_55_ram[2726] = 192;
    exp_55_ram[2727] = 196;
    exp_55_ram[2728] = 7;
    exp_55_ram[2729] = 132;
    exp_55_ram[2730] = 196;
    exp_55_ram[2731] = 7;
    exp_55_ram[2732] = 7;
    exp_55_ram[2733] = 193;
    exp_55_ram[2734] = 129;
    exp_55_ram[2735] = 65;
    exp_55_ram[2736] = 1;
    exp_55_ram[2737] = 193;
    exp_55_ram[2738] = 1;
    exp_55_ram[2739] = 0;
    exp_55_ram[2740] = 1;
    exp_55_ram[2741] = 17;
    exp_55_ram[2742] = 129;
    exp_55_ram[2743] = 33;
    exp_55_ram[2744] = 49;
    exp_55_ram[2745] = 65;
    exp_55_ram[2746] = 81;
    exp_55_ram[2747] = 97;
    exp_55_ram[2748] = 113;
    exp_55_ram[2749] = 1;
    exp_55_ram[2750] = 164;
    exp_55_ram[2751] = 143;
    exp_55_ram[2752] = 5;
    exp_55_ram[2753] = 5;
    exp_55_ram[2754] = 0;
    exp_55_ram[2755] = 6;
    exp_55_ram[2756] = 6;
    exp_55_ram[2757] = 0;
    exp_55_ram[2758] = 10;
    exp_55_ram[2759] = 10;
    exp_55_ram[2760] = 7;
    exp_55_ram[2761] = 7;
    exp_55_ram[2762] = 79;
    exp_55_ram[2763] = 5;
    exp_55_ram[2764] = 5;
    exp_55_ram[2765] = 228;
    exp_55_ram[2766] = 0;
    exp_55_ram[2767] = 135;
    exp_55_ram[2768] = 199;
    exp_55_ram[2769] = 196;
    exp_55_ram[2770] = 231;
    exp_55_ram[2771] = 244;
    exp_55_ram[2772] = 196;
    exp_55_ram[2773] = 7;
    exp_55_ram[2774] = 196;
    exp_55_ram[2775] = 7;
    exp_55_ram[2776] = 0;
    exp_55_ram[2777] = 196;
    exp_55_ram[2778] = 39;
    exp_55_ram[2779] = 55;
    exp_55_ram[2780] = 196;
    exp_55_ram[2781] = 7;
    exp_55_ram[2782] = 0;
    exp_55_ram[2783] = 11;
    exp_55_ram[2784] = 11;
    exp_55_ram[2785] = 7;
    exp_55_ram[2786] = 7;
    exp_55_ram[2787] = 193;
    exp_55_ram[2788] = 129;
    exp_55_ram[2789] = 65;
    exp_55_ram[2790] = 1;
    exp_55_ram[2791] = 193;
    exp_55_ram[2792] = 129;
    exp_55_ram[2793] = 65;
    exp_55_ram[2794] = 1;
    exp_55_ram[2795] = 1;
    exp_55_ram[2796] = 0;
    exp_55_ram[2797] = 1;
    exp_55_ram[2798] = 17;
    exp_55_ram[2799] = 129;
    exp_55_ram[2800] = 33;
    exp_55_ram[2801] = 49;
    exp_55_ram[2802] = 1;
    exp_55_ram[2803] = 164;
    exp_55_ram[2804] = 180;
    exp_55_ram[2805] = 15;
    exp_55_ram[2806] = 5;
    exp_55_ram[2807] = 5;
    exp_55_ram[2808] = 0;
    exp_55_ram[2809] = 6;
    exp_55_ram[2810] = 6;
    exp_55_ram[2811] = 0;
    exp_55_ram[2812] = 9;
    exp_55_ram[2813] = 9;
    exp_55_ram[2814] = 7;
    exp_55_ram[2815] = 7;
    exp_55_ram[2816] = 207;
    exp_55_ram[2817] = 5;
    exp_55_ram[2818] = 5;
    exp_55_ram[2819] = 228;
    exp_55_ram[2820] = 244;
    exp_55_ram[2821] = 132;
    exp_55_ram[2822] = 196;
    exp_55_ram[2823] = 132;
    exp_55_ram[2824] = 196;
    exp_55_ram[2825] = 167;
    exp_55_ram[2826] = 6;
    exp_55_ram[2827] = 7;
    exp_55_ram[2828] = 183;
    exp_55_ram[2829] = 6;
    exp_55_ram[2830] = 7;
    exp_55_ram[2831] = 6;
    exp_55_ram[2832] = 6;
    exp_55_ram[2833] = 0;
    exp_55_ram[2834] = 230;
    exp_55_ram[2835] = 246;
    exp_55_ram[2836] = 0;
    exp_55_ram[2837] = 193;
    exp_55_ram[2838] = 129;
    exp_55_ram[2839] = 65;
    exp_55_ram[2840] = 1;
    exp_55_ram[2841] = 1;
    exp_55_ram[2842] = 0;
    exp_55_ram[2843] = 1;
    exp_55_ram[2844] = 17;
    exp_55_ram[2845] = 129;
    exp_55_ram[2846] = 1;
    exp_55_ram[2847] = 164;
    exp_55_ram[2848] = 0;
    exp_55_ram[2849] = 135;
    exp_55_ram[2850] = 7;
    exp_55_ram[2851] = 71;
    exp_55_ram[2852] = 135;
    exp_55_ram[2853] = 199;
    exp_55_ram[2854] = 7;
    exp_55_ram[2855] = 164;
    exp_55_ram[2856] = 180;
    exp_55_ram[2857] = 196;
    exp_55_ram[2858] = 212;
    exp_55_ram[2859] = 228;
    exp_55_ram[2860] = 71;
    exp_55_ram[2861] = 244;
    exp_55_ram[2862] = 0;
    exp_55_ram[2863] = 7;
    exp_55_ram[2864] = 7;
    exp_55_ram[2865] = 71;
    exp_55_ram[2866] = 135;
    exp_55_ram[2867] = 199;
    exp_55_ram[2868] = 7;
    exp_55_ram[2869] = 71;
    exp_55_ram[2870] = 135;
    exp_55_ram[2871] = 199;
    exp_55_ram[2872] = 7;
    exp_55_ram[2873] = 196;
    exp_55_ram[2874] = 100;
    exp_55_ram[2875] = 20;
    exp_55_ram[2876] = 4;
    exp_55_ram[2877] = 164;
    exp_55_ram[2878] = 180;
    exp_55_ram[2879] = 196;
    exp_55_ram[2880] = 212;
    exp_55_ram[2881] = 228;
    exp_55_ram[2882] = 71;
    exp_55_ram[2883] = 244;
    exp_55_ram[2884] = 4;
    exp_55_ram[2885] = 192;
    exp_55_ram[2886] = 196;
    exp_55_ram[2887] = 135;
    exp_55_ram[2888] = 7;
    exp_55_ram[2889] = 23;
    exp_55_ram[2890] = 231;
    exp_55_ram[2891] = 196;
    exp_55_ram[2892] = 247;
    exp_55_ram[2893] = 4;
    exp_55_ram[2894] = 247;
    exp_55_ram[2895] = 71;
    exp_55_ram[2896] = 0;
    exp_55_ram[2897] = 7;
    exp_55_ram[2898] = 196;
    exp_55_ram[2899] = 246;
    exp_55_ram[2900] = 231;
    exp_55_ram[2901] = 196;
    exp_55_ram[2902] = 23;
    exp_55_ram[2903] = 244;
    exp_55_ram[2904] = 196;
    exp_55_ram[2905] = 32;
    exp_55_ram[2906] = 231;
    exp_55_ram[2907] = 0;
    exp_55_ram[2908] = 7;
    exp_55_ram[2909] = 0;
    exp_55_ram[2910] = 231;
    exp_55_ram[2911] = 4;
    exp_55_ram[2912] = 0;
    exp_55_ram[2913] = 196;
    exp_55_ram[2914] = 7;
    exp_55_ram[2915] = 7;
    exp_55_ram[2916] = 23;
    exp_55_ram[2917] = 231;
    exp_55_ram[2918] = 196;
    exp_55_ram[2919] = 247;
    exp_55_ram[2920] = 196;
    exp_55_ram[2921] = 71;
    exp_55_ram[2922] = 4;
    exp_55_ram[2923] = 230;
    exp_55_ram[2924] = 199;
    exp_55_ram[2925] = 0;
    exp_55_ram[2926] = 6;
    exp_55_ram[2927] = 246;
    exp_55_ram[2928] = 231;
    exp_55_ram[2929] = 196;
    exp_55_ram[2930] = 23;
    exp_55_ram[2931] = 244;
    exp_55_ram[2932] = 196;
    exp_55_ram[2933] = 32;
    exp_55_ram[2934] = 231;
    exp_55_ram[2935] = 0;
    exp_55_ram[2936] = 7;
    exp_55_ram[2937] = 0;
    exp_55_ram[2938] = 231;
    exp_55_ram[2939] = 196;
    exp_55_ram[2940] = 199;
    exp_55_ram[2941] = 160;
    exp_55_ram[2942] = 7;
    exp_55_ram[2943] = 128;
    exp_55_ram[2944] = 5;
    exp_55_ram[2945] = 5;
    exp_55_ram[2946] = 228;
    exp_55_ram[2947] = 244;
    exp_55_ram[2948] = 68;
    exp_55_ram[2949] = 247;
    exp_55_ram[2950] = 7;
    exp_55_ram[2951] = 247;
    exp_55_ram[2952] = 0;
    exp_55_ram[2953] = 7;
    exp_55_ram[2954] = 231;
    exp_55_ram[2955] = 132;
    exp_55_ram[2956] = 247;
    exp_55_ram[2957] = 7;
    exp_55_ram[2958] = 247;
    exp_55_ram[2959] = 0;
    exp_55_ram[2960] = 7;
    exp_55_ram[2961] = 231;
    exp_55_ram[2962] = 0;
    exp_55_ram[2963] = 7;
    exp_55_ram[2964] = 0;
    exp_55_ram[2965] = 231;
    exp_55_ram[2966] = 196;
    exp_55_ram[2967] = 135;
    exp_55_ram[2968] = 160;
    exp_55_ram[2969] = 7;
    exp_55_ram[2970] = 192;
    exp_55_ram[2971] = 5;
    exp_55_ram[2972] = 5;
    exp_55_ram[2973] = 228;
    exp_55_ram[2974] = 244;
    exp_55_ram[2975] = 68;
    exp_55_ram[2976] = 247;
    exp_55_ram[2977] = 7;
    exp_55_ram[2978] = 247;
    exp_55_ram[2979] = 0;
    exp_55_ram[2980] = 7;
    exp_55_ram[2981] = 231;
    exp_55_ram[2982] = 132;
    exp_55_ram[2983] = 247;
    exp_55_ram[2984] = 7;
    exp_55_ram[2985] = 247;
    exp_55_ram[2986] = 0;
    exp_55_ram[2987] = 7;
    exp_55_ram[2988] = 231;
    exp_55_ram[2989] = 0;
    exp_55_ram[2990] = 7;
    exp_55_ram[2991] = 160;
    exp_55_ram[2992] = 231;
    exp_55_ram[2993] = 196;
    exp_55_ram[2994] = 71;
    exp_55_ram[2995] = 160;
    exp_55_ram[2996] = 7;
    exp_55_ram[2997] = 0;
    exp_55_ram[2998] = 5;
    exp_55_ram[2999] = 5;
    exp_55_ram[3000] = 228;
    exp_55_ram[3001] = 244;
    exp_55_ram[3002] = 68;
    exp_55_ram[3003] = 247;
    exp_55_ram[3004] = 7;
    exp_55_ram[3005] = 247;
    exp_55_ram[3006] = 0;
    exp_55_ram[3007] = 7;
    exp_55_ram[3008] = 231;
    exp_55_ram[3009] = 132;
    exp_55_ram[3010] = 247;
    exp_55_ram[3011] = 7;
    exp_55_ram[3012] = 247;
    exp_55_ram[3013] = 0;
    exp_55_ram[3014] = 7;
    exp_55_ram[3015] = 231;
    exp_55_ram[3016] = 0;
    exp_55_ram[3017] = 7;
    exp_55_ram[3018] = 160;
    exp_55_ram[3019] = 231;
    exp_55_ram[3020] = 196;
    exp_55_ram[3021] = 7;
    exp_55_ram[3022] = 160;
    exp_55_ram[3023] = 7;
    exp_55_ram[3024] = 64;
    exp_55_ram[3025] = 5;
    exp_55_ram[3026] = 5;
    exp_55_ram[3027] = 228;
    exp_55_ram[3028] = 244;
    exp_55_ram[3029] = 68;
    exp_55_ram[3030] = 247;
    exp_55_ram[3031] = 7;
    exp_55_ram[3032] = 247;
    exp_55_ram[3033] = 0;
    exp_55_ram[3034] = 7;
    exp_55_ram[3035] = 231;
    exp_55_ram[3036] = 132;
    exp_55_ram[3037] = 247;
    exp_55_ram[3038] = 7;
    exp_55_ram[3039] = 247;
    exp_55_ram[3040] = 0;
    exp_55_ram[3041] = 7;
    exp_55_ram[3042] = 231;
    exp_55_ram[3043] = 0;
    exp_55_ram[3044] = 7;
    exp_55_ram[3045] = 0;
    exp_55_ram[3046] = 231;
    exp_55_ram[3047] = 196;
    exp_55_ram[3048] = 71;
    exp_55_ram[3049] = 199;
    exp_55_ram[3050] = 128;
    exp_55_ram[3051] = 7;
    exp_55_ram[3052] = 64;
    exp_55_ram[3053] = 5;
    exp_55_ram[3054] = 5;
    exp_55_ram[3055] = 228;
    exp_55_ram[3056] = 244;
    exp_55_ram[3057] = 68;
    exp_55_ram[3058] = 247;
    exp_55_ram[3059] = 7;
    exp_55_ram[3060] = 247;
    exp_55_ram[3061] = 0;
    exp_55_ram[3062] = 7;
    exp_55_ram[3063] = 231;
    exp_55_ram[3064] = 132;
    exp_55_ram[3065] = 64;
    exp_55_ram[3066] = 7;
    exp_55_ram[3067] = 128;
    exp_55_ram[3068] = 5;
    exp_55_ram[3069] = 5;
    exp_55_ram[3070] = 228;
    exp_55_ram[3071] = 244;
    exp_55_ram[3072] = 68;
    exp_55_ram[3073] = 247;
    exp_55_ram[3074] = 7;
    exp_55_ram[3075] = 247;
    exp_55_ram[3076] = 0;
    exp_55_ram[3077] = 7;
    exp_55_ram[3078] = 231;
    exp_55_ram[3079] = 132;
    exp_55_ram[3080] = 160;
    exp_55_ram[3081] = 7;
    exp_55_ram[3082] = 192;
    exp_55_ram[3083] = 5;
    exp_55_ram[3084] = 5;
    exp_55_ram[3085] = 228;
    exp_55_ram[3086] = 244;
    exp_55_ram[3087] = 68;
    exp_55_ram[3088] = 247;
    exp_55_ram[3089] = 7;
    exp_55_ram[3090] = 247;
    exp_55_ram[3091] = 0;
    exp_55_ram[3092] = 7;
    exp_55_ram[3093] = 231;
    exp_55_ram[3094] = 132;
    exp_55_ram[3095] = 247;
    exp_55_ram[3096] = 7;
    exp_55_ram[3097] = 247;
    exp_55_ram[3098] = 0;
    exp_55_ram[3099] = 7;
    exp_55_ram[3100] = 231;
    exp_55_ram[3101] = 0;
    exp_55_ram[3102] = 7;
    exp_55_ram[3103] = 160;
    exp_55_ram[3104] = 231;
    exp_55_ram[3105] = 0;
    exp_55_ram[3106] = 7;
    exp_55_ram[3107] = 7;
    exp_55_ram[3108] = 0;
    exp_55_ram[3109] = 7;
    exp_55_ram[3110] = 7;
    exp_55_ram[3111] = 193;
    exp_55_ram[3112] = 129;
    exp_55_ram[3113] = 1;
    exp_55_ram[3114] = 0;
    exp_55_ram[3115] = 1;
    exp_55_ram[3116] = 17;
    exp_55_ram[3117] = 129;
    exp_55_ram[3118] = 1;
    exp_55_ram[3119] = 164;
    exp_55_ram[3120] = 196;
    exp_55_ram[3121] = 64;
    exp_55_ram[3122] = 5;
    exp_55_ram[3123] = 7;
    exp_55_ram[3124] = 223;
    exp_55_ram[3125] = 5;
    exp_55_ram[3126] = 7;
    exp_55_ram[3127] = 193;
    exp_55_ram[3128] = 129;
    exp_55_ram[3129] = 1;
    exp_55_ram[3130] = 0;
    exp_55_ram[3131] = 1;
    exp_55_ram[3132] = 17;
    exp_55_ram[3133] = 129;
    exp_55_ram[3134] = 33;
    exp_55_ram[3135] = 49;
    exp_55_ram[3136] = 65;
    exp_55_ram[3137] = 81;
    exp_55_ram[3138] = 97;
    exp_55_ram[3139] = 113;
    exp_55_ram[3140] = 129;
    exp_55_ram[3141] = 145;
    exp_55_ram[3142] = 1;
    exp_55_ram[3143] = 164;
    exp_55_ram[3144] = 180;
    exp_55_ram[3145] = 196;
    exp_55_ram[3146] = 32;
    exp_55_ram[3147] = 244;
    exp_55_ram[3148] = 64;
    exp_55_ram[3149] = 244;
    exp_55_ram[3150] = 132;
    exp_55_ram[3151] = 7;
    exp_55_ram[3152] = 207;
    exp_55_ram[3153] = 164;
    exp_55_ram[3154] = 196;
    exp_55_ram[3155] = 1;
    exp_55_ram[3156] = 7;
    exp_55_ram[3157] = 247;
    exp_55_ram[3158] = 244;
    exp_55_ram[3159] = 132;
    exp_55_ram[3160] = 7;
    exp_55_ram[3161] = 0;
    exp_55_ram[3162] = 68;
    exp_55_ram[3163] = 12;
    exp_55_ram[3164] = 231;
    exp_55_ram[3165] = 68;
    exp_55_ram[3166] = 12;
    exp_55_ram[3167] = 231;
    exp_55_ram[3168] = 4;
    exp_55_ram[3169] = 12;
    exp_55_ram[3170] = 231;
    exp_55_ram[3171] = 132;
    exp_55_ram[3172] = 23;
    exp_55_ram[3173] = 244;
    exp_55_ram[3174] = 196;
    exp_55_ram[3175] = 7;
    exp_55_ram[3176] = 196;
    exp_55_ram[3177] = 247;
    exp_55_ram[3178] = 244;
    exp_55_ram[3179] = 132;
    exp_55_ram[3180] = 7;
    exp_55_ram[3181] = 0;
    exp_55_ram[3182] = 4;
    exp_55_ram[3183] = 68;
    exp_55_ram[3184] = 70;
    exp_55_ram[3185] = 7;
    exp_55_ram[3186] = 182;
    exp_55_ram[3187] = 86;
    exp_55_ram[3188] = 183;
    exp_55_ram[3189] = 6;
    exp_55_ram[3190] = 228;
    exp_55_ram[3191] = 244;
    exp_55_ram[3192] = 159;
    exp_55_ram[3193] = 0;
    exp_55_ram[3194] = 4;
    exp_55_ram[3195] = 4;
    exp_55_ram[3196] = 132;
    exp_55_ram[3197] = 7;
    exp_55_ram[3198] = 68;
    exp_55_ram[3199] = 7;
    exp_55_ram[3200] = 7;
    exp_55_ram[3201] = 207;
    exp_55_ram[3202] = 164;
    exp_55_ram[3203] = 196;
    exp_55_ram[3204] = 1;
    exp_55_ram[3205] = 7;
    exp_55_ram[3206] = 247;
    exp_55_ram[3207] = 244;
    exp_55_ram[3208] = 132;
    exp_55_ram[3209] = 7;
    exp_55_ram[3210] = 0;
    exp_55_ram[3211] = 68;
    exp_55_ram[3212] = 11;
    exp_55_ram[3213] = 231;
    exp_55_ram[3214] = 68;
    exp_55_ram[3215] = 11;
    exp_55_ram[3216] = 231;
    exp_55_ram[3217] = 4;
    exp_55_ram[3218] = 11;
    exp_55_ram[3219] = 231;
    exp_55_ram[3220] = 68;
    exp_55_ram[3221] = 23;
    exp_55_ram[3222] = 244;
    exp_55_ram[3223] = 196;
    exp_55_ram[3224] = 7;
    exp_55_ram[3225] = 196;
    exp_55_ram[3226] = 247;
    exp_55_ram[3227] = 244;
    exp_55_ram[3228] = 4;
    exp_55_ram[3229] = 7;
    exp_55_ram[3230] = 196;
    exp_55_ram[3231] = 247;
    exp_55_ram[3232] = 244;
    exp_55_ram[3233] = 132;
    exp_55_ram[3234] = 7;
    exp_55_ram[3235] = 0;
    exp_55_ram[3236] = 4;
    exp_55_ram[3237] = 68;
    exp_55_ram[3238] = 38;
    exp_55_ram[3239] = 7;
    exp_55_ram[3240] = 182;
    exp_55_ram[3241] = 54;
    exp_55_ram[3242] = 183;
    exp_55_ram[3243] = 6;
    exp_55_ram[3244] = 228;
    exp_55_ram[3245] = 244;
    exp_55_ram[3246] = 159;
    exp_55_ram[3247] = 0;
    exp_55_ram[3248] = 132;
    exp_55_ram[3249] = 71;
    exp_55_ram[3250] = 244;
    exp_55_ram[3251] = 4;
    exp_55_ram[3252] = 1;
    exp_55_ram[3253] = 7;
    exp_55_ram[3254] = 7;
    exp_55_ram[3255] = 144;
    exp_55_ram[3256] = 5;
    exp_55_ram[3257] = 5;
    exp_55_ram[3258] = 228;
    exp_55_ram[3259] = 244;
    exp_55_ram[3260] = 196;
    exp_55_ram[3261] = 23;
    exp_55_ram[3262] = 244;
    exp_55_ram[3263] = 196;
    exp_55_ram[3264] = 196;
    exp_55_ram[3265] = 247;
    exp_55_ram[3266] = 244;
    exp_55_ram[3267] = 196;
    exp_55_ram[3268] = 112;
    exp_55_ram[3269] = 247;
    exp_55_ram[3270] = 244;
    exp_55_ram[3271] = 4;
    exp_55_ram[3272] = 196;
    exp_55_ram[3273] = 247;
    exp_55_ram[3274] = 244;
    exp_55_ram[3275] = 4;
    exp_55_ram[3276] = 244;
    exp_55_ram[3277] = 247;
    exp_55_ram[3278] = 244;
    exp_55_ram[3279] = 4;
    exp_55_ram[3280] = 0;
    exp_55_ram[3281] = 7;
    exp_55_ram[3282] = 7;
    exp_55_ram[3283] = 144;
    exp_55_ram[3284] = 5;
    exp_55_ram[3285] = 5;
    exp_55_ram[3286] = 228;
    exp_55_ram[3287] = 244;
    exp_55_ram[3288] = 196;
    exp_55_ram[3289] = 244;
    exp_55_ram[3290] = 4;
    exp_55_ram[3291] = 244;
    exp_55_ram[3292] = 247;
    exp_55_ram[3293] = 244;
    exp_55_ram[3294] = 4;
    exp_55_ram[3295] = 192;
    exp_55_ram[3296] = 7;
    exp_55_ram[3297] = 16;
    exp_55_ram[3298] = 5;
    exp_55_ram[3299] = 5;
    exp_55_ram[3300] = 228;
    exp_55_ram[3301] = 244;
    exp_55_ram[3302] = 196;
    exp_55_ram[3303] = 244;
    exp_55_ram[3304] = 4;
    exp_55_ram[3305] = 244;
    exp_55_ram[3306] = 247;
    exp_55_ram[3307] = 244;
    exp_55_ram[3308] = 4;
    exp_55_ram[3309] = 244;
    exp_55_ram[3310] = 196;
    exp_55_ram[3311] = 68;
    exp_55_ram[3312] = 132;
    exp_55_ram[3313] = 196;
    exp_55_ram[3314] = 4;
    exp_55_ram[3315] = 68;
    exp_55_ram[3316] = 132;
    exp_55_ram[3317] = 196;
    exp_55_ram[3318] = 4;
    exp_55_ram[3319] = 68;
    exp_55_ram[3320] = 199;
    exp_55_ram[3321] = 103;
    exp_55_ram[3322] = 23;
    exp_55_ram[3323] = 7;
    exp_55_ram[3324] = 167;
    exp_55_ram[3325] = 183;
    exp_55_ram[3326] = 199;
    exp_55_ram[3327] = 215;
    exp_55_ram[3328] = 231;
    exp_55_ram[3329] = 196;
    exp_55_ram[3330] = 193;
    exp_55_ram[3331] = 129;
    exp_55_ram[3332] = 65;
    exp_55_ram[3333] = 1;
    exp_55_ram[3334] = 193;
    exp_55_ram[3335] = 129;
    exp_55_ram[3336] = 65;
    exp_55_ram[3337] = 1;
    exp_55_ram[3338] = 193;
    exp_55_ram[3339] = 129;
    exp_55_ram[3340] = 1;
    exp_55_ram[3341] = 0;
    exp_55_ram[3342] = 1;
    exp_55_ram[3343] = 17;
    exp_55_ram[3344] = 129;
    exp_55_ram[3345] = 145;
    exp_55_ram[3346] = 33;
    exp_55_ram[3347] = 49;
    exp_55_ram[3348] = 1;
    exp_55_ram[3349] = 164;
    exp_55_ram[3350] = 0;
    exp_55_ram[3351] = 0;
    exp_55_ram[3352] = 244;
    exp_55_ram[3353] = 4;
    exp_55_ram[3354] = 196;
    exp_55_ram[3355] = 7;
    exp_55_ram[3356] = 71;
    exp_55_ram[3357] = 228;
    exp_55_ram[3358] = 244;
    exp_55_ram[3359] = 4;
    exp_55_ram[3360] = 68;
    exp_55_ram[3361] = 159;
    exp_55_ram[3362] = 5;
    exp_55_ram[3363] = 7;
    exp_55_ram[3364] = 0;
    exp_55_ram[3365] = 7;
    exp_55_ram[3366] = 0;
    exp_55_ram[3367] = 228;
    exp_55_ram[3368] = 244;
    exp_55_ram[3369] = 0;
    exp_55_ram[3370] = 7;
    exp_55_ram[3371] = 7;
    exp_55_ram[3372] = 247;
    exp_55_ram[3373] = 7;
    exp_55_ram[3374] = 4;
    exp_55_ram[3375] = 68;
    exp_55_ram[3376] = 201;
    exp_55_ram[3377] = 7;
    exp_55_ram[3378] = 37;
    exp_55_ram[3379] = 217;
    exp_55_ram[3380] = 245;
    exp_55_ram[3381] = 6;
    exp_55_ram[3382] = 7;
    exp_55_ram[3383] = 7;
    exp_55_ram[3384] = 132;
    exp_55_ram[3385] = 196;
    exp_55_ram[3386] = 166;
    exp_55_ram[3387] = 7;
    exp_55_ram[3388] = 200;
    exp_55_ram[3389] = 182;
    exp_55_ram[3390] = 248;
    exp_55_ram[3391] = 6;
    exp_55_ram[3392] = 228;
    exp_55_ram[3393] = 244;
    exp_55_ram[3394] = 0;
    exp_55_ram[3395] = 199;
    exp_55_ram[3396] = 4;
    exp_55_ram[3397] = 132;
    exp_55_ram[3398] = 196;
    exp_55_ram[3399] = 7;
    exp_55_ram[3400] = 223;
    exp_55_ram[3401] = 4;
    exp_55_ram[3402] = 68;
    exp_55_ram[3403] = 132;
    exp_55_ram[3404] = 196;
    exp_55_ram[3405] = 4;
    exp_55_ram[3406] = 68;
    exp_55_ram[3407] = 132;
    exp_55_ram[3408] = 196;
    exp_55_ram[3409] = 4;
    exp_55_ram[3410] = 100;
    exp_55_ram[3411] = 20;
    exp_55_ram[3412] = 4;
    exp_55_ram[3413] = 164;
    exp_55_ram[3414] = 180;
    exp_55_ram[3415] = 196;
    exp_55_ram[3416] = 212;
    exp_55_ram[3417] = 228;
    exp_55_ram[3418] = 244;
    exp_55_ram[3419] = 4;
    exp_55_ram[3420] = 68;
    exp_55_ram[3421] = 159;
    exp_55_ram[3422] = 5;
    exp_55_ram[3423] = 0;
    exp_55_ram[3424] = 199;
    exp_55_ram[3425] = 231;
    exp_55_ram[3426] = 0;
    exp_55_ram[3427] = 199;
    exp_55_ram[3428] = 7;
    exp_55_ram[3429] = 193;
    exp_55_ram[3430] = 129;
    exp_55_ram[3431] = 65;
    exp_55_ram[3432] = 1;
    exp_55_ram[3433] = 193;
    exp_55_ram[3434] = 1;
    exp_55_ram[3435] = 0;
    exp_55_ram[3436] = 1;
    exp_55_ram[3437] = 17;
    exp_55_ram[3438] = 129;
    exp_55_ram[3439] = 1;
    exp_55_ram[3440] = 164;
    exp_55_ram[3441] = 4;
    exp_55_ram[3442] = 196;
    exp_55_ram[3443] = 79;
    exp_55_ram[3444] = 5;
    exp_55_ram[3445] = 244;
    exp_55_ram[3446] = 180;
    exp_55_ram[3447] = 7;
    exp_55_ram[3448] = 144;
    exp_55_ram[3449] = 231;
    exp_55_ram[3450] = 196;
    exp_55_ram[3451] = 7;
    exp_55_ram[3452] = 39;
    exp_55_ram[3453] = 231;
    exp_55_ram[3454] = 23;
    exp_55_ram[3455] = 244;
    exp_55_ram[3456] = 180;
    exp_55_ram[3457] = 196;
    exp_55_ram[3458] = 247;
    exp_55_ram[3459] = 7;
    exp_55_ram[3460] = 244;
    exp_55_ram[3461] = 95;
    exp_55_ram[3462] = 0;
    exp_55_ram[3463] = 196;
    exp_55_ram[3464] = 7;
    exp_55_ram[3465] = 193;
    exp_55_ram[3466] = 129;
    exp_55_ram[3467] = 1;
    exp_55_ram[3468] = 0;
    exp_55_ram[3469] = 1;
    exp_55_ram[3470] = 17;
    exp_55_ram[3471] = 129;
    exp_55_ram[3472] = 1;
    exp_55_ram[3473] = 0;
    exp_55_ram[3474] = 71;
    exp_55_ram[3475] = 7;
    exp_55_ram[3476] = 31;
    exp_55_ram[3477] = 5;
    exp_55_ram[3478] = 7;
    exp_55_ram[3479] = 193;
    exp_55_ram[3480] = 129;
    exp_55_ram[3481] = 1;
    exp_55_ram[3482] = 0;
    exp_55_ram[3483] = 1;
    exp_55_ram[3484] = 17;
    exp_55_ram[3485] = 129;
    exp_55_ram[3486] = 33;
    exp_55_ram[3487] = 49;
    exp_55_ram[3488] = 1;
    exp_55_ram[3489] = 164;
    exp_55_ram[3490] = 223;
    exp_55_ram[3491] = 164;
    exp_55_ram[3492] = 180;
    exp_55_ram[3493] = 0;
    exp_55_ram[3494] = 223;
    exp_55_ram[3495] = 5;
    exp_55_ram[3496] = 5;
    exp_55_ram[3497] = 132;
    exp_55_ram[3498] = 196;
    exp_55_ram[3499] = 166;
    exp_55_ram[3500] = 7;
    exp_55_ram[3501] = 6;
    exp_55_ram[3502] = 182;
    exp_55_ram[3503] = 7;
    exp_55_ram[3504] = 6;
    exp_55_ram[3505] = 196;
    exp_55_ram[3506] = 6;
    exp_55_ram[3507] = 0;
    exp_55_ram[3508] = 9;
    exp_55_ram[3509] = 7;
    exp_55_ram[3510] = 198;
    exp_55_ram[3511] = 9;
    exp_55_ram[3512] = 7;
    exp_55_ram[3513] = 214;
    exp_55_ram[3514] = 9;
    exp_55_ram[3515] = 7;
    exp_55_ram[3516] = 215;
    exp_55_ram[3517] = 0;
    exp_55_ram[3518] = 7;
    exp_55_ram[3519] = 193;
    exp_55_ram[3520] = 129;
    exp_55_ram[3521] = 65;
    exp_55_ram[3522] = 1;
    exp_55_ram[3523] = 1;
    exp_55_ram[3524] = 0;
    exp_55_ram[3525] = 1;
    exp_55_ram[3526] = 17;
    exp_55_ram[3527] = 129;
    exp_55_ram[3528] = 1;
    exp_55_ram[3529] = 0;
    exp_55_ram[3530] = 135;
    exp_55_ram[3531] = 207;
    exp_55_ram[3532] = 0;
    exp_55_ram[3533] = 193;
    exp_55_ram[3534] = 129;
    exp_55_ram[3535] = 1;
    exp_55_ram[3536] = 0;
    exp_55_ram[3537] = 1;
    exp_55_ram[3538] = 17;
    exp_55_ram[3539] = 129;
    exp_55_ram[3540] = 1;
    exp_55_ram[3541] = 0;
    exp_55_ram[3542] = 135;
    exp_55_ram[3543] = 207;
    exp_55_ram[3544] = 16;
    exp_55_ram[3545] = 244;
    exp_55_ram[3546] = 4;
    exp_55_ram[3547] = 0;
    exp_55_ram[3548] = 132;
    exp_55_ram[3549] = 0;
    exp_55_ram[3550] = 135;
    exp_55_ram[3551] = 207;
    exp_55_ram[3552] = 192;
    exp_55_ram[3553] = 196;
    exp_55_ram[3554] = 23;
    exp_55_ram[3555] = 244;
    exp_55_ram[3556] = 0;
    exp_55_ram[3557] = 199;
    exp_55_ram[3558] = 7;
    exp_55_ram[3559] = 196;
    exp_55_ram[3560] = 15;
    exp_55_ram[3561] = 0;
    exp_55_ram[3562] = 7;
    exp_55_ram[3563] = 160;
    exp_55_ram[3564] = 247;
    exp_55_ram[3565] = 7;
    exp_55_ram[3566] = 95;
    exp_55_ram[3567] = 196;
    exp_55_ram[3568] = 240;
    exp_55_ram[3569] = 231;
    exp_55_ram[3570] = 192;
    exp_55_ram[3571] = 196;
    exp_55_ram[3572] = 23;
    exp_55_ram[3573] = 244;
    exp_55_ram[3574] = 0;
    exp_55_ram[3575] = 199;
    exp_55_ram[3576] = 7;
    exp_55_ram[3577] = 196;
    exp_55_ram[3578] = 143;
    exp_55_ram[3579] = 0;
    exp_55_ram[3580] = 7;
    exp_55_ram[3581] = 160;
    exp_55_ram[3582] = 247;
    exp_55_ram[3583] = 7;
    exp_55_ram[3584] = 223;
    exp_55_ram[3585] = 196;
    exp_55_ram[3586] = 16;
    exp_55_ram[3587] = 231;
    exp_55_ram[3588] = 132;
    exp_55_ram[3589] = 23;
    exp_55_ram[3590] = 244;
    exp_55_ram[3591] = 132;
    exp_55_ram[3592] = 144;
    exp_55_ram[3593] = 231;
    exp_55_ram[3594] = 0;
    exp_55_ram[3595] = 199;
    exp_55_ram[3596] = 7;
    exp_55_ram[3597] = 0;
    exp_55_ram[3598] = 143;
    exp_55_ram[3599] = 0;
    exp_55_ram[3600] = 193;
    exp_55_ram[3601] = 129;
    exp_55_ram[3602] = 1;
    exp_55_ram[3603] = 0;
    exp_55_ram[3604] = 1;
    exp_55_ram[3605] = 17;
    exp_55_ram[3606] = 129;
    exp_55_ram[3607] = 33;
    exp_55_ram[3608] = 49;
    exp_55_ram[3609] = 65;
    exp_55_ram[3610] = 81;
    exp_55_ram[3611] = 97;
    exp_55_ram[3612] = 113;
    exp_55_ram[3613] = 129;
    exp_55_ram[3614] = 145;
    exp_55_ram[3615] = 161;
    exp_55_ram[3616] = 177;
    exp_55_ram[3617] = 1;
    exp_55_ram[3618] = 16;
    exp_55_ram[3619] = 244;
    exp_55_ram[3620] = 16;
    exp_55_ram[3621] = 0;
    exp_55_ram[3622] = 228;
    exp_55_ram[3623] = 244;
    exp_55_ram[3624] = 95;
    exp_55_ram[3625] = 164;
    exp_55_ram[3626] = 180;
    exp_55_ram[3627] = 4;
    exp_55_ram[3628] = 0;
    exp_55_ram[3629] = 196;
    exp_55_ram[3630] = 52;
    exp_55_ram[3631] = 135;
    exp_55_ram[3632] = 247;
    exp_55_ram[3633] = 244;
    exp_55_ram[3634] = 196;
    exp_55_ram[3635] = 52;
    exp_55_ram[3636] = 135;
    exp_55_ram[3637] = 247;
    exp_55_ram[3638] = 244;
    exp_55_ram[3639] = 196;
    exp_55_ram[3640] = 52;
    exp_55_ram[3641] = 135;
    exp_55_ram[3642] = 247;
    exp_55_ram[3643] = 244;
    exp_55_ram[3644] = 196;
    exp_55_ram[3645] = 52;
    exp_55_ram[3646] = 135;
    exp_55_ram[3647] = 247;
    exp_55_ram[3648] = 244;
    exp_55_ram[3649] = 196;
    exp_55_ram[3650] = 71;
    exp_55_ram[3651] = 244;
    exp_55_ram[3652] = 95;
    exp_55_ram[3653] = 5;
    exp_55_ram[3654] = 5;
    exp_55_ram[3655] = 4;
    exp_55_ram[3656] = 68;
    exp_55_ram[3657] = 166;
    exp_55_ram[3658] = 7;
    exp_55_ram[3659] = 6;
    exp_55_ram[3660] = 182;
    exp_55_ram[3661] = 7;
    exp_55_ram[3662] = 6;
    exp_55_ram[3663] = 0;
    exp_55_ram[3664] = 6;
    exp_55_ram[3665] = 212;
    exp_55_ram[3666] = 4;
    exp_55_ram[3667] = 132;
    exp_55_ram[3668] = 196;
    exp_55_ram[3669] = 5;
    exp_55_ram[3670] = 7;
    exp_55_ram[3671] = 198;
    exp_55_ram[3672] = 5;
    exp_55_ram[3673] = 7;
    exp_55_ram[3674] = 214;
    exp_55_ram[3675] = 5;
    exp_55_ram[3676] = 7;
    exp_55_ram[3677] = 215;
    exp_55_ram[3678] = 196;
    exp_55_ram[3679] = 0;
    exp_55_ram[3680] = 199;
    exp_55_ram[3681] = 79;
    exp_55_ram[3682] = 223;
    exp_55_ram[3683] = 164;
    exp_55_ram[3684] = 180;
    exp_55_ram[3685] = 4;
    exp_55_ram[3686] = 0;
    exp_55_ram[3687] = 4;
    exp_55_ram[3688] = 68;
    exp_55_ram[3689] = 52;
    exp_55_ram[3690] = 134;
    exp_55_ram[3691] = 215;
    exp_55_ram[3692] = 0;
    exp_55_ram[3693] = 215;
    exp_55_ram[3694] = 214;
    exp_55_ram[3695] = 52;
    exp_55_ram[3696] = 134;
    exp_55_ram[3697] = 215;
    exp_55_ram[3698] = 215;
    exp_55_ram[3699] = 5;
    exp_55_ram[3700] = 54;
    exp_55_ram[3701] = 7;
    exp_55_ram[3702] = 36;
    exp_55_ram[3703] = 52;
    exp_55_ram[3704] = 4;
    exp_55_ram[3705] = 68;
    exp_55_ram[3706] = 52;
    exp_55_ram[3707] = 134;
    exp_55_ram[3708] = 215;
    exp_55_ram[3709] = 0;
    exp_55_ram[3710] = 215;
    exp_55_ram[3711] = 214;
    exp_55_ram[3712] = 52;
    exp_55_ram[3713] = 134;
    exp_55_ram[3714] = 215;
    exp_55_ram[3715] = 215;
    exp_55_ram[3716] = 5;
    exp_55_ram[3717] = 86;
    exp_55_ram[3718] = 7;
    exp_55_ram[3719] = 68;
    exp_55_ram[3720] = 84;
    exp_55_ram[3721] = 4;
    exp_55_ram[3722] = 68;
    exp_55_ram[3723] = 52;
    exp_55_ram[3724] = 134;
    exp_55_ram[3725] = 215;
    exp_55_ram[3726] = 0;
    exp_55_ram[3727] = 215;
    exp_55_ram[3728] = 214;
    exp_55_ram[3729] = 52;
    exp_55_ram[3730] = 134;
    exp_55_ram[3731] = 215;
    exp_55_ram[3732] = 215;
    exp_55_ram[3733] = 5;
    exp_55_ram[3734] = 118;
    exp_55_ram[3735] = 7;
    exp_55_ram[3736] = 100;
    exp_55_ram[3737] = 116;
    exp_55_ram[3738] = 4;
    exp_55_ram[3739] = 68;
    exp_55_ram[3740] = 52;
    exp_55_ram[3741] = 134;
    exp_55_ram[3742] = 215;
    exp_55_ram[3743] = 0;
    exp_55_ram[3744] = 215;
    exp_55_ram[3745] = 214;
    exp_55_ram[3746] = 52;
    exp_55_ram[3747] = 134;
    exp_55_ram[3748] = 215;
    exp_55_ram[3749] = 215;
    exp_55_ram[3750] = 5;
    exp_55_ram[3751] = 150;
    exp_55_ram[3752] = 7;
    exp_55_ram[3753] = 132;
    exp_55_ram[3754] = 148;
    exp_55_ram[3755] = 196;
    exp_55_ram[3756] = 71;
    exp_55_ram[3757] = 244;
    exp_55_ram[3758] = 223;
    exp_55_ram[3759] = 5;
    exp_55_ram[3760] = 5;
    exp_55_ram[3761] = 4;
    exp_55_ram[3762] = 68;
    exp_55_ram[3763] = 166;
    exp_55_ram[3764] = 7;
    exp_55_ram[3765] = 6;
    exp_55_ram[3766] = 182;
    exp_55_ram[3767] = 7;
    exp_55_ram[3768] = 6;
    exp_55_ram[3769] = 0;
    exp_55_ram[3770] = 6;
    exp_55_ram[3771] = 212;
    exp_55_ram[3772] = 4;
    exp_55_ram[3773] = 4;
    exp_55_ram[3774] = 68;
    exp_55_ram[3775] = 5;
    exp_55_ram[3776] = 7;
    exp_55_ram[3777] = 198;
    exp_55_ram[3778] = 5;
    exp_55_ram[3779] = 7;
    exp_55_ram[3780] = 214;
    exp_55_ram[3781] = 5;
    exp_55_ram[3782] = 7;
    exp_55_ram[3783] = 215;
    exp_55_ram[3784] = 196;
    exp_55_ram[3785] = 0;
    exp_55_ram[3786] = 135;
    exp_55_ram[3787] = 207;
    exp_55_ram[3788] = 79;
    exp_55_ram[3789] = 164;
    exp_55_ram[3790] = 180;
    exp_55_ram[3791] = 4;
    exp_55_ram[3792] = 0;
    exp_55_ram[3793] = 196;
    exp_55_ram[3794] = 52;
    exp_55_ram[3795] = 135;
    exp_55_ram[3796] = 247;
    exp_55_ram[3797] = 244;
    exp_55_ram[3798] = 196;
    exp_55_ram[3799] = 52;
    exp_55_ram[3800] = 135;
    exp_55_ram[3801] = 247;
    exp_55_ram[3802] = 244;
    exp_55_ram[3803] = 196;
    exp_55_ram[3804] = 52;
    exp_55_ram[3805] = 135;
    exp_55_ram[3806] = 247;
    exp_55_ram[3807] = 244;
    exp_55_ram[3808] = 196;
    exp_55_ram[3809] = 52;
    exp_55_ram[3810] = 135;
    exp_55_ram[3811] = 247;
    exp_55_ram[3812] = 244;
    exp_55_ram[3813] = 196;
    exp_55_ram[3814] = 71;
    exp_55_ram[3815] = 244;
    exp_55_ram[3816] = 79;
    exp_55_ram[3817] = 5;
    exp_55_ram[3818] = 5;
    exp_55_ram[3819] = 4;
    exp_55_ram[3820] = 68;
    exp_55_ram[3821] = 166;
    exp_55_ram[3822] = 7;
    exp_55_ram[3823] = 6;
    exp_55_ram[3824] = 182;
    exp_55_ram[3825] = 7;
    exp_55_ram[3826] = 6;
    exp_55_ram[3827] = 0;
    exp_55_ram[3828] = 6;
    exp_55_ram[3829] = 212;
    exp_55_ram[3830] = 4;
    exp_55_ram[3831] = 132;
    exp_55_ram[3832] = 196;
    exp_55_ram[3833] = 5;
    exp_55_ram[3834] = 7;
    exp_55_ram[3835] = 198;
    exp_55_ram[3836] = 5;
    exp_55_ram[3837] = 7;
    exp_55_ram[3838] = 214;
    exp_55_ram[3839] = 5;
    exp_55_ram[3840] = 7;
    exp_55_ram[3841] = 215;
    exp_55_ram[3842] = 196;
    exp_55_ram[3843] = 0;
    exp_55_ram[3844] = 71;
    exp_55_ram[3845] = 79;
    exp_55_ram[3846] = 207;
    exp_55_ram[3847] = 164;
    exp_55_ram[3848] = 180;
    exp_55_ram[3849] = 4;
    exp_55_ram[3850] = 0;
    exp_55_ram[3851] = 4;
    exp_55_ram[3852] = 68;
    exp_55_ram[3853] = 52;
    exp_55_ram[3854] = 134;
    exp_55_ram[3855] = 0;
    exp_55_ram[3856] = 7;
    exp_55_ram[3857] = 7;
    exp_55_ram[3858] = 79;
    exp_55_ram[3859] = 5;
    exp_55_ram[3860] = 5;
    exp_55_ram[3861] = 228;
    exp_55_ram[3862] = 244;
    exp_55_ram[3863] = 4;
    exp_55_ram[3864] = 68;
    exp_55_ram[3865] = 52;
    exp_55_ram[3866] = 134;
    exp_55_ram[3867] = 0;
    exp_55_ram[3868] = 7;
    exp_55_ram[3869] = 7;
    exp_55_ram[3870] = 79;
    exp_55_ram[3871] = 5;
    exp_55_ram[3872] = 5;
    exp_55_ram[3873] = 228;
    exp_55_ram[3874] = 244;
    exp_55_ram[3875] = 4;
    exp_55_ram[3876] = 68;
    exp_55_ram[3877] = 52;
    exp_55_ram[3878] = 134;
    exp_55_ram[3879] = 0;
    exp_55_ram[3880] = 7;
    exp_55_ram[3881] = 7;
    exp_55_ram[3882] = 79;
    exp_55_ram[3883] = 5;
    exp_55_ram[3884] = 5;
    exp_55_ram[3885] = 228;
    exp_55_ram[3886] = 244;
    exp_55_ram[3887] = 4;
    exp_55_ram[3888] = 68;
    exp_55_ram[3889] = 52;
    exp_55_ram[3890] = 134;
    exp_55_ram[3891] = 0;
    exp_55_ram[3892] = 7;
    exp_55_ram[3893] = 7;
    exp_55_ram[3894] = 79;
    exp_55_ram[3895] = 5;
    exp_55_ram[3896] = 5;
    exp_55_ram[3897] = 228;
    exp_55_ram[3898] = 244;
    exp_55_ram[3899] = 196;
    exp_55_ram[3900] = 71;
    exp_55_ram[3901] = 244;
    exp_55_ram[3902] = 207;
    exp_55_ram[3903] = 5;
    exp_55_ram[3904] = 5;
    exp_55_ram[3905] = 4;
    exp_55_ram[3906] = 68;
    exp_55_ram[3907] = 166;
    exp_55_ram[3908] = 7;
    exp_55_ram[3909] = 6;
    exp_55_ram[3910] = 182;
    exp_55_ram[3911] = 7;
    exp_55_ram[3912] = 6;
    exp_55_ram[3913] = 0;
    exp_55_ram[3914] = 6;
    exp_55_ram[3915] = 6;
    exp_55_ram[3916] = 0;
    exp_55_ram[3917] = 13;
    exp_55_ram[3918] = 7;
    exp_55_ram[3919] = 198;
    exp_55_ram[3920] = 13;
    exp_55_ram[3921] = 7;
    exp_55_ram[3922] = 214;
    exp_55_ram[3923] = 13;
    exp_55_ram[3924] = 7;
    exp_55_ram[3925] = 215;
    exp_55_ram[3926] = 196;
    exp_55_ram[3927] = 0;
    exp_55_ram[3928] = 199;
    exp_55_ram[3929] = 79;
    exp_55_ram[3930] = 0;
    exp_55_ram[3931] = 193;
    exp_55_ram[3932] = 129;
    exp_55_ram[3933] = 65;
    exp_55_ram[3934] = 1;
    exp_55_ram[3935] = 193;
    exp_55_ram[3936] = 129;
    exp_55_ram[3937] = 65;
    exp_55_ram[3938] = 1;
    exp_55_ram[3939] = 193;
    exp_55_ram[3940] = 129;
    exp_55_ram[3941] = 65;
    exp_55_ram[3942] = 1;
    exp_55_ram[3943] = 1;
    exp_55_ram[3944] = 0;
    exp_55_ram[3945] = 1;
    exp_55_ram[3946] = 17;
    exp_55_ram[3947] = 129;
    exp_55_ram[3948] = 33;
    exp_55_ram[3949] = 49;
    exp_55_ram[3950] = 65;
    exp_55_ram[3951] = 81;
    exp_55_ram[3952] = 1;
    exp_55_ram[3953] = 0;
    exp_55_ram[3954] = 71;
    exp_55_ram[3955] = 207;
    exp_55_ram[3956] = 95;
    exp_55_ram[3957] = 5;
    exp_55_ram[3958] = 71;
    exp_55_ram[3959] = 244;
    exp_55_ram[3960] = 0;
    exp_55_ram[3961] = 199;
    exp_55_ram[3962] = 15;
    exp_55_ram[3963] = 159;
    exp_55_ram[3964] = 5;
    exp_55_ram[3965] = 247;
    exp_55_ram[3966] = 244;
    exp_55_ram[3967] = 0;
    exp_55_ram[3968] = 71;
    exp_55_ram[3969] = 79;
    exp_55_ram[3970] = 223;
    exp_55_ram[3971] = 5;
    exp_55_ram[3972] = 244;
    exp_55_ram[3973] = 0;
    exp_55_ram[3974] = 199;
    exp_55_ram[3975] = 207;
    exp_55_ram[3976] = 95;
    exp_55_ram[3977] = 5;
    exp_55_ram[3978] = 244;
    exp_55_ram[3979] = 0;
    exp_55_ram[3980] = 71;
    exp_55_ram[3981] = 79;
    exp_55_ram[3982] = 207;
    exp_55_ram[3983] = 5;
    exp_55_ram[3984] = 244;
    exp_55_ram[3985] = 112;
    exp_55_ram[3986] = 244;
    exp_55_ram[3987] = 16;
    exp_55_ram[3988] = 244;
    exp_55_ram[3989] = 4;
    exp_55_ram[3990] = 7;
    exp_55_ram[3991] = 31;
    exp_55_ram[3992] = 5;
    exp_55_ram[3993] = 5;
    exp_55_ram[3994] = 228;
    exp_55_ram[3995] = 244;
    exp_55_ram[3996] = 132;
    exp_55_ram[3997] = 196;
    exp_55_ram[3998] = 7;
    exp_55_ram[3999] = 7;
    exp_55_ram[4000] = 95;
    exp_55_ram[4001] = 15;
    exp_55_ram[4002] = 164;
    exp_55_ram[4003] = 180;
    exp_55_ram[4004] = 4;
    exp_55_ram[4005] = 128;
    exp_55_ram[4006] = 0;
    exp_55_ram[4007] = 143;
    exp_55_ram[4008] = 5;
    exp_55_ram[4009] = 5;
    exp_55_ram[4010] = 132;
    exp_55_ram[4011] = 196;
    exp_55_ram[4012] = 7;
    exp_55_ram[4013] = 7;
    exp_55_ram[4014] = 15;
    exp_55_ram[4015] = 5;
    exp_55_ram[4016] = 5;
    exp_55_ram[4017] = 0;
    exp_55_ram[4018] = 7;
    exp_55_ram[4019] = 7;
    exp_55_ram[4020] = 79;
    exp_55_ram[4021] = 5;
    exp_55_ram[4022] = 5;
    exp_55_ram[4023] = 7;
    exp_55_ram[4024] = 7;
    exp_55_ram[4025] = 10;
    exp_55_ram[4026] = 10;
    exp_55_ram[4027] = 79;
    exp_55_ram[4028] = 5;
    exp_55_ram[4029] = 7;
    exp_55_ram[4030] = 0;
    exp_55_ram[4031] = 7;
    exp_55_ram[4032] = 7;
    exp_55_ram[4033] = 0;
    exp_55_ram[4034] = 132;
    exp_55_ram[4035] = 196;
    exp_55_ram[4036] = 38;
    exp_55_ram[4037] = 7;
    exp_55_ram[4038] = 197;
    exp_55_ram[4039] = 54;
    exp_55_ram[4040] = 245;
    exp_55_ram[4041] = 6;
    exp_55_ram[4042] = 228;
    exp_55_ram[4043] = 244;
    exp_55_ram[4044] = 0;
    exp_55_ram[4045] = 223;
    exp_55_ram[4046] = 5;
    exp_55_ram[4047] = 5;
    exp_55_ram[4048] = 228;
    exp_55_ram[4049] = 244;
    exp_55_ram[4050] = 132;
    exp_55_ram[4051] = 7;
    exp_55_ram[4052] = 207;
    exp_55_ram[4053] = 5;
    exp_55_ram[4054] = 7;
    exp_55_ram[4055] = 159;
    exp_55_ram[4056] = 68;
    exp_55_ram[4057] = 23;
    exp_55_ram[4058] = 244;
    exp_55_ram[4059] = 68;
    exp_55_ram[4060] = 48;
    exp_55_ram[4061] = 231;
    exp_55_ram[4062] = 0;
    exp_55_ram[4063] = 0;
    exp_55_ram[4064] = 193;
    exp_55_ram[4065] = 129;
    exp_55_ram[4066] = 65;
    exp_55_ram[4067] = 1;
    exp_55_ram[4068] = 193;
    exp_55_ram[4069] = 129;
    exp_55_ram[4070] = 1;
    exp_55_ram[4071] = 0;
    exp_55_ram[4072] = 1;
    exp_55_ram[4073] = 17;
    exp_55_ram[4074] = 129;
    exp_55_ram[4075] = 1;
    exp_55_ram[4076] = 0;
    exp_55_ram[4077] = 7;
    exp_55_ram[4078] = 31;
    exp_55_ram[4079] = 0;
    exp_55_ram[4080] = 7;
    exp_55_ram[4081] = 95;
    exp_55_ram[4082] = 0;
    exp_55_ram[4083] = 71;
    exp_55_ram[4084] = 159;
    exp_55_ram[4085] = 0;
    exp_55_ram[4086] = 135;
    exp_55_ram[4087] = 223;
    exp_55_ram[4088] = 0;
    exp_55_ram[4089] = 7;
    exp_55_ram[4090] = 31;
    exp_55_ram[4091] = 31;
    exp_55_ram[4092] = 5;
    exp_55_ram[4093] = 244;
    exp_55_ram[4094] = 244;
    exp_55_ram[4095] = 64;
    exp_55_ram[4096] = 231;
    exp_55_ram[4097] = 64;
    exp_55_ram[4098] = 247;
    exp_55_ram[4099] = 48;
    exp_55_ram[4100] = 231;
    exp_55_ram[4101] = 48;
    exp_55_ram[4102] = 247;
    exp_55_ram[4103] = 16;
    exp_55_ram[4104] = 231;
    exp_55_ram[4105] = 32;
    exp_55_ram[4106] = 231;
    exp_55_ram[4107] = 64;
    exp_55_ram[4108] = 79;
    exp_55_ram[4109] = 192;
    exp_55_ram[4110] = 207;
    exp_55_ram[4111] = 64;
    exp_55_ram[4112] = 31;
    exp_55_ram[4113] = 192;
    exp_55_ram[4114] = 223;
    exp_55_ram[4115] = 0;
    exp_55_ram[4116] = 31;
    exp_55_ram[4117] = 5;
    exp_55_ram[4118] = 5;
    exp_55_ram[4119] = 181;
    exp_55_ram[4120] = 1;
    exp_55_ram[4121] = 183;
    exp_55_ram[4122] = 7;
    exp_55_ram[4123] = 5;
    exp_55_ram[4124] = 21;
    exp_55_ram[4125] = 245;
    exp_55_ram[4126] = 1;
    exp_55_ram[4127] = 0;
    exp_55_ram[4128] = 176;
    exp_55_ram[4129] = 245;
    exp_55_ram[4130] = 245;
    exp_55_ram[4131] = 223;
    exp_55_ram[4132] = 250;
    exp_55_ram[4133] = 0;
    exp_55_ram[4134] = 0;
    exp_55_ram[4135] = 0;
    exp_55_ram[4136] = 0;
    exp_55_ram[4137] = 0;
    exp_55_ram[4138] = 0;
    exp_55_ram[4139] = 0;
    exp_55_ram[4140] = 0;
    exp_55_ram[4141] = 0;
    exp_55_ram[4142] = 0;
    exp_55_ram[4143] = 0;
    exp_55_ram[4144] = 0;
    exp_55_ram[4145] = 0;
    exp_55_ram[4146] = 0;
    exp_55_ram[4147] = 0;
    exp_55_ram[4148] = 0;
    exp_55_ram[4149] = 0;
    exp_55_ram[4150] = 0;
    exp_55_ram[4151] = 0;
    exp_55_ram[4152] = 0;
    exp_55_ram[4153] = 0;
    exp_55_ram[4154] = 0;
    exp_55_ram[4155] = 0;
    exp_55_ram[4156] = 0;
    exp_55_ram[4157] = 0;
    exp_55_ram[4158] = 0;
    exp_55_ram[4159] = 0;
    exp_55_ram[4160] = 0;
    exp_55_ram[4161] = 0;
    exp_55_ram[4162] = 0;
    exp_55_ram[4163] = 0;
    exp_55_ram[4164] = 0;
    exp_55_ram[4165] = 0;
    exp_55_ram[4166] = 0;
    exp_55_ram[4167] = 0;
    exp_55_ram[4168] = 0;
    exp_55_ram[4169] = 0;
    exp_55_ram[4170] = 0;
    exp_55_ram[4171] = 0;
    exp_55_ram[4172] = 0;
    exp_55_ram[4173] = 0;
    exp_55_ram[4174] = 0;
    exp_55_ram[4175] = 0;
    exp_55_ram[4176] = 0;
    exp_55_ram[4177] = 0;
    exp_55_ram[4178] = 0;
    exp_55_ram[4179] = 0;
    exp_55_ram[4180] = 0;
    exp_55_ram[4181] = 0;
    exp_55_ram[4182] = 0;
    exp_55_ram[4183] = 0;
    exp_55_ram[4184] = 0;
    exp_55_ram[4185] = 0;
    exp_55_ram[4186] = 0;
    exp_55_ram[4187] = 0;
    exp_55_ram[4188] = 0;
    exp_55_ram[4189] = 0;
    exp_55_ram[4190] = 0;
    exp_55_ram[4191] = 0;
    exp_55_ram[4192] = 0;
    exp_55_ram[4193] = 0;
    exp_55_ram[4194] = 0;
    exp_55_ram[4195] = 0;
    exp_55_ram[4196] = 0;
    exp_55_ram[4197] = 0;
    exp_55_ram[4198] = 0;
    exp_55_ram[4199] = 0;
    exp_55_ram[4200] = 0;
    exp_55_ram[4201] = 0;
    exp_55_ram[4202] = 0;
    exp_55_ram[4203] = 0;
    exp_55_ram[4204] = 0;
    exp_55_ram[4205] = 0;
    exp_55_ram[4206] = 0;
    exp_55_ram[4207] = 0;
    exp_55_ram[4208] = 0;
    exp_55_ram[4209] = 0;
    exp_55_ram[4210] = 0;
    exp_55_ram[4211] = 0;
    exp_55_ram[4212] = 0;
    exp_55_ram[4213] = 0;
    exp_55_ram[4214] = 0;
    exp_55_ram[4215] = 0;
    exp_55_ram[4216] = 0;
    exp_55_ram[4217] = 0;
    exp_55_ram[4218] = 0;
    exp_55_ram[4219] = 0;
    exp_55_ram[4220] = 0;
    exp_55_ram[4221] = 0;
    exp_55_ram[4222] = 0;
    exp_55_ram[4223] = 0;
    exp_55_ram[4224] = 0;
    exp_55_ram[4225] = 0;
    exp_55_ram[4226] = 0;
    exp_55_ram[4227] = 0;
    exp_55_ram[4228] = 0;
    exp_55_ram[4229] = 0;
    exp_55_ram[4230] = 0;
    exp_55_ram[4231] = 0;
    exp_55_ram[4232] = 0;
    exp_55_ram[4233] = 0;
    exp_55_ram[4234] = 0;
    exp_55_ram[4235] = 0;
    exp_55_ram[4236] = 0;
    exp_55_ram[4237] = 0;
    exp_55_ram[4238] = 0;
    exp_55_ram[4239] = 0;
    exp_55_ram[4240] = 0;
    exp_55_ram[4241] = 0;
    exp_55_ram[4242] = 0;
    exp_55_ram[4243] = 0;
    exp_55_ram[4244] = 0;
    exp_55_ram[4245] = 0;
    exp_55_ram[4246] = 0;
    exp_55_ram[4247] = 0;
    exp_55_ram[4248] = 0;
    exp_55_ram[4249] = 0;
    exp_55_ram[4250] = 0;
    exp_55_ram[4251] = 0;
    exp_55_ram[4252] = 0;
    exp_55_ram[4253] = 0;
    exp_55_ram[4254] = 0;
    exp_55_ram[4255] = 0;
    exp_55_ram[4256] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_53) begin
      exp_55_ram[exp_49] <= exp_51;
    end
  end
  assign exp_55 = exp_55_ram[exp_50];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_81) begin
        exp_55_ram[exp_77] <= exp_79;
    end
  end
  assign exp_83 = exp_55_ram[exp_78];
  assign exp_82 = exp_96;
  assign exp_96 = 1;
  assign exp_78 = exp_95;
  assign exp_95 = exp_16[31:2];
  assign exp_81 = exp_92;
  assign exp_92 = 0;
  assign exp_77 = exp_91;
  assign exp_91 = 0;
  assign exp_79 = exp_91;
  assign exp_54 = exp_131;
  assign exp_131 = 1;
  assign exp_50 = exp_130;
  assign exp_130 = exp_18[31:2];
  assign exp_53 = exp_119;
  assign exp_119 = exp_117 & exp_118;
  assign exp_117 = exp_22 & exp_23;
  assign exp_118 = exp_24[2:2];
  assign exp_49 = exp_115;
  assign exp_115 = exp_18[31:2];
  assign exp_51 = exp_116;
  assign exp_116 = exp_19[23:16];

  //Create RAM
  reg [7:0] exp_48_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_48_ram[0] = 0;
    exp_48_ram[1] = 1;
    exp_48_ram[2] = 1;
    exp_48_ram[3] = 2;
    exp_48_ram[4] = 2;
    exp_48_ram[5] = 3;
    exp_48_ram[6] = 3;
    exp_48_ram[7] = 4;
    exp_48_ram[8] = 4;
    exp_48_ram[9] = 5;
    exp_48_ram[10] = 5;
    exp_48_ram[11] = 6;
    exp_48_ram[12] = 6;
    exp_48_ram[13] = 7;
    exp_48_ram[14] = 7;
    exp_48_ram[15] = 8;
    exp_48_ram[16] = 8;
    exp_48_ram[17] = 9;
    exp_48_ram[18] = 9;
    exp_48_ram[19] = 10;
    exp_48_ram[20] = 10;
    exp_48_ram[21] = 11;
    exp_48_ram[22] = 11;
    exp_48_ram[23] = 12;
    exp_48_ram[24] = 12;
    exp_48_ram[25] = 13;
    exp_48_ram[26] = 13;
    exp_48_ram[27] = 14;
    exp_48_ram[28] = 14;
    exp_48_ram[29] = 15;
    exp_48_ram[30] = 15;
    exp_48_ram[31] = 81;
    exp_48_ram[32] = 1;
    exp_48_ram[33] = 48;
    exp_48_ram[34] = 0;
    exp_48_ram[35] = 8;
    exp_48_ram[36] = 135;
    exp_48_ram[37] = 8;
    exp_48_ram[38] = 133;
    exp_48_ram[39] = 131;
    exp_48_ram[40] = 148;
    exp_48_ram[41] = 22;
    exp_48_ram[42] = 134;
    exp_48_ram[43] = 246;
    exp_48_ram[44] = 7;
    exp_48_ram[45] = 120;
    exp_48_ram[46] = 7;
    exp_48_ram[47] = 55;
    exp_48_ram[48] = 23;
    exp_48_ram[49] = 85;
    exp_48_ram[50] = 134;
    exp_48_ram[51] = 198;
    exp_48_ram[52] = 5;
    exp_48_ram[53] = 135;
    exp_48_ram[54] = 6;
    exp_48_ram[55] = 12;
    exp_48_ram[56] = 149;
    exp_48_ram[57] = 215;
    exp_48_ram[58] = 24;
    exp_48_ram[59] = 101;
    exp_48_ram[60] = 147;
    exp_48_ram[61] = 88;
    exp_48_ram[62] = 214;
    exp_48_ram[63] = 22;
    exp_48_ram[64] = 86;
    exp_48_ram[65] = 87;
    exp_48_ram[66] = 247;
    exp_48_ram[67] = 133;
    exp_48_ram[68] = 5;
    exp_48_ram[69] = 23;
    exp_48_ram[70] = 103;
    exp_48_ram[71] = 254;
    exp_48_ram[72] = 135;
    exp_48_ram[73] = 133;
    exp_48_ram[74] = 232;
    exp_48_ram[75] = 246;
    exp_48_ram[76] = 133;
    exp_48_ram[77] = 135;
    exp_48_ram[78] = 135;
    exp_48_ram[79] = 247;
    exp_48_ram[80] = 19;
    exp_48_ram[81] = 83;
    exp_48_ram[82] = 215;
    exp_48_ram[83] = 23;
    exp_48_ram[84] = 99;
    exp_48_ram[85] = 6;
    exp_48_ram[86] = 134;
    exp_48_ram[87] = 124;
    exp_48_ram[88] = 3;
    exp_48_ram[89] = 134;
    exp_48_ram[90] = 102;
    exp_48_ram[91] = 116;
    exp_48_ram[92] = 134;
    exp_48_ram[93] = 21;
    exp_48_ram[94] = 101;
    exp_48_ram[95] = 5;
    exp_48_ram[96] = 0;
    exp_48_ram[97] = 5;
    exp_48_ram[98] = 7;
    exp_48_ram[99] = 108;
    exp_48_ram[100] = 7;
    exp_48_ram[101] = 240;
    exp_48_ram[102] = 22;
    exp_48_ram[103] = 7;
    exp_48_ram[104] = 88;
    exp_48_ram[105] = 7;
    exp_48_ram[106] = 112;
    exp_48_ram[107] = 7;
    exp_48_ram[108] = 116;
    exp_48_ram[109] = 5;
    exp_48_ram[110] = 87;
    exp_48_ram[111] = 134;
    exp_48_ram[112] = 199;
    exp_48_ram[113] = 6;
    exp_48_ram[114] = 7;
    exp_48_ram[115] = 6;
    exp_48_ram[116] = 22;
    exp_48_ram[117] = 135;
    exp_48_ram[118] = 5;
    exp_48_ram[119] = 88;
    exp_48_ram[120] = 22;
    exp_48_ram[121] = 86;
    exp_48_ram[122] = 87;
    exp_48_ram[123] = 246;
    exp_48_ram[124] = 215;
    exp_48_ram[125] = 150;
    exp_48_ram[126] = 231;
    exp_48_ram[127] = 14;
    exp_48_ram[128] = 133;
    exp_48_ram[129] = 126;
    exp_48_ram[130] = 7;
    exp_48_ram[131] = 133;
    exp_48_ram[132] = 104;
    exp_48_ram[133] = 118;
    exp_48_ram[134] = 133;
    exp_48_ram[135] = 7;
    exp_48_ram[136] = 7;
    exp_48_ram[137] = 119;
    exp_48_ram[138] = 19;
    exp_48_ram[139] = 83;
    exp_48_ram[140] = 87;
    exp_48_ram[141] = 151;
    exp_48_ram[142] = 227;
    exp_48_ram[143] = 6;
    exp_48_ram[144] = 6;
    exp_48_ram[145] = 124;
    exp_48_ram[146] = 3;
    exp_48_ram[147] = 6;
    exp_48_ram[148] = 102;
    exp_48_ram[149] = 116;
    exp_48_ram[150] = 6;
    exp_48_ram[151] = 21;
    exp_48_ram[152] = 101;
    exp_48_ram[153] = 128;
    exp_48_ram[154] = 7;
    exp_48_ram[155] = 5;
    exp_48_ram[156] = 100;
    exp_48_ram[157] = 5;
    exp_48_ram[158] = 240;
    exp_48_ram[159] = 24;
    exp_48_ram[160] = 213;
    exp_48_ram[161] = 147;
    exp_48_ram[162] = 151;
    exp_48_ram[163] = 215;
    exp_48_ram[164] = 88;
    exp_48_ram[165] = 102;
    exp_48_ram[166] = 119;
    exp_48_ram[167] = 23;
    exp_48_ram[168] = 215;
    exp_48_ram[169] = 85;
    exp_48_ram[170] = 85;
    exp_48_ram[171] = 23;
    exp_48_ram[172] = 103;
    exp_48_ram[173] = 134;
    exp_48_ram[174] = 5;
    exp_48_ram[175] = 126;
    exp_48_ram[176] = 7;
    exp_48_ram[177] = 5;
    exp_48_ram[178] = 104;
    exp_48_ram[179] = 118;
    exp_48_ram[180] = 5;
    exp_48_ram[181] = 7;
    exp_48_ram[182] = 6;
    exp_48_ram[183] = 247;
    exp_48_ram[184] = 22;
    exp_48_ram[185] = 86;
    exp_48_ram[186] = 214;
    exp_48_ram[187] = 23;
    exp_48_ram[188] = 133;
    exp_48_ram[189] = 103;
    exp_48_ram[190] = 135;
    exp_48_ram[191] = 254;
    exp_48_ram[192] = 135;
    exp_48_ram[193] = 135;
    exp_48_ram[194] = 232;
    exp_48_ram[195] = 246;
    exp_48_ram[196] = 135;
    exp_48_ram[197] = 135;
    exp_48_ram[198] = 149;
    exp_48_ram[199] = 135;
    exp_48_ram[200] = 229;
    exp_48_ram[201] = 240;
    exp_48_ram[202] = 230;
    exp_48_ram[203] = 7;
    exp_48_ram[204] = 244;
    exp_48_ram[205] = 7;
    exp_48_ram[206] = 53;
    exp_48_ram[207] = 149;
    exp_48_ram[208] = 23;
    exp_48_ram[209] = 213;
    exp_48_ram[210] = 7;
    exp_48_ram[211] = 7;
    exp_48_ram[212] = 71;
    exp_48_ram[213] = 5;
    exp_48_ram[214] = 7;
    exp_48_ram[215] = 5;
    exp_48_ram[216] = 22;
    exp_48_ram[217] = 5;
    exp_48_ram[218] = 238;
    exp_48_ram[219] = 181;
    exp_48_ram[220] = 69;
    exp_48_ram[221] = 240;
    exp_48_ram[222] = 7;
    exp_48_ram[223] = 5;
    exp_48_ram[224] = 224;
    exp_48_ram[225] = 5;
    exp_48_ram[226] = 240;
    exp_48_ram[227] = 88;
    exp_48_ram[228] = 150;
    exp_48_ram[229] = 104;
    exp_48_ram[230] = 222;
    exp_48_ram[231] = 94;
    exp_48_ram[232] = 118;
    exp_48_ram[233] = 151;
    exp_48_ram[234] = 215;
    exp_48_ram[235] = 19;
    exp_48_ram[236] = 102;
    exp_48_ram[237] = 23;
    exp_48_ram[238] = 215;
    exp_48_ram[239] = 87;
    exp_48_ram[240] = 94;
    exp_48_ram[241] = 150;
    exp_48_ram[242] = 231;
    exp_48_ram[243] = 143;
    exp_48_ram[244] = 5;
    exp_48_ram[245] = 126;
    exp_48_ram[246] = 7;
    exp_48_ram[247] = 5;
    exp_48_ram[248] = 104;
    exp_48_ram[249] = 118;
    exp_48_ram[250] = 5;
    exp_48_ram[251] = 7;
    exp_48_ram[252] = 7;
    exp_48_ram[253] = 118;
    exp_48_ram[254] = 87;
    exp_48_ram[255] = 150;
    exp_48_ram[256] = 142;
    exp_48_ram[257] = 23;
    exp_48_ram[258] = 215;
    exp_48_ram[259] = 231;
    exp_48_ram[260] = 6;
    exp_48_ram[261] = 254;
    exp_48_ram[262] = 135;
    exp_48_ram[263] = 6;
    exp_48_ram[264] = 232;
    exp_48_ram[265] = 246;
    exp_48_ram[266] = 6;
    exp_48_ram[267] = 135;
    exp_48_ram[268] = 21;
    exp_48_ram[269] = 14;
    exp_48_ram[270] = 101;
    exp_48_ram[271] = 134;
    exp_48_ram[272] = 120;
    exp_48_ram[273] = 86;
    exp_48_ram[274] = 118;
    exp_48_ram[275] = 83;
    exp_48_ram[276] = 135;
    exp_48_ram[277] = 14;
    exp_48_ram[278] = 6;
    exp_48_ram[279] = 87;
    exp_48_ram[280] = 8;
    exp_48_ram[281] = 8;
    exp_48_ram[282] = 7;
    exp_48_ram[283] = 6;
    exp_48_ram[284] = 116;
    exp_48_ram[285] = 6;
    exp_48_ram[286] = 86;
    exp_48_ram[287] = 134;
    exp_48_ram[288] = 230;
    exp_48_ram[289] = 156;
    exp_48_ram[290] = 7;
    exp_48_ram[291] = 135;
    exp_48_ram[292] = 119;
    exp_48_ram[293] = 23;
    exp_48_ram[294] = 126;
    exp_48_ram[295] = 152;
    exp_48_ram[296] = 7;
    exp_48_ram[297] = 5;
    exp_48_ram[298] = 254;
    exp_48_ram[299] = 5;
    exp_48_ram[300] = 240;
    exp_48_ram[301] = 5;
    exp_48_ram[302] = 5;
    exp_48_ram[303] = 240;
    exp_48_ram[304] = 7;
    exp_48_ram[305] = 7;
    exp_48_ram[306] = 216;
    exp_48_ram[307] = 120;
    exp_48_ram[308] = 7;
    exp_48_ram[309] = 3;
    exp_48_ram[310] = 120;
    exp_48_ram[311] = 213;
    exp_48_ram[312] = 14;
    exp_48_ram[313] = 213;
    exp_48_ram[314] = 119;
    exp_48_ram[315] = 14;
    exp_48_ram[316] = 245;
    exp_48_ram[317] = 214;
    exp_48_ram[318] = 26;
    exp_48_ram[319] = 238;
    exp_48_ram[320] = 138;
    exp_48_ram[321] = 5;
    exp_48_ram[322] = 128;
    exp_48_ram[323] = 150;
    exp_48_ram[324] = 110;
    exp_48_ram[325] = 152;
    exp_48_ram[326] = 16;
    exp_48_ram[327] = 231;
    exp_48_ram[328] = 183;
    exp_48_ram[329] = 150;
    exp_48_ram[330] = 102;
    exp_48_ram[331] = 12;
    exp_48_ram[332] = 156;
    exp_48_ram[333] = 20;
    exp_48_ram[334] = 208;
    exp_48_ram[335] = 0;
    exp_48_ram[336] = 5;
    exp_48_ram[337] = 128;
    exp_48_ram[338] = 5;
    exp_48_ram[339] = 138;
    exp_48_ram[340] = 133;
    exp_48_ram[341] = 128;
    exp_48_ram[342] = 86;
    exp_48_ram[343] = 2;
    exp_48_ram[344] = 128;
    exp_48_ram[345] = 108;
    exp_48_ram[346] = 146;
    exp_48_ram[347] = 104;
    exp_48_ram[348] = 102;
    exp_48_ram[349] = 5;
    exp_48_ram[350] = 128;
    exp_48_ram[351] = 5;
    exp_48_ram[352] = 128;
    exp_48_ram[353] = 152;
    exp_48_ram[354] = 240;
    exp_48_ram[355] = 232;
    exp_48_ram[356] = 240;
    exp_48_ram[357] = 142;
    exp_48_ram[358] = 158;
    exp_48_ram[359] = 7;
    exp_48_ram[360] = 240;
    exp_48_ram[361] = 1;
    exp_48_ram[362] = 36;
    exp_48_ram[363] = 38;
    exp_48_ram[364] = 4;
    exp_48_ram[365] = 2;
    exp_48_ram[366] = 0;
    exp_48_ram[367] = 7;
    exp_48_ram[368] = 7;
    exp_48_ram[369] = 7;
    exp_48_ram[370] = 192;
    exp_48_ram[371] = 7;
    exp_48_ram[372] = 135;
    exp_48_ram[373] = 5;
    exp_48_ram[374] = 87;
    exp_48_ram[375] = 20;
    exp_48_ram[376] = 32;
    exp_48_ram[377] = 5;
    exp_48_ram[378] = 151;
    exp_48_ram[379] = 36;
    exp_48_ram[380] = 23;
    exp_48_ram[381] = 215;
    exp_48_ram[382] = 102;
    exp_48_ram[383] = 133;
    exp_48_ram[384] = 1;
    exp_48_ram[385] = 128;
    exp_48_ram[386] = 7;
    exp_48_ram[387] = 23;
    exp_48_ram[388] = 4;
    exp_48_ram[389] = 240;
    exp_48_ram[390] = 7;
    exp_48_ram[391] = 7;
    exp_48_ram[392] = 240;
    exp_48_ram[393] = 1;
    exp_48_ram[394] = 46;
    exp_48_ram[395] = 44;
    exp_48_ram[396] = 42;
    exp_48_ram[397] = 40;
    exp_48_ram[398] = 38;
    exp_48_ram[399] = 36;
    exp_48_ram[400] = 103;
    exp_48_ram[401] = 140;
    exp_48_ram[402] = 4;
    exp_48_ram[403] = 137;
    exp_48_ram[404] = 132;
    exp_48_ram[405] = 132;
    exp_48_ram[406] = 133;
    exp_48_ram[407] = 0;
    exp_48_ram[408] = 9;
    exp_48_ram[409] = 10;
    exp_48_ram[410] = 10;
    exp_48_ram[411] = 7;
    exp_48_ram[412] = 196;
    exp_48_ram[413] = 7;
    exp_48_ram[414] = 7;
    exp_48_ram[415] = 84;
    exp_48_ram[416] = 7;
    exp_48_ram[417] = 66;
    exp_48_ram[418] = 4;
    exp_48_ram[419] = 135;
    exp_48_ram[420] = 132;
    exp_48_ram[421] = 84;
    exp_48_ram[422] = 21;
    exp_48_ram[423] = 228;
    exp_48_ram[424] = 23;
    exp_48_ram[425] = 32;
    exp_48_ram[426] = 36;
    exp_48_ram[427] = 149;
    exp_48_ram[428] = 26;
    exp_48_ram[429] = 213;
    exp_48_ram[430] = 103;
    exp_48_ram[431] = 36;
    exp_48_ram[432] = 41;
    exp_48_ram[433] = 41;
    exp_48_ram[434] = 42;
    exp_48_ram[435] = 133;
    exp_48_ram[436] = 5;
    exp_48_ram[437] = 1;
    exp_48_ram[438] = 128;
    exp_48_ram[439] = 0;
    exp_48_ram[440] = 9;
    exp_48_ram[441] = 240;
    exp_48_ram[442] = 133;
    exp_48_ram[443] = 20;
    exp_48_ram[444] = 7;
    exp_48_ram[445] = 240;
    exp_48_ram[446] = 7;
    exp_48_ram[447] = 220;
    exp_48_ram[448] = 134;
    exp_48_ram[449] = 5;
    exp_48_ram[450] = 5;
    exp_48_ram[451] = 0;
    exp_48_ram[452] = 101;
    exp_48_ram[453] = 6;
    exp_48_ram[454] = 52;
    exp_48_ram[455] = 5;
    exp_48_ram[456] = 5;
    exp_48_ram[457] = 6;
    exp_48_ram[458] = 0;
    exp_48_ram[459] = 228;
    exp_48_ram[460] = 137;
    exp_48_ram[461] = 7;
    exp_48_ram[462] = 7;
    exp_48_ram[463] = 5;
    exp_48_ram[464] = 84;
    exp_48_ram[465] = 7;
    exp_48_ram[466] = 66;
    exp_48_ram[467] = 135;
    exp_48_ram[468] = 21;
    exp_48_ram[469] = 9;
    exp_48_ram[470] = 9;
    exp_48_ram[471] = 89;
    exp_48_ram[472] = 101;
    exp_48_ram[473] = 23;
    exp_48_ram[474] = 7;
    exp_48_ram[475] = 7;
    exp_48_ram[476] = 245;
    exp_48_ram[477] = 247;
    exp_48_ram[478] = 0;
    exp_48_ram[479] = 247;
    exp_48_ram[480] = 6;
    exp_48_ram[481] = 10;
    exp_48_ram[482] = 135;
    exp_48_ram[483] = 55;
    exp_48_ram[484] = 133;
    exp_48_ram[485] = 7;
    exp_48_ram[486] = 7;
    exp_48_ram[487] = 247;
    exp_48_ram[488] = 12;
    exp_48_ram[489] = 7;
    exp_48_ram[490] = 7;
    exp_48_ram[491] = 10;
    exp_48_ram[492] = 245;
    exp_48_ram[493] = 10;
    exp_48_ram[494] = 215;
    exp_48_ram[495] = 149;
    exp_48_ram[496] = 103;
    exp_48_ram[497] = 212;
    exp_48_ram[498] = 240;
    exp_48_ram[499] = 133;
    exp_48_ram[500] = 21;
    exp_48_ram[501] = 7;
    exp_48_ram[502] = 240;
    exp_48_ram[503] = 4;
    exp_48_ram[504] = 7;
    exp_48_ram[505] = 10;
    exp_48_ram[506] = 240;
    exp_48_ram[507] = 0;
    exp_48_ram[508] = 7;
    exp_48_ram[509] = 135;
    exp_48_ram[510] = 76;
    exp_48_ram[511] = 5;
    exp_48_ram[512] = 7;
    exp_48_ram[513] = 213;
    exp_48_ram[514] = 5;
    exp_48_ram[515] = 128;
    exp_48_ram[516] = 215;
    exp_48_ram[517] = 85;
    exp_48_ram[518] = 149;
    exp_48_ram[519] = 101;
    exp_48_ram[520] = 240;
    exp_48_ram[521] = 0;
    exp_48_ram[522] = 7;
    exp_48_ram[523] = 135;
    exp_48_ram[524] = 76;
    exp_48_ram[525] = 5;
    exp_48_ram[526] = 7;
    exp_48_ram[527] = 21;
    exp_48_ram[528] = 5;
    exp_48_ram[529] = 128;
    exp_48_ram[530] = 23;
    exp_48_ram[531] = 149;
    exp_48_ram[532] = 85;
    exp_48_ram[533] = 229;
    exp_48_ram[534] = 240;
    exp_48_ram[535] = 7;
    exp_48_ram[536] = 122;
    exp_48_ram[537] = 7;
    exp_48_ram[538] = 183;
    exp_48_ram[539] = 151;
    exp_48_ram[540] = 23;
    exp_48_ram[541] = 6;
    exp_48_ram[542] = 134;
    exp_48_ram[543] = 85;
    exp_48_ram[544] = 7;
    exp_48_ram[545] = 133;
    exp_48_ram[546] = 69;
    exp_48_ram[547] = 133;
    exp_48_ram[548] = 128;
    exp_48_ram[549] = 7;
    exp_48_ram[550] = 7;
    exp_48_ram[551] = 106;
    exp_48_ram[552] = 7;
    exp_48_ram[553] = 240;
    exp_48_ram[554] = 117;
    exp_48_ram[555] = 110;
    exp_48_ram[556] = 87;
    exp_48_ram[557] = 104;
    exp_48_ram[558] = 105;
    exp_48_ram[559] = 0;
    exp_48_ram[560] = 97;
    exp_48_ram[561] = 98;
    exp_48_ram[562] = 65;
    exp_48_ram[563] = 97;
    exp_48_ram[564] = 110;
    exp_48_ram[565] = 65;
    exp_48_ram[566] = 101;
    exp_48_ram[567] = 116;
    exp_48_ram[568] = 68;
    exp_48_ram[569] = 0;
    exp_48_ram[570] = 101;
    exp_48_ram[571] = 32;
    exp_48_ram[572] = 108;
    exp_48_ram[573] = 0;
    exp_48_ram[574] = 117;
    exp_48_ram[575] = 110;
    exp_48_ram[576] = 110;
    exp_48_ram[577] = 116;
    exp_48_ram[578] = 100;
    exp_48_ram[579] = 100;
    exp_48_ram[580] = 46;
    exp_48_ram[581] = 0;
    exp_48_ram[582] = 117;
    exp_48_ram[583] = 117;
    exp_48_ram[584] = 45;
    exp_48_ram[585] = 32;
    exp_48_ram[586] = 101;
    exp_48_ram[587] = 32;
    exp_48_ram[588] = 116;
    exp_48_ram[589] = 105;
    exp_48_ram[590] = 105;
    exp_48_ram[591] = 32;
    exp_48_ram[592] = 111;
    exp_48_ram[593] = 0;
    exp_48_ram[594] = 117;
    exp_48_ram[595] = 45;
    exp_48_ram[596] = 32;
    exp_48_ram[597] = 101;
    exp_48_ram[598] = 32;
    exp_48_ram[599] = 116;
    exp_48_ram[600] = 105;
    exp_48_ram[601] = 105;
    exp_48_ram[602] = 32;
    exp_48_ram[603] = 111;
    exp_48_ram[604] = 0;
    exp_48_ram[605] = 117;
    exp_48_ram[606] = 45;
    exp_48_ram[607] = 32;
    exp_48_ram[608] = 101;
    exp_48_ram[609] = 32;
    exp_48_ram[610] = 105;
    exp_48_ram[611] = 32;
    exp_48_ram[612] = 49;
    exp_48_ram[613] = 99;
    exp_48_ram[614] = 10;
    exp_48_ram[615] = 117;
    exp_48_ram[616] = 45;
    exp_48_ram[617] = 32;
    exp_48_ram[618] = 101;
    exp_48_ram[619] = 32;
    exp_48_ram[620] = 105;
    exp_48_ram[621] = 32;
    exp_48_ram[622] = 49;
    exp_48_ram[623] = 99;
    exp_48_ram[624] = 10;
    exp_48_ram[625] = 101;
    exp_48_ram[626] = 10;
    exp_48_ram[627] = 111;
    exp_48_ram[628] = 58;
    exp_48_ram[629] = 97;
    exp_48_ram[630] = 0;
    exp_48_ram[631] = 111;
    exp_48_ram[632] = 10;
    exp_48_ram[633] = 105;
    exp_48_ram[634] = 101;
    exp_48_ram[635] = 0;
    exp_48_ram[636] = 67;
    exp_48_ram[637] = 115;
    exp_48_ram[638] = 68;
    exp_48_ram[639] = 10;
    exp_48_ram[640] = 97;
    exp_48_ram[641] = 101;
    exp_48_ram[642] = 32;
    exp_48_ram[643] = 108;
    exp_48_ram[644] = 0;
    exp_48_ram[645] = 41;
    exp_48_ram[646] = 105;
    exp_48_ram[647] = 32;
    exp_48_ram[648] = 101;
    exp_48_ram[649] = 0;
    exp_48_ram[650] = 41;
    exp_48_ram[651] = 115;
    exp_48_ram[652] = 117;
    exp_48_ram[653] = 112;
    exp_48_ram[654] = 97;
    exp_48_ram[655] = 110;
    exp_48_ram[656] = 41;
    exp_48_ram[657] = 108;
    exp_48_ram[658] = 108;
    exp_48_ram[659] = 10;
    exp_48_ram[660] = 1;
    exp_48_ram[661] = 3;
    exp_48_ram[662] = 4;
    exp_48_ram[663] = 4;
    exp_48_ram[664] = 5;
    exp_48_ram[665] = 5;
    exp_48_ram[666] = 5;
    exp_48_ram[667] = 5;
    exp_48_ram[668] = 6;
    exp_48_ram[669] = 6;
    exp_48_ram[670] = 6;
    exp_48_ram[671] = 6;
    exp_48_ram[672] = 6;
    exp_48_ram[673] = 6;
    exp_48_ram[674] = 6;
    exp_48_ram[675] = 6;
    exp_48_ram[676] = 7;
    exp_48_ram[677] = 7;
    exp_48_ram[678] = 7;
    exp_48_ram[679] = 7;
    exp_48_ram[680] = 7;
    exp_48_ram[681] = 7;
    exp_48_ram[682] = 7;
    exp_48_ram[683] = 7;
    exp_48_ram[684] = 7;
    exp_48_ram[685] = 7;
    exp_48_ram[686] = 7;
    exp_48_ram[687] = 7;
    exp_48_ram[688] = 7;
    exp_48_ram[689] = 7;
    exp_48_ram[690] = 7;
    exp_48_ram[691] = 7;
    exp_48_ram[692] = 8;
    exp_48_ram[693] = 8;
    exp_48_ram[694] = 8;
    exp_48_ram[695] = 8;
    exp_48_ram[696] = 8;
    exp_48_ram[697] = 8;
    exp_48_ram[698] = 8;
    exp_48_ram[699] = 8;
    exp_48_ram[700] = 8;
    exp_48_ram[701] = 8;
    exp_48_ram[702] = 8;
    exp_48_ram[703] = 8;
    exp_48_ram[704] = 8;
    exp_48_ram[705] = 8;
    exp_48_ram[706] = 8;
    exp_48_ram[707] = 8;
    exp_48_ram[708] = 8;
    exp_48_ram[709] = 8;
    exp_48_ram[710] = 8;
    exp_48_ram[711] = 8;
    exp_48_ram[712] = 8;
    exp_48_ram[713] = 8;
    exp_48_ram[714] = 8;
    exp_48_ram[715] = 8;
    exp_48_ram[716] = 8;
    exp_48_ram[717] = 8;
    exp_48_ram[718] = 8;
    exp_48_ram[719] = 8;
    exp_48_ram[720] = 8;
    exp_48_ram[721] = 8;
    exp_48_ram[722] = 8;
    exp_48_ram[723] = 8;
    exp_48_ram[724] = 1;
    exp_48_ram[725] = 38;
    exp_48_ram[726] = 4;
    exp_48_ram[727] = 46;
    exp_48_ram[728] = 39;
    exp_48_ram[729] = 38;
    exp_48_ram[730] = 39;
    exp_48_ram[731] = 167;
    exp_48_ram[732] = 133;
    exp_48_ram[733] = 36;
    exp_48_ram[734] = 1;
    exp_48_ram[735] = 128;
    exp_48_ram[736] = 1;
    exp_48_ram[737] = 38;
    exp_48_ram[738] = 4;
    exp_48_ram[739] = 46;
    exp_48_ram[740] = 44;
    exp_48_ram[741] = 39;
    exp_48_ram[742] = 38;
    exp_48_ram[743] = 39;
    exp_48_ram[744] = 39;
    exp_48_ram[745] = 160;
    exp_48_ram[746] = 39;
    exp_48_ram[747] = 133;
    exp_48_ram[748] = 36;
    exp_48_ram[749] = 1;
    exp_48_ram[750] = 128;
    exp_48_ram[751] = 1;
    exp_48_ram[752] = 38;
    exp_48_ram[753] = 36;
    exp_48_ram[754] = 4;
    exp_48_ram[755] = 71;
    exp_48_ram[756] = 167;
    exp_48_ram[757] = 133;
    exp_48_ram[758] = 240;
    exp_48_ram[759] = 7;
    exp_48_ram[760] = 133;
    exp_48_ram[761] = 32;
    exp_48_ram[762] = 36;
    exp_48_ram[763] = 1;
    exp_48_ram[764] = 128;
    exp_48_ram[765] = 1;
    exp_48_ram[766] = 38;
    exp_48_ram[767] = 36;
    exp_48_ram[768] = 4;
    exp_48_ram[769] = 46;
    exp_48_ram[770] = 44;
    exp_48_ram[771] = 38;
    exp_48_ram[772] = 0;
    exp_48_ram[773] = 39;
    exp_48_ram[774] = 135;
    exp_48_ram[775] = 38;
    exp_48_ram[776] = 39;
    exp_48_ram[777] = 7;
    exp_48_ram[778] = 199;
    exp_48_ram[779] = 37;
    exp_48_ram[780] = 133;
    exp_48_ram[781] = 240;
    exp_48_ram[782] = 39;
    exp_48_ram[783] = 39;
    exp_48_ram[784] = 7;
    exp_48_ram[785] = 199;
    exp_48_ram[786] = 150;
    exp_48_ram[787] = 39;
    exp_48_ram[788] = 133;
    exp_48_ram[789] = 32;
    exp_48_ram[790] = 36;
    exp_48_ram[791] = 1;
    exp_48_ram[792] = 128;
    exp_48_ram[793] = 1;
    exp_48_ram[794] = 46;
    exp_48_ram[795] = 44;
    exp_48_ram[796] = 4;
    exp_48_ram[797] = 38;
    exp_48_ram[798] = 71;
    exp_48_ram[799] = 167;
    exp_48_ram[800] = 133;
    exp_48_ram[801] = 37;
    exp_48_ram[802] = 240;
    exp_48_ram[803] = 71;
    exp_48_ram[804] = 167;
    exp_48_ram[805] = 133;
    exp_48_ram[806] = 5;
    exp_48_ram[807] = 240;
    exp_48_ram[808] = 7;
    exp_48_ram[809] = 133;
    exp_48_ram[810] = 32;
    exp_48_ram[811] = 36;
    exp_48_ram[812] = 1;
    exp_48_ram[813] = 128;
    exp_48_ram[814] = 1;
    exp_48_ram[815] = 46;
    exp_48_ram[816] = 4;
    exp_48_ram[817] = 7;
    exp_48_ram[818] = 36;
    exp_48_ram[819] = 34;
    exp_48_ram[820] = 32;
    exp_48_ram[821] = 7;
    exp_48_ram[822] = 0;
    exp_48_ram[823] = 36;
    exp_48_ram[824] = 1;
    exp_48_ram[825] = 128;
    exp_48_ram[826] = 1;
    exp_48_ram[827] = 46;
    exp_48_ram[828] = 44;
    exp_48_ram[829] = 4;
    exp_48_ram[830] = 7;
    exp_48_ram[831] = 36;
    exp_48_ram[832] = 34;
    exp_48_ram[833] = 32;
    exp_48_ram[834] = 7;
    exp_48_ram[835] = 71;
    exp_48_ram[836] = 136;
    exp_48_ram[837] = 71;
    exp_48_ram[838] = 133;
    exp_48_ram[839] = 16;
    exp_48_ram[840] = 0;
    exp_48_ram[841] = 32;
    exp_48_ram[842] = 36;
    exp_48_ram[843] = 1;
    exp_48_ram[844] = 128;
    exp_48_ram[845] = 1;
    exp_48_ram[846] = 38;
    exp_48_ram[847] = 4;
    exp_48_ram[848] = 46;
    exp_48_ram[849] = 44;
    exp_48_ram[850] = 39;
    exp_48_ram[851] = 38;
    exp_48_ram[852] = 0;
    exp_48_ram[853] = 39;
    exp_48_ram[854] = 135;
    exp_48_ram[855] = 38;
    exp_48_ram[856] = 39;
    exp_48_ram[857] = 199;
    exp_48_ram[858] = 138;
    exp_48_ram[859] = 39;
    exp_48_ram[860] = 135;
    exp_48_ram[861] = 44;
    exp_48_ram[862] = 158;
    exp_48_ram[863] = 39;
    exp_48_ram[864] = 39;
    exp_48_ram[865] = 7;
    exp_48_ram[866] = 133;
    exp_48_ram[867] = 36;
    exp_48_ram[868] = 1;
    exp_48_ram[869] = 128;
    exp_48_ram[870] = 1;
    exp_48_ram[871] = 46;
    exp_48_ram[872] = 4;
    exp_48_ram[873] = 7;
    exp_48_ram[874] = 7;
    exp_48_ram[875] = 71;
    exp_48_ram[876] = 7;
    exp_48_ram[877] = 252;
    exp_48_ram[878] = 71;
    exp_48_ram[879] = 7;
    exp_48_ram[880] = 230;
    exp_48_ram[881] = 7;
    exp_48_ram[882] = 0;
    exp_48_ram[883] = 7;
    exp_48_ram[884] = 247;
    exp_48_ram[885] = 247;
    exp_48_ram[886] = 133;
    exp_48_ram[887] = 36;
    exp_48_ram[888] = 1;
    exp_48_ram[889] = 128;
    exp_48_ram[890] = 1;
    exp_48_ram[891] = 38;
    exp_48_ram[892] = 36;
    exp_48_ram[893] = 4;
    exp_48_ram[894] = 46;
    exp_48_ram[895] = 38;
    exp_48_ram[896] = 0;
    exp_48_ram[897] = 39;
    exp_48_ram[898] = 7;
    exp_48_ram[899] = 151;
    exp_48_ram[900] = 135;
    exp_48_ram[901] = 151;
    exp_48_ram[902] = 134;
    exp_48_ram[903] = 39;
    exp_48_ram[904] = 167;
    exp_48_ram[905] = 134;
    exp_48_ram[906] = 39;
    exp_48_ram[907] = 32;
    exp_48_ram[908] = 199;
    exp_48_ram[909] = 7;
    exp_48_ram[910] = 135;
    exp_48_ram[911] = 38;
    exp_48_ram[912] = 39;
    exp_48_ram[913] = 167;
    exp_48_ram[914] = 199;
    exp_48_ram[915] = 133;
    exp_48_ram[916] = 240;
    exp_48_ram[917] = 7;
    exp_48_ram[918] = 150;
    exp_48_ram[919] = 39;
    exp_48_ram[920] = 133;
    exp_48_ram[921] = 32;
    exp_48_ram[922] = 36;
    exp_48_ram[923] = 1;
    exp_48_ram[924] = 128;
    exp_48_ram[925] = 1;
    exp_48_ram[926] = 46;
    exp_48_ram[927] = 44;
    exp_48_ram[928] = 4;
    exp_48_ram[929] = 46;
    exp_48_ram[930] = 44;
    exp_48_ram[931] = 42;
    exp_48_ram[932] = 40;
    exp_48_ram[933] = 38;
    exp_48_ram[934] = 36;
    exp_48_ram[935] = 34;
    exp_48_ram[936] = 32;
    exp_48_ram[937] = 39;
    exp_48_ram[938] = 36;
    exp_48_ram[939] = 39;
    exp_48_ram[940] = 247;
    exp_48_ram[941] = 156;
    exp_48_ram[942] = 39;
    exp_48_ram[943] = 247;
    exp_48_ram[944] = 150;
    exp_48_ram[945] = 39;
    exp_48_ram[946] = 38;
    exp_48_ram[947] = 0;
    exp_48_ram[948] = 39;
    exp_48_ram[949] = 135;
    exp_48_ram[950] = 42;
    exp_48_ram[951] = 39;
    exp_48_ram[952] = 38;
    exp_48_ram[953] = 134;
    exp_48_ram[954] = 37;
    exp_48_ram[955] = 5;
    exp_48_ram[956] = 0;
    exp_48_ram[957] = 39;
    exp_48_ram[958] = 135;
    exp_48_ram[959] = 38;
    exp_48_ram[960] = 39;
    exp_48_ram[961] = 39;
    exp_48_ram[962] = 100;
    exp_48_ram[963] = 0;
    exp_48_ram[964] = 39;
    exp_48_ram[965] = 135;
    exp_48_ram[966] = 36;
    exp_48_ram[967] = 39;
    exp_48_ram[968] = 39;
    exp_48_ram[969] = 7;
    exp_48_ram[970] = 197;
    exp_48_ram[971] = 39;
    exp_48_ram[972] = 135;
    exp_48_ram[973] = 42;
    exp_48_ram[974] = 39;
    exp_48_ram[975] = 38;
    exp_48_ram[976] = 134;
    exp_48_ram[977] = 37;
    exp_48_ram[978] = 0;
    exp_48_ram[979] = 39;
    exp_48_ram[980] = 144;
    exp_48_ram[981] = 39;
    exp_48_ram[982] = 247;
    exp_48_ram[983] = 128;
    exp_48_ram[984] = 0;
    exp_48_ram[985] = 39;
    exp_48_ram[986] = 135;
    exp_48_ram[987] = 42;
    exp_48_ram[988] = 39;
    exp_48_ram[989] = 38;
    exp_48_ram[990] = 134;
    exp_48_ram[991] = 37;
    exp_48_ram[992] = 5;
    exp_48_ram[993] = 0;
    exp_48_ram[994] = 39;
    exp_48_ram[995] = 39;
    exp_48_ram[996] = 7;
    exp_48_ram[997] = 39;
    exp_48_ram[998] = 230;
    exp_48_ram[999] = 39;
    exp_48_ram[1000] = 133;
    exp_48_ram[1001] = 32;
    exp_48_ram[1002] = 36;
    exp_48_ram[1003] = 1;
    exp_48_ram[1004] = 128;
    exp_48_ram[1005] = 1;
    exp_48_ram[1006] = 38;
    exp_48_ram[1007] = 36;
    exp_48_ram[1008] = 4;
    exp_48_ram[1009] = 38;
    exp_48_ram[1010] = 36;
    exp_48_ram[1011] = 34;
    exp_48_ram[1012] = 32;
    exp_48_ram[1013] = 46;
    exp_48_ram[1014] = 44;
    exp_48_ram[1015] = 7;
    exp_48_ram[1016] = 40;
    exp_48_ram[1017] = 11;
    exp_48_ram[1018] = 39;
    exp_48_ram[1019] = 247;
    exp_48_ram[1020] = 154;
    exp_48_ram[1021] = 39;
    exp_48_ram[1022] = 136;
    exp_48_ram[1023] = 39;
    exp_48_ram[1024] = 247;
    exp_48_ram[1025] = 130;
    exp_48_ram[1026] = 71;
    exp_48_ram[1027] = 152;
    exp_48_ram[1028] = 39;
    exp_48_ram[1029] = 247;
    exp_48_ram[1030] = 136;
    exp_48_ram[1031] = 39;
    exp_48_ram[1032] = 135;
    exp_48_ram[1033] = 34;
    exp_48_ram[1034] = 0;
    exp_48_ram[1035] = 39;
    exp_48_ram[1036] = 135;
    exp_48_ram[1037] = 44;
    exp_48_ram[1038] = 39;
    exp_48_ram[1039] = 7;
    exp_48_ram[1040] = 7;
    exp_48_ram[1041] = 128;
    exp_48_ram[1042] = 39;
    exp_48_ram[1043] = 39;
    exp_48_ram[1044] = 120;
    exp_48_ram[1045] = 39;
    exp_48_ram[1046] = 7;
    exp_48_ram[1047] = 248;
    exp_48_ram[1048] = 0;
    exp_48_ram[1049] = 39;
    exp_48_ram[1050] = 135;
    exp_48_ram[1051] = 44;
    exp_48_ram[1052] = 39;
    exp_48_ram[1053] = 7;
    exp_48_ram[1054] = 7;
    exp_48_ram[1055] = 128;
    exp_48_ram[1056] = 39;
    exp_48_ram[1057] = 247;
    exp_48_ram[1058] = 142;
    exp_48_ram[1059] = 39;
    exp_48_ram[1060] = 39;
    exp_48_ram[1061] = 120;
    exp_48_ram[1062] = 39;
    exp_48_ram[1063] = 7;
    exp_48_ram[1064] = 242;
    exp_48_ram[1065] = 39;
    exp_48_ram[1066] = 247;
    exp_48_ram[1067] = 128;
    exp_48_ram[1068] = 39;
    exp_48_ram[1069] = 247;
    exp_48_ram[1070] = 152;
    exp_48_ram[1071] = 39;
    exp_48_ram[1072] = 132;
    exp_48_ram[1073] = 39;
    exp_48_ram[1074] = 39;
    exp_48_ram[1075] = 8;
    exp_48_ram[1076] = 39;
    exp_48_ram[1077] = 39;
    exp_48_ram[1078] = 24;
    exp_48_ram[1079] = 39;
    exp_48_ram[1080] = 135;
    exp_48_ram[1081] = 44;
    exp_48_ram[1082] = 39;
    exp_48_ram[1083] = 142;
    exp_48_ram[1084] = 39;
    exp_48_ram[1085] = 7;
    exp_48_ram[1086] = 24;
    exp_48_ram[1087] = 39;
    exp_48_ram[1088] = 135;
    exp_48_ram[1089] = 44;
    exp_48_ram[1090] = 39;
    exp_48_ram[1091] = 7;
    exp_48_ram[1092] = 30;
    exp_48_ram[1093] = 39;
    exp_48_ram[1094] = 247;
    exp_48_ram[1095] = 152;
    exp_48_ram[1096] = 39;
    exp_48_ram[1097] = 7;
    exp_48_ram[1098] = 226;
    exp_48_ram[1099] = 39;
    exp_48_ram[1100] = 135;
    exp_48_ram[1101] = 44;
    exp_48_ram[1102] = 39;
    exp_48_ram[1103] = 7;
    exp_48_ram[1104] = 7;
    exp_48_ram[1105] = 128;
    exp_48_ram[1106] = 0;
    exp_48_ram[1107] = 39;
    exp_48_ram[1108] = 7;
    exp_48_ram[1109] = 30;
    exp_48_ram[1110] = 39;
    exp_48_ram[1111] = 247;
    exp_48_ram[1112] = 136;
    exp_48_ram[1113] = 39;
    exp_48_ram[1114] = 7;
    exp_48_ram[1115] = 226;
    exp_48_ram[1116] = 39;
    exp_48_ram[1117] = 135;
    exp_48_ram[1118] = 44;
    exp_48_ram[1119] = 39;
    exp_48_ram[1120] = 7;
    exp_48_ram[1121] = 7;
    exp_48_ram[1122] = 128;
    exp_48_ram[1123] = 0;
    exp_48_ram[1124] = 39;
    exp_48_ram[1125] = 7;
    exp_48_ram[1126] = 22;
    exp_48_ram[1127] = 39;
    exp_48_ram[1128] = 7;
    exp_48_ram[1129] = 224;
    exp_48_ram[1130] = 39;
    exp_48_ram[1131] = 135;
    exp_48_ram[1132] = 44;
    exp_48_ram[1133] = 39;
    exp_48_ram[1134] = 7;
    exp_48_ram[1135] = 7;
    exp_48_ram[1136] = 128;
    exp_48_ram[1137] = 39;
    exp_48_ram[1138] = 7;
    exp_48_ram[1139] = 224;
    exp_48_ram[1140] = 39;
    exp_48_ram[1141] = 135;
    exp_48_ram[1142] = 44;
    exp_48_ram[1143] = 39;
    exp_48_ram[1144] = 7;
    exp_48_ram[1145] = 7;
    exp_48_ram[1146] = 128;
    exp_48_ram[1147] = 39;
    exp_48_ram[1148] = 7;
    exp_48_ram[1149] = 224;
    exp_48_ram[1150] = 71;
    exp_48_ram[1151] = 130;
    exp_48_ram[1152] = 39;
    exp_48_ram[1153] = 135;
    exp_48_ram[1154] = 44;
    exp_48_ram[1155] = 39;
    exp_48_ram[1156] = 7;
    exp_48_ram[1157] = 7;
    exp_48_ram[1158] = 128;
    exp_48_ram[1159] = 0;
    exp_48_ram[1160] = 39;
    exp_48_ram[1161] = 247;
    exp_48_ram[1162] = 130;
    exp_48_ram[1163] = 39;
    exp_48_ram[1164] = 135;
    exp_48_ram[1165] = 44;
    exp_48_ram[1166] = 39;
    exp_48_ram[1167] = 7;
    exp_48_ram[1168] = 7;
    exp_48_ram[1169] = 128;
    exp_48_ram[1170] = 0;
    exp_48_ram[1171] = 39;
    exp_48_ram[1172] = 247;
    exp_48_ram[1173] = 128;
    exp_48_ram[1174] = 39;
    exp_48_ram[1175] = 135;
    exp_48_ram[1176] = 44;
    exp_48_ram[1177] = 39;
    exp_48_ram[1178] = 7;
    exp_48_ram[1179] = 7;
    exp_48_ram[1180] = 128;
    exp_48_ram[1181] = 40;
    exp_48_ram[1182] = 40;
    exp_48_ram[1183] = 39;
    exp_48_ram[1184] = 39;
    exp_48_ram[1185] = 38;
    exp_48_ram[1186] = 38;
    exp_48_ram[1187] = 37;
    exp_48_ram[1188] = 37;
    exp_48_ram[1189] = 240;
    exp_48_ram[1190] = 7;
    exp_48_ram[1191] = 133;
    exp_48_ram[1192] = 32;
    exp_48_ram[1193] = 36;
    exp_48_ram[1194] = 1;
    exp_48_ram[1195] = 128;
    exp_48_ram[1196] = 1;
    exp_48_ram[1197] = 38;
    exp_48_ram[1198] = 36;
    exp_48_ram[1199] = 4;
    exp_48_ram[1200] = 46;
    exp_48_ram[1201] = 44;
    exp_48_ram[1202] = 42;
    exp_48_ram[1203] = 40;
    exp_48_ram[1204] = 38;
    exp_48_ram[1205] = 34;
    exp_48_ram[1206] = 32;
    exp_48_ram[1207] = 5;
    exp_48_ram[1208] = 38;
    exp_48_ram[1209] = 39;
    exp_48_ram[1210] = 152;
    exp_48_ram[1211] = 39;
    exp_48_ram[1212] = 247;
    exp_48_ram[1213] = 34;
    exp_48_ram[1214] = 39;
    exp_48_ram[1215] = 247;
    exp_48_ram[1216] = 134;
    exp_48_ram[1217] = 39;
    exp_48_ram[1218] = 140;
    exp_48_ram[1219] = 39;
    exp_48_ram[1220] = 39;
    exp_48_ram[1221] = 119;
    exp_48_ram[1222] = 5;
    exp_48_ram[1223] = 71;
    exp_48_ram[1224] = 7;
    exp_48_ram[1225] = 234;
    exp_48_ram[1226] = 71;
    exp_48_ram[1227] = 135;
    exp_48_ram[1228] = 247;
    exp_48_ram[1229] = 0;
    exp_48_ram[1230] = 39;
    exp_48_ram[1231] = 247;
    exp_48_ram[1232] = 134;
    exp_48_ram[1233] = 7;
    exp_48_ram[1234] = 0;
    exp_48_ram[1235] = 7;
    exp_48_ram[1236] = 71;
    exp_48_ram[1237] = 135;
    exp_48_ram[1238] = 247;
    exp_48_ram[1239] = 135;
    exp_48_ram[1240] = 247;
    exp_48_ram[1241] = 39;
    exp_48_ram[1242] = 6;
    exp_48_ram[1243] = 38;
    exp_48_ram[1244] = 6;
    exp_48_ram[1245] = 135;
    exp_48_ram[1246] = 12;
    exp_48_ram[1247] = 39;
    exp_48_ram[1248] = 39;
    exp_48_ram[1249] = 87;
    exp_48_ram[1250] = 38;
    exp_48_ram[1251] = 39;
    exp_48_ram[1252] = 136;
    exp_48_ram[1253] = 39;
    exp_48_ram[1254] = 7;
    exp_48_ram[1255] = 248;
    exp_48_ram[1256] = 70;
    exp_48_ram[1257] = 7;
    exp_48_ram[1258] = 39;
    exp_48_ram[1259] = 36;
    exp_48_ram[1260] = 39;
    exp_48_ram[1261] = 34;
    exp_48_ram[1262] = 39;
    exp_48_ram[1263] = 32;
    exp_48_ram[1264] = 40;
    exp_48_ram[1265] = 136;
    exp_48_ram[1266] = 39;
    exp_48_ram[1267] = 38;
    exp_48_ram[1268] = 38;
    exp_48_ram[1269] = 37;
    exp_48_ram[1270] = 37;
    exp_48_ram[1271] = 240;
    exp_48_ram[1272] = 7;
    exp_48_ram[1273] = 133;
    exp_48_ram[1274] = 32;
    exp_48_ram[1275] = 36;
    exp_48_ram[1276] = 1;
    exp_48_ram[1277] = 128;
    exp_48_ram[1278] = 1;
    exp_48_ram[1279] = 46;
    exp_48_ram[1280] = 44;
    exp_48_ram[1281] = 4;
    exp_48_ram[1282] = 38;
    exp_48_ram[1283] = 36;
    exp_48_ram[1284] = 34;
    exp_48_ram[1285] = 32;
    exp_48_ram[1286] = 46;
    exp_48_ram[1287] = 46;
    exp_48_ram[1288] = 39;
    exp_48_ram[1289] = 158;
    exp_48_ram[1290] = 23;
    exp_48_ram[1291] = 135;
    exp_48_ram[1292] = 38;
    exp_48_ram[1293] = 0;
    exp_48_ram[1294] = 39;
    exp_48_ram[1295] = 199;
    exp_48_ram[1296] = 7;
    exp_48_ram[1297] = 14;
    exp_48_ram[1298] = 39;
    exp_48_ram[1299] = 197;
    exp_48_ram[1300] = 39;
    exp_48_ram[1301] = 135;
    exp_48_ram[1302] = 46;
    exp_48_ram[1303] = 39;
    exp_48_ram[1304] = 38;
    exp_48_ram[1305] = 134;
    exp_48_ram[1306] = 37;
    exp_48_ram[1307] = 0;
    exp_48_ram[1308] = 39;
    exp_48_ram[1309] = 135;
    exp_48_ram[1310] = 32;
    exp_48_ram[1311] = 0;
    exp_48_ram[1312] = 39;
    exp_48_ram[1313] = 135;
    exp_48_ram[1314] = 32;
    exp_48_ram[1315] = 38;
    exp_48_ram[1316] = 39;
    exp_48_ram[1317] = 199;
    exp_48_ram[1318] = 135;
    exp_48_ram[1319] = 7;
    exp_48_ram[1320] = 104;
    exp_48_ram[1321] = 151;
    exp_48_ram[1322] = 71;
    exp_48_ram[1323] = 135;
    exp_48_ram[1324] = 7;
    exp_48_ram[1325] = 167;
    exp_48_ram[1326] = 128;
    exp_48_ram[1327] = 39;
    exp_48_ram[1328] = 231;
    exp_48_ram[1329] = 38;
    exp_48_ram[1330] = 39;
    exp_48_ram[1331] = 135;
    exp_48_ram[1332] = 32;
    exp_48_ram[1333] = 7;
    exp_48_ram[1334] = 32;
    exp_48_ram[1335] = 0;
    exp_48_ram[1336] = 39;
    exp_48_ram[1337] = 231;
    exp_48_ram[1338] = 38;
    exp_48_ram[1339] = 39;
    exp_48_ram[1340] = 135;
    exp_48_ram[1341] = 32;
    exp_48_ram[1342] = 7;
    exp_48_ram[1343] = 32;
    exp_48_ram[1344] = 0;
    exp_48_ram[1345] = 39;
    exp_48_ram[1346] = 231;
    exp_48_ram[1347] = 38;
    exp_48_ram[1348] = 39;
    exp_48_ram[1349] = 135;
    exp_48_ram[1350] = 32;
    exp_48_ram[1351] = 7;
    exp_48_ram[1352] = 32;
    exp_48_ram[1353] = 0;
    exp_48_ram[1354] = 39;
    exp_48_ram[1355] = 231;
    exp_48_ram[1356] = 38;
    exp_48_ram[1357] = 39;
    exp_48_ram[1358] = 135;
    exp_48_ram[1359] = 32;
    exp_48_ram[1360] = 7;
    exp_48_ram[1361] = 32;
    exp_48_ram[1362] = 0;
    exp_48_ram[1363] = 39;
    exp_48_ram[1364] = 231;
    exp_48_ram[1365] = 38;
    exp_48_ram[1366] = 39;
    exp_48_ram[1367] = 135;
    exp_48_ram[1368] = 32;
    exp_48_ram[1369] = 7;
    exp_48_ram[1370] = 32;
    exp_48_ram[1371] = 0;
    exp_48_ram[1372] = 32;
    exp_48_ram[1373] = 0;
    exp_48_ram[1374] = 39;
    exp_48_ram[1375] = 154;
    exp_48_ram[1376] = 36;
    exp_48_ram[1377] = 39;
    exp_48_ram[1378] = 199;
    exp_48_ram[1379] = 133;
    exp_48_ram[1380] = 240;
    exp_48_ram[1381] = 7;
    exp_48_ram[1382] = 140;
    exp_48_ram[1383] = 7;
    exp_48_ram[1384] = 133;
    exp_48_ram[1385] = 240;
    exp_48_ram[1386] = 36;
    exp_48_ram[1387] = 0;
    exp_48_ram[1388] = 39;
    exp_48_ram[1389] = 199;
    exp_48_ram[1390] = 7;
    exp_48_ram[1391] = 24;
    exp_48_ram[1392] = 39;
    exp_48_ram[1393] = 135;
    exp_48_ram[1394] = 46;
    exp_48_ram[1395] = 167;
    exp_48_ram[1396] = 36;
    exp_48_ram[1397] = 39;
    exp_48_ram[1398] = 208;
    exp_48_ram[1399] = 39;
    exp_48_ram[1400] = 231;
    exp_48_ram[1401] = 38;
    exp_48_ram[1402] = 39;
    exp_48_ram[1403] = 7;
    exp_48_ram[1404] = 36;
    exp_48_ram[1405] = 0;
    exp_48_ram[1406] = 39;
    exp_48_ram[1407] = 36;
    exp_48_ram[1408] = 39;
    exp_48_ram[1409] = 135;
    exp_48_ram[1410] = 32;
    exp_48_ram[1411] = 34;
    exp_48_ram[1412] = 39;
    exp_48_ram[1413] = 199;
    exp_48_ram[1414] = 7;
    exp_48_ram[1415] = 20;
    exp_48_ram[1416] = 39;
    exp_48_ram[1417] = 231;
    exp_48_ram[1418] = 38;
    exp_48_ram[1419] = 39;
    exp_48_ram[1420] = 135;
    exp_48_ram[1421] = 32;
    exp_48_ram[1422] = 39;
    exp_48_ram[1423] = 199;
    exp_48_ram[1424] = 133;
    exp_48_ram[1425] = 240;
    exp_48_ram[1426] = 7;
    exp_48_ram[1427] = 140;
    exp_48_ram[1428] = 7;
    exp_48_ram[1429] = 133;
    exp_48_ram[1430] = 240;
    exp_48_ram[1431] = 34;
    exp_48_ram[1432] = 0;
    exp_48_ram[1433] = 39;
    exp_48_ram[1434] = 199;
    exp_48_ram[1435] = 7;
    exp_48_ram[1436] = 26;
    exp_48_ram[1437] = 39;
    exp_48_ram[1438] = 135;
    exp_48_ram[1439] = 46;
    exp_48_ram[1440] = 167;
    exp_48_ram[1441] = 34;
    exp_48_ram[1442] = 39;
    exp_48_ram[1443] = 212;
    exp_48_ram[1444] = 7;
    exp_48_ram[1445] = 34;
    exp_48_ram[1446] = 39;
    exp_48_ram[1447] = 135;
    exp_48_ram[1448] = 32;
    exp_48_ram[1449] = 39;
    exp_48_ram[1450] = 199;
    exp_48_ram[1451] = 135;
    exp_48_ram[1452] = 7;
    exp_48_ram[1453] = 108;
    exp_48_ram[1454] = 151;
    exp_48_ram[1455] = 71;
    exp_48_ram[1456] = 135;
    exp_48_ram[1457] = 7;
    exp_48_ram[1458] = 167;
    exp_48_ram[1459] = 128;
    exp_48_ram[1460] = 39;
    exp_48_ram[1461] = 231;
    exp_48_ram[1462] = 38;
    exp_48_ram[1463] = 39;
    exp_48_ram[1464] = 135;
    exp_48_ram[1465] = 32;
    exp_48_ram[1466] = 39;
    exp_48_ram[1467] = 199;
    exp_48_ram[1468] = 7;
    exp_48_ram[1469] = 16;
    exp_48_ram[1470] = 39;
    exp_48_ram[1471] = 231;
    exp_48_ram[1472] = 38;
    exp_48_ram[1473] = 39;
    exp_48_ram[1474] = 135;
    exp_48_ram[1475] = 32;
    exp_48_ram[1476] = 0;
    exp_48_ram[1477] = 39;
    exp_48_ram[1478] = 231;
    exp_48_ram[1479] = 38;
    exp_48_ram[1480] = 39;
    exp_48_ram[1481] = 135;
    exp_48_ram[1482] = 32;
    exp_48_ram[1483] = 39;
    exp_48_ram[1484] = 199;
    exp_48_ram[1485] = 7;
    exp_48_ram[1486] = 18;
    exp_48_ram[1487] = 39;
    exp_48_ram[1488] = 231;
    exp_48_ram[1489] = 38;
    exp_48_ram[1490] = 39;
    exp_48_ram[1491] = 135;
    exp_48_ram[1492] = 32;
    exp_48_ram[1493] = 0;
    exp_48_ram[1494] = 39;
    exp_48_ram[1495] = 231;
    exp_48_ram[1496] = 38;
    exp_48_ram[1497] = 39;
    exp_48_ram[1498] = 135;
    exp_48_ram[1499] = 32;
    exp_48_ram[1500] = 0;
    exp_48_ram[1501] = 39;
    exp_48_ram[1502] = 231;
    exp_48_ram[1503] = 38;
    exp_48_ram[1504] = 39;
    exp_48_ram[1505] = 135;
    exp_48_ram[1506] = 32;
    exp_48_ram[1507] = 0;
    exp_48_ram[1508] = 39;
    exp_48_ram[1509] = 231;
    exp_48_ram[1510] = 38;
    exp_48_ram[1511] = 39;
    exp_48_ram[1512] = 135;
    exp_48_ram[1513] = 32;
    exp_48_ram[1514] = 0;
    exp_48_ram[1515] = 0;
    exp_48_ram[1516] = 0;
    exp_48_ram[1517] = 0;
    exp_48_ram[1518] = 0;
    exp_48_ram[1519] = 0;
    exp_48_ram[1520] = 39;
    exp_48_ram[1521] = 199;
    exp_48_ram[1522] = 135;
    exp_48_ram[1523] = 7;
    exp_48_ram[1524] = 108;
    exp_48_ram[1525] = 151;
    exp_48_ram[1526] = 71;
    exp_48_ram[1527] = 135;
    exp_48_ram[1528] = 7;
    exp_48_ram[1529] = 167;
    exp_48_ram[1530] = 128;
    exp_48_ram[1531] = 39;
    exp_48_ram[1532] = 199;
    exp_48_ram[1533] = 7;
    exp_48_ram[1534] = 10;
    exp_48_ram[1535] = 39;
    exp_48_ram[1536] = 199;
    exp_48_ram[1537] = 7;
    exp_48_ram[1538] = 24;
    exp_48_ram[1539] = 7;
    exp_48_ram[1540] = 44;
    exp_48_ram[1541] = 0;
    exp_48_ram[1542] = 39;
    exp_48_ram[1543] = 199;
    exp_48_ram[1544] = 7;
    exp_48_ram[1545] = 24;
    exp_48_ram[1546] = 7;
    exp_48_ram[1547] = 44;
    exp_48_ram[1548] = 0;
    exp_48_ram[1549] = 39;
    exp_48_ram[1550] = 199;
    exp_48_ram[1551] = 7;
    exp_48_ram[1552] = 24;
    exp_48_ram[1553] = 7;
    exp_48_ram[1554] = 44;
    exp_48_ram[1555] = 0;
    exp_48_ram[1556] = 7;
    exp_48_ram[1557] = 44;
    exp_48_ram[1558] = 39;
    exp_48_ram[1559] = 247;
    exp_48_ram[1560] = 38;
    exp_48_ram[1561] = 39;
    exp_48_ram[1562] = 199;
    exp_48_ram[1563] = 7;
    exp_48_ram[1564] = 24;
    exp_48_ram[1565] = 39;
    exp_48_ram[1566] = 231;
    exp_48_ram[1567] = 38;
    exp_48_ram[1568] = 39;
    exp_48_ram[1569] = 199;
    exp_48_ram[1570] = 7;
    exp_48_ram[1571] = 0;
    exp_48_ram[1572] = 39;
    exp_48_ram[1573] = 199;
    exp_48_ram[1574] = 7;
    exp_48_ram[1575] = 8;
    exp_48_ram[1576] = 39;
    exp_48_ram[1577] = 247;
    exp_48_ram[1578] = 38;
    exp_48_ram[1579] = 39;
    exp_48_ram[1580] = 247;
    exp_48_ram[1581] = 136;
    exp_48_ram[1582] = 39;
    exp_48_ram[1583] = 247;
    exp_48_ram[1584] = 38;
    exp_48_ram[1585] = 39;
    exp_48_ram[1586] = 199;
    exp_48_ram[1587] = 7;
    exp_48_ram[1588] = 10;
    exp_48_ram[1589] = 39;
    exp_48_ram[1590] = 199;
    exp_48_ram[1591] = 7;
    exp_48_ram[1592] = 24;
    exp_48_ram[1593] = 39;
    exp_48_ram[1594] = 247;
    exp_48_ram[1595] = 158;
    exp_48_ram[1596] = 39;
    exp_48_ram[1597] = 247;
    exp_48_ram[1598] = 140;
    exp_48_ram[1599] = 39;
    exp_48_ram[1600] = 135;
    exp_48_ram[1601] = 46;
    exp_48_ram[1602] = 167;
    exp_48_ram[1603] = 44;
    exp_48_ram[1604] = 39;
    exp_48_ram[1605] = 215;
    exp_48_ram[1606] = 39;
    exp_48_ram[1607] = 71;
    exp_48_ram[1608] = 135;
    exp_48_ram[1609] = 134;
    exp_48_ram[1610] = 39;
    exp_48_ram[1611] = 215;
    exp_48_ram[1612] = 247;
    exp_48_ram[1613] = 39;
    exp_48_ram[1614] = 34;
    exp_48_ram[1615] = 39;
    exp_48_ram[1616] = 32;
    exp_48_ram[1617] = 40;
    exp_48_ram[1618] = 40;
    exp_48_ram[1619] = 7;
    exp_48_ram[1620] = 135;
    exp_48_ram[1621] = 38;
    exp_48_ram[1622] = 38;
    exp_48_ram[1623] = 37;
    exp_48_ram[1624] = 37;
    exp_48_ram[1625] = 240;
    exp_48_ram[1626] = 46;
    exp_48_ram[1627] = 0;
    exp_48_ram[1628] = 39;
    exp_48_ram[1629] = 247;
    exp_48_ram[1630] = 142;
    exp_48_ram[1631] = 39;
    exp_48_ram[1632] = 135;
    exp_48_ram[1633] = 46;
    exp_48_ram[1634] = 167;
    exp_48_ram[1635] = 247;
    exp_48_ram[1636] = 0;
    exp_48_ram[1637] = 39;
    exp_48_ram[1638] = 247;
    exp_48_ram[1639] = 128;
    exp_48_ram[1640] = 39;
    exp_48_ram[1641] = 135;
    exp_48_ram[1642] = 46;
    exp_48_ram[1643] = 167;
    exp_48_ram[1644] = 151;
    exp_48_ram[1645] = 215;
    exp_48_ram[1646] = 0;
    exp_48_ram[1647] = 39;
    exp_48_ram[1648] = 135;
    exp_48_ram[1649] = 46;
    exp_48_ram[1650] = 167;
    exp_48_ram[1651] = 46;
    exp_48_ram[1652] = 39;
    exp_48_ram[1653] = 215;
    exp_48_ram[1654] = 39;
    exp_48_ram[1655] = 71;
    exp_48_ram[1656] = 135;
    exp_48_ram[1657] = 134;
    exp_48_ram[1658] = 39;
    exp_48_ram[1659] = 215;
    exp_48_ram[1660] = 247;
    exp_48_ram[1661] = 39;
    exp_48_ram[1662] = 34;
    exp_48_ram[1663] = 39;
    exp_48_ram[1664] = 32;
    exp_48_ram[1665] = 40;
    exp_48_ram[1666] = 40;
    exp_48_ram[1667] = 7;
    exp_48_ram[1668] = 135;
    exp_48_ram[1669] = 38;
    exp_48_ram[1670] = 38;
    exp_48_ram[1671] = 37;
    exp_48_ram[1672] = 37;
    exp_48_ram[1673] = 240;
    exp_48_ram[1674] = 46;
    exp_48_ram[1675] = 0;
    exp_48_ram[1676] = 39;
    exp_48_ram[1677] = 247;
    exp_48_ram[1678] = 152;
    exp_48_ram[1679] = 39;
    exp_48_ram[1680] = 247;
    exp_48_ram[1681] = 134;
    exp_48_ram[1682] = 39;
    exp_48_ram[1683] = 135;
    exp_48_ram[1684] = 46;
    exp_48_ram[1685] = 167;
    exp_48_ram[1686] = 39;
    exp_48_ram[1687] = 34;
    exp_48_ram[1688] = 39;
    exp_48_ram[1689] = 32;
    exp_48_ram[1690] = 40;
    exp_48_ram[1691] = 40;
    exp_48_ram[1692] = 7;
    exp_48_ram[1693] = 38;
    exp_48_ram[1694] = 38;
    exp_48_ram[1695] = 37;
    exp_48_ram[1696] = 37;
    exp_48_ram[1697] = 240;
    exp_48_ram[1698] = 46;
    exp_48_ram[1699] = 0;
    exp_48_ram[1700] = 39;
    exp_48_ram[1701] = 247;
    exp_48_ram[1702] = 142;
    exp_48_ram[1703] = 39;
    exp_48_ram[1704] = 135;
    exp_48_ram[1705] = 46;
    exp_48_ram[1706] = 167;
    exp_48_ram[1707] = 247;
    exp_48_ram[1708] = 0;
    exp_48_ram[1709] = 39;
    exp_48_ram[1710] = 247;
    exp_48_ram[1711] = 128;
    exp_48_ram[1712] = 39;
    exp_48_ram[1713] = 135;
    exp_48_ram[1714] = 46;
    exp_48_ram[1715] = 167;
    exp_48_ram[1716] = 151;
    exp_48_ram[1717] = 215;
    exp_48_ram[1718] = 0;
    exp_48_ram[1719] = 39;
    exp_48_ram[1720] = 135;
    exp_48_ram[1721] = 46;
    exp_48_ram[1722] = 167;
    exp_48_ram[1723] = 32;
    exp_48_ram[1724] = 39;
    exp_48_ram[1725] = 34;
    exp_48_ram[1726] = 39;
    exp_48_ram[1727] = 32;
    exp_48_ram[1728] = 40;
    exp_48_ram[1729] = 40;
    exp_48_ram[1730] = 7;
    exp_48_ram[1731] = 39;
    exp_48_ram[1732] = 38;
    exp_48_ram[1733] = 38;
    exp_48_ram[1734] = 37;
    exp_48_ram[1735] = 37;
    exp_48_ram[1736] = 240;
    exp_48_ram[1737] = 46;
    exp_48_ram[1738] = 39;
    exp_48_ram[1739] = 135;
    exp_48_ram[1740] = 32;
    exp_48_ram[1741] = 0;
    exp_48_ram[1742] = 7;
    exp_48_ram[1743] = 42;
    exp_48_ram[1744] = 39;
    exp_48_ram[1745] = 247;
    exp_48_ram[1746] = 144;
    exp_48_ram[1747] = 0;
    exp_48_ram[1748] = 39;
    exp_48_ram[1749] = 135;
    exp_48_ram[1750] = 46;
    exp_48_ram[1751] = 39;
    exp_48_ram[1752] = 38;
    exp_48_ram[1753] = 134;
    exp_48_ram[1754] = 37;
    exp_48_ram[1755] = 5;
    exp_48_ram[1756] = 0;
    exp_48_ram[1757] = 39;
    exp_48_ram[1758] = 135;
    exp_48_ram[1759] = 42;
    exp_48_ram[1760] = 39;
    exp_48_ram[1761] = 230;
    exp_48_ram[1762] = 39;
    exp_48_ram[1763] = 135;
    exp_48_ram[1764] = 46;
    exp_48_ram[1765] = 167;
    exp_48_ram[1766] = 245;
    exp_48_ram[1767] = 39;
    exp_48_ram[1768] = 135;
    exp_48_ram[1769] = 46;
    exp_48_ram[1770] = 39;
    exp_48_ram[1771] = 38;
    exp_48_ram[1772] = 134;
    exp_48_ram[1773] = 37;
    exp_48_ram[1774] = 0;
    exp_48_ram[1775] = 39;
    exp_48_ram[1776] = 247;
    exp_48_ram[1777] = 128;
    exp_48_ram[1778] = 0;
    exp_48_ram[1779] = 39;
    exp_48_ram[1780] = 135;
    exp_48_ram[1781] = 46;
    exp_48_ram[1782] = 39;
    exp_48_ram[1783] = 38;
    exp_48_ram[1784] = 134;
    exp_48_ram[1785] = 37;
    exp_48_ram[1786] = 5;
    exp_48_ram[1787] = 0;
    exp_48_ram[1788] = 39;
    exp_48_ram[1789] = 135;
    exp_48_ram[1790] = 42;
    exp_48_ram[1791] = 39;
    exp_48_ram[1792] = 230;
    exp_48_ram[1793] = 39;
    exp_48_ram[1794] = 135;
    exp_48_ram[1795] = 32;
    exp_48_ram[1796] = 0;
    exp_48_ram[1797] = 39;
    exp_48_ram[1798] = 135;
    exp_48_ram[1799] = 46;
    exp_48_ram[1800] = 167;
    exp_48_ram[1801] = 40;
    exp_48_ram[1802] = 39;
    exp_48_ram[1803] = 134;
    exp_48_ram[1804] = 39;
    exp_48_ram[1805] = 0;
    exp_48_ram[1806] = 7;
    exp_48_ram[1807] = 133;
    exp_48_ram[1808] = 37;
    exp_48_ram[1809] = 240;
    exp_48_ram[1810] = 38;
    exp_48_ram[1811] = 39;
    exp_48_ram[1812] = 247;
    exp_48_ram[1813] = 140;
    exp_48_ram[1814] = 39;
    exp_48_ram[1815] = 39;
    exp_48_ram[1816] = 116;
    exp_48_ram[1817] = 7;
    exp_48_ram[1818] = 38;
    exp_48_ram[1819] = 39;
    exp_48_ram[1820] = 247;
    exp_48_ram[1821] = 154;
    exp_48_ram[1822] = 0;
    exp_48_ram[1823] = 39;
    exp_48_ram[1824] = 135;
    exp_48_ram[1825] = 46;
    exp_48_ram[1826] = 39;
    exp_48_ram[1827] = 38;
    exp_48_ram[1828] = 134;
    exp_48_ram[1829] = 37;
    exp_48_ram[1830] = 5;
    exp_48_ram[1831] = 0;
    exp_48_ram[1832] = 39;
    exp_48_ram[1833] = 135;
    exp_48_ram[1834] = 38;
    exp_48_ram[1835] = 39;
    exp_48_ram[1836] = 230;
    exp_48_ram[1837] = 0;
    exp_48_ram[1838] = 39;
    exp_48_ram[1839] = 135;
    exp_48_ram[1840] = 40;
    exp_48_ram[1841] = 197;
    exp_48_ram[1842] = 39;
    exp_48_ram[1843] = 135;
    exp_48_ram[1844] = 46;
    exp_48_ram[1845] = 39;
    exp_48_ram[1846] = 38;
    exp_48_ram[1847] = 134;
    exp_48_ram[1848] = 37;
    exp_48_ram[1849] = 0;
    exp_48_ram[1850] = 39;
    exp_48_ram[1851] = 199;
    exp_48_ram[1852] = 128;
    exp_48_ram[1853] = 39;
    exp_48_ram[1854] = 247;
    exp_48_ram[1855] = 142;
    exp_48_ram[1856] = 39;
    exp_48_ram[1857] = 135;
    exp_48_ram[1858] = 34;
    exp_48_ram[1859] = 150;
    exp_48_ram[1860] = 39;
    exp_48_ram[1861] = 247;
    exp_48_ram[1862] = 128;
    exp_48_ram[1863] = 0;
    exp_48_ram[1864] = 39;
    exp_48_ram[1865] = 135;
    exp_48_ram[1866] = 46;
    exp_48_ram[1867] = 39;
    exp_48_ram[1868] = 38;
    exp_48_ram[1869] = 134;
    exp_48_ram[1870] = 37;
    exp_48_ram[1871] = 5;
    exp_48_ram[1872] = 0;
    exp_48_ram[1873] = 39;
    exp_48_ram[1874] = 135;
    exp_48_ram[1875] = 38;
    exp_48_ram[1876] = 39;
    exp_48_ram[1877] = 230;
    exp_48_ram[1878] = 39;
    exp_48_ram[1879] = 135;
    exp_48_ram[1880] = 32;
    exp_48_ram[1881] = 0;
    exp_48_ram[1882] = 7;
    exp_48_ram[1883] = 36;
    exp_48_ram[1884] = 39;
    exp_48_ram[1885] = 231;
    exp_48_ram[1886] = 38;
    exp_48_ram[1887] = 39;
    exp_48_ram[1888] = 135;
    exp_48_ram[1889] = 46;
    exp_48_ram[1890] = 167;
    exp_48_ram[1891] = 135;
    exp_48_ram[1892] = 39;
    exp_48_ram[1893] = 34;
    exp_48_ram[1894] = 39;
    exp_48_ram[1895] = 32;
    exp_48_ram[1896] = 40;
    exp_48_ram[1897] = 8;
    exp_48_ram[1898] = 7;
    exp_48_ram[1899] = 38;
    exp_48_ram[1900] = 38;
    exp_48_ram[1901] = 37;
    exp_48_ram[1902] = 37;
    exp_48_ram[1903] = 240;
    exp_48_ram[1904] = 46;
    exp_48_ram[1905] = 39;
    exp_48_ram[1906] = 135;
    exp_48_ram[1907] = 32;
    exp_48_ram[1908] = 0;
    exp_48_ram[1909] = 39;
    exp_48_ram[1910] = 135;
    exp_48_ram[1911] = 46;
    exp_48_ram[1912] = 39;
    exp_48_ram[1913] = 38;
    exp_48_ram[1914] = 134;
    exp_48_ram[1915] = 37;
    exp_48_ram[1916] = 5;
    exp_48_ram[1917] = 0;
    exp_48_ram[1918] = 39;
    exp_48_ram[1919] = 135;
    exp_48_ram[1920] = 32;
    exp_48_ram[1921] = 0;
    exp_48_ram[1922] = 39;
    exp_48_ram[1923] = 197;
    exp_48_ram[1924] = 39;
    exp_48_ram[1925] = 135;
    exp_48_ram[1926] = 46;
    exp_48_ram[1927] = 39;
    exp_48_ram[1928] = 38;
    exp_48_ram[1929] = 134;
    exp_48_ram[1930] = 37;
    exp_48_ram[1931] = 0;
    exp_48_ram[1932] = 39;
    exp_48_ram[1933] = 135;
    exp_48_ram[1934] = 32;
    exp_48_ram[1935] = 0;
    exp_48_ram[1936] = 39;
    exp_48_ram[1937] = 199;
    exp_48_ram[1938] = 152;
    exp_48_ram[1939] = 39;
    exp_48_ram[1940] = 39;
    exp_48_ram[1941] = 104;
    exp_48_ram[1942] = 39;
    exp_48_ram[1943] = 135;
    exp_48_ram[1944] = 0;
    exp_48_ram[1945] = 39;
    exp_48_ram[1946] = 39;
    exp_48_ram[1947] = 38;
    exp_48_ram[1948] = 134;
    exp_48_ram[1949] = 37;
    exp_48_ram[1950] = 5;
    exp_48_ram[1951] = 0;
    exp_48_ram[1952] = 39;
    exp_48_ram[1953] = 133;
    exp_48_ram[1954] = 32;
    exp_48_ram[1955] = 36;
    exp_48_ram[1956] = 1;
    exp_48_ram[1957] = 128;
    exp_48_ram[1958] = 1;
    exp_48_ram[1959] = 38;
    exp_48_ram[1960] = 36;
    exp_48_ram[1961] = 4;
    exp_48_ram[1962] = 46;
    exp_48_ram[1963] = 34;
    exp_48_ram[1964] = 36;
    exp_48_ram[1965] = 38;
    exp_48_ram[1966] = 40;
    exp_48_ram[1967] = 42;
    exp_48_ram[1968] = 44;
    exp_48_ram[1969] = 46;
    exp_48_ram[1970] = 7;
    exp_48_ram[1971] = 44;
    exp_48_ram[1972] = 39;
    exp_48_ram[1973] = 135;
    exp_48_ram[1974] = 36;
    exp_48_ram[1975] = 39;
    exp_48_ram[1976] = 7;
    exp_48_ram[1977] = 38;
    exp_48_ram[1978] = 6;
    exp_48_ram[1979] = 133;
    exp_48_ram[1980] = 23;
    exp_48_ram[1981] = 133;
    exp_48_ram[1982] = 240;
    exp_48_ram[1983] = 38;
    exp_48_ram[1984] = 39;
    exp_48_ram[1985] = 133;
    exp_48_ram[1986] = 32;
    exp_48_ram[1987] = 36;
    exp_48_ram[1988] = 1;
    exp_48_ram[1989] = 128;
    exp_48_ram[1990] = 1;
    exp_48_ram[1991] = 46;
    exp_48_ram[1992] = 44;
    exp_48_ram[1993] = 4;
    exp_48_ram[1994] = 7;
    exp_48_ram[1995] = 7;
    exp_48_ram[1996] = 71;
    exp_48_ram[1997] = 71;
    exp_48_ram[1998] = 167;
    exp_48_ram[1999] = 133;
    exp_48_ram[2000] = 5;
    exp_48_ram[2001] = 224;
    exp_48_ram[2002] = 0;
    exp_48_ram[2003] = 32;
    exp_48_ram[2004] = 36;
    exp_48_ram[2005] = 1;
    exp_48_ram[2006] = 128;
    exp_48_ram[2007] = 1;
    exp_48_ram[2008] = 46;
    exp_48_ram[2009] = 44;
    exp_48_ram[2010] = 42;
    exp_48_ram[2011] = 4;
    exp_48_ram[2012] = 4;
    exp_48_ram[2013] = 167;
    exp_48_ram[2014] = 36;
    exp_48_ram[2015] = 7;
    exp_48_ram[2016] = 34;
    exp_48_ram[2017] = 7;
    exp_48_ram[2018] = 32;
    exp_48_ram[2019] = 7;
    exp_48_ram[2020] = 46;
    exp_48_ram[2021] = 44;
    exp_48_ram[2022] = 42;
    exp_48_ram[2023] = 42;
    exp_48_ram[2024] = 35;
    exp_48_ram[2025] = 40;
    exp_48_ram[2026] = 40;
    exp_48_ram[2027] = 37;
    exp_48_ram[2028] = 37;
    exp_48_ram[2029] = 38;
    exp_48_ram[2030] = 38;
    exp_48_ram[2031] = 39;
    exp_48_ram[2032] = 39;
    exp_48_ram[2033] = 32;
    exp_48_ram[2034] = 34;
    exp_48_ram[2035] = 36;
    exp_48_ram[2036] = 38;
    exp_48_ram[2037] = 40;
    exp_48_ram[2038] = 42;
    exp_48_ram[2039] = 44;
    exp_48_ram[2040] = 46;
    exp_48_ram[2041] = 32;
    exp_48_ram[2042] = 7;
    exp_48_ram[2043] = 133;
    exp_48_ram[2044] = 0;
    exp_48_ram[2045] = 36;
    exp_48_ram[2046] = 38;
    exp_48_ram[2047] = 7;
    exp_48_ram[2048] = 37;
    exp_48_ram[2049] = 38;
    exp_48_ram[2050] = 133;
    exp_48_ram[2051] = 16;
    exp_48_ram[2052] = 39;
    exp_48_ram[2053] = 39;
    exp_48_ram[2054] = 7;
    exp_48_ram[2055] = 32;
    exp_48_ram[2056] = 35;
    exp_48_ram[2057] = 40;
    exp_48_ram[2058] = 40;
    exp_48_ram[2059] = 37;
    exp_48_ram[2060] = 37;
    exp_48_ram[2061] = 38;
    exp_48_ram[2062] = 38;
    exp_48_ram[2063] = 39;
    exp_48_ram[2064] = 39;
    exp_48_ram[2065] = 32;
    exp_48_ram[2066] = 34;
    exp_48_ram[2067] = 36;
    exp_48_ram[2068] = 38;
    exp_48_ram[2069] = 40;
    exp_48_ram[2070] = 42;
    exp_48_ram[2071] = 44;
    exp_48_ram[2072] = 46;
    exp_48_ram[2073] = 32;
    exp_48_ram[2074] = 7;
    exp_48_ram[2075] = 133;
    exp_48_ram[2076] = 0;
    exp_48_ram[2077] = 36;
    exp_48_ram[2078] = 38;
    exp_48_ram[2079] = 167;
    exp_48_ram[2080] = 34;
    exp_48_ram[2081] = 7;
    exp_48_ram[2082] = 32;
    exp_48_ram[2083] = 7;
    exp_48_ram[2084] = 46;
    exp_48_ram[2085] = 7;
    exp_48_ram[2086] = 44;
    exp_48_ram[2087] = 42;
    exp_48_ram[2088] = 40;
    exp_48_ram[2089] = 42;
    exp_48_ram[2090] = 35;
    exp_48_ram[2091] = 40;
    exp_48_ram[2092] = 40;
    exp_48_ram[2093] = 37;
    exp_48_ram[2094] = 37;
    exp_48_ram[2095] = 38;
    exp_48_ram[2096] = 38;
    exp_48_ram[2097] = 39;
    exp_48_ram[2098] = 39;
    exp_48_ram[2099] = 32;
    exp_48_ram[2100] = 34;
    exp_48_ram[2101] = 36;
    exp_48_ram[2102] = 38;
    exp_48_ram[2103] = 40;
    exp_48_ram[2104] = 42;
    exp_48_ram[2105] = 44;
    exp_48_ram[2106] = 46;
    exp_48_ram[2107] = 32;
    exp_48_ram[2108] = 7;
    exp_48_ram[2109] = 133;
    exp_48_ram[2110] = 0;
    exp_48_ram[2111] = 32;
    exp_48_ram[2112] = 34;
    exp_48_ram[2113] = 7;
    exp_48_ram[2114] = 37;
    exp_48_ram[2115] = 38;
    exp_48_ram[2116] = 133;
    exp_48_ram[2117] = 0;
    exp_48_ram[2118] = 39;
    exp_48_ram[2119] = 39;
    exp_48_ram[2120] = 7;
    exp_48_ram[2121] = 46;
    exp_48_ram[2122] = 35;
    exp_48_ram[2123] = 40;
    exp_48_ram[2124] = 40;
    exp_48_ram[2125] = 37;
    exp_48_ram[2126] = 37;
    exp_48_ram[2127] = 38;
    exp_48_ram[2128] = 38;
    exp_48_ram[2129] = 39;
    exp_48_ram[2130] = 39;
    exp_48_ram[2131] = 32;
    exp_48_ram[2132] = 34;
    exp_48_ram[2133] = 36;
    exp_48_ram[2134] = 38;
    exp_48_ram[2135] = 40;
    exp_48_ram[2136] = 42;
    exp_48_ram[2137] = 44;
    exp_48_ram[2138] = 46;
    exp_48_ram[2139] = 32;
    exp_48_ram[2140] = 7;
    exp_48_ram[2141] = 133;
    exp_48_ram[2142] = 0;
    exp_48_ram[2143] = 32;
    exp_48_ram[2144] = 34;
    exp_48_ram[2145] = 163;
    exp_48_ram[2146] = 168;
    exp_48_ram[2147] = 168;
    exp_48_ram[2148] = 165;
    exp_48_ram[2149] = 165;
    exp_48_ram[2150] = 166;
    exp_48_ram[2151] = 166;
    exp_48_ram[2152] = 167;
    exp_48_ram[2153] = 167;
    exp_48_ram[2154] = 32;
    exp_48_ram[2155] = 34;
    exp_48_ram[2156] = 36;
    exp_48_ram[2157] = 38;
    exp_48_ram[2158] = 40;
    exp_48_ram[2159] = 42;
    exp_48_ram[2160] = 44;
    exp_48_ram[2161] = 46;
    exp_48_ram[2162] = 32;
    exp_48_ram[2163] = 7;
    exp_48_ram[2164] = 133;
    exp_48_ram[2165] = 0;
    exp_48_ram[2166] = 44;
    exp_48_ram[2167] = 46;
    exp_48_ram[2168] = 39;
    exp_48_ram[2169] = 39;
    exp_48_ram[2170] = 228;
    exp_48_ram[2171] = 39;
    exp_48_ram[2172] = 39;
    exp_48_ram[2173] = 24;
    exp_48_ram[2174] = 39;
    exp_48_ram[2175] = 39;
    exp_48_ram[2176] = 232;
    exp_48_ram[2177] = 39;
    exp_48_ram[2178] = 39;
    exp_48_ram[2179] = 238;
    exp_48_ram[2180] = 39;
    exp_48_ram[2181] = 39;
    exp_48_ram[2182] = 28;
    exp_48_ram[2183] = 39;
    exp_48_ram[2184] = 39;
    exp_48_ram[2185] = 246;
    exp_48_ram[2186] = 7;
    exp_48_ram[2187] = 0;
    exp_48_ram[2188] = 7;
    exp_48_ram[2189] = 133;
    exp_48_ram[2190] = 32;
    exp_48_ram[2191] = 36;
    exp_48_ram[2192] = 36;
    exp_48_ram[2193] = 1;
    exp_48_ram[2194] = 128;
    exp_48_ram[2195] = 1;
    exp_48_ram[2196] = 46;
    exp_48_ram[2197] = 44;
    exp_48_ram[2198] = 4;
    exp_48_ram[2199] = 44;
    exp_48_ram[2200] = 46;
    exp_48_ram[2201] = 7;
    exp_48_ram[2202] = 37;
    exp_48_ram[2203] = 38;
    exp_48_ram[2204] = 133;
    exp_48_ram[2205] = 0;
    exp_48_ram[2206] = 35;
    exp_48_ram[2207] = 40;
    exp_48_ram[2208] = 40;
    exp_48_ram[2209] = 37;
    exp_48_ram[2210] = 37;
    exp_48_ram[2211] = 38;
    exp_48_ram[2212] = 38;
    exp_48_ram[2213] = 39;
    exp_48_ram[2214] = 39;
    exp_48_ram[2215] = 32;
    exp_48_ram[2216] = 34;
    exp_48_ram[2217] = 36;
    exp_48_ram[2218] = 38;
    exp_48_ram[2219] = 40;
    exp_48_ram[2220] = 42;
    exp_48_ram[2221] = 44;
    exp_48_ram[2222] = 46;
    exp_48_ram[2223] = 32;
    exp_48_ram[2224] = 7;
    exp_48_ram[2225] = 133;
    exp_48_ram[2226] = 240;
    exp_48_ram[2227] = 7;
    exp_48_ram[2228] = 133;
    exp_48_ram[2229] = 32;
    exp_48_ram[2230] = 36;
    exp_48_ram[2231] = 1;
    exp_48_ram[2232] = 128;
    exp_48_ram[2233] = 1;
    exp_48_ram[2234] = 46;
    exp_48_ram[2235] = 4;
    exp_48_ram[2236] = 6;
    exp_48_ram[2237] = 38;
    exp_48_ram[2238] = 6;
    exp_48_ram[2239] = 134;
    exp_48_ram[2240] = 36;
    exp_48_ram[2241] = 38;
    exp_48_ram[2242] = 166;
    exp_48_ram[2243] = 32;
    exp_48_ram[2244] = 34;
    exp_48_ram[2245] = 38;
    exp_48_ram[2246] = 150;
    exp_48_ram[2247] = 34;
    exp_48_ram[2248] = 32;
    exp_48_ram[2249] = 38;
    exp_48_ram[2250] = 166;
    exp_48_ram[2251] = 135;
    exp_48_ram[2252] = 7;
    exp_48_ram[2253] = 38;
    exp_48_ram[2254] = 230;
    exp_48_ram[2255] = 32;
    exp_48_ram[2256] = 38;
    exp_48_ram[2257] = 231;
    exp_48_ram[2258] = 34;
    exp_48_ram[2259] = 39;
    exp_48_ram[2260] = 39;
    exp_48_ram[2261] = 5;
    exp_48_ram[2262] = 133;
    exp_48_ram[2263] = 36;
    exp_48_ram[2264] = 1;
    exp_48_ram[2265] = 128;
    exp_48_ram[2266] = 1;
    exp_48_ram[2267] = 46;
    exp_48_ram[2268] = 44;
    exp_48_ram[2269] = 4;
    exp_48_ram[2270] = 36;
    exp_48_ram[2271] = 38;
    exp_48_ram[2272] = 32;
    exp_48_ram[2273] = 34;
    exp_48_ram[2274] = 39;
    exp_48_ram[2275] = 39;
    exp_48_ram[2276] = 37;
    exp_48_ram[2277] = 37;
    exp_48_ram[2278] = 6;
    exp_48_ram[2279] = 8;
    exp_48_ram[2280] = 56;
    exp_48_ram[2281] = 134;
    exp_48_ram[2282] = 135;
    exp_48_ram[2283] = 134;
    exp_48_ram[2284] = 7;
    exp_48_ram[2285] = 135;
    exp_48_ram[2286] = 5;
    exp_48_ram[2287] = 133;
    exp_48_ram[2288] = 224;
    exp_48_ram[2289] = 7;
    exp_48_ram[2290] = 135;
    exp_48_ram[2291] = 5;
    exp_48_ram[2292] = 133;
    exp_48_ram[2293] = 32;
    exp_48_ram[2294] = 36;
    exp_48_ram[2295] = 1;
    exp_48_ram[2296] = 128;
    exp_48_ram[2297] = 1;
    exp_48_ram[2298] = 46;
    exp_48_ram[2299] = 4;
    exp_48_ram[2300] = 38;
    exp_48_ram[2301] = 39;
    exp_48_ram[2302] = 247;
    exp_48_ram[2303] = 150;
    exp_48_ram[2304] = 39;
    exp_48_ram[2305] = 7;
    exp_48_ram[2306] = 119;
    exp_48_ram[2307] = 154;
    exp_48_ram[2308] = 39;
    exp_48_ram[2309] = 7;
    exp_48_ram[2310] = 119;
    exp_48_ram[2311] = 150;
    exp_48_ram[2312] = 7;
    exp_48_ram[2313] = 0;
    exp_48_ram[2314] = 7;
    exp_48_ram[2315] = 133;
    exp_48_ram[2316] = 36;
    exp_48_ram[2317] = 1;
    exp_48_ram[2318] = 128;
    exp_48_ram[2319] = 1;
    exp_48_ram[2320] = 46;
    exp_48_ram[2321] = 44;
    exp_48_ram[2322] = 4;
    exp_48_ram[2323] = 38;
    exp_48_ram[2324] = 37;
    exp_48_ram[2325] = 240;
    exp_48_ram[2326] = 7;
    exp_48_ram[2327] = 134;
    exp_48_ram[2328] = 7;
    exp_48_ram[2329] = 0;
    exp_48_ram[2330] = 7;
    exp_48_ram[2331] = 133;
    exp_48_ram[2332] = 32;
    exp_48_ram[2333] = 36;
    exp_48_ram[2334] = 1;
    exp_48_ram[2335] = 128;
    exp_48_ram[2336] = 1;
    exp_48_ram[2337] = 46;
    exp_48_ram[2338] = 44;
    exp_48_ram[2339] = 4;
    exp_48_ram[2340] = 38;
    exp_48_ram[2341] = 36;
    exp_48_ram[2342] = 39;
    exp_48_ram[2343] = 7;
    exp_48_ram[2344] = 4;
    exp_48_ram[2345] = 39;
    exp_48_ram[2346] = 7;
    exp_48_ram[2347] = 14;
    exp_48_ram[2348] = 39;
    exp_48_ram[2349] = 7;
    exp_48_ram[2350] = 8;
    exp_48_ram[2351] = 39;
    exp_48_ram[2352] = 7;
    exp_48_ram[2353] = 22;
    exp_48_ram[2354] = 7;
    exp_48_ram[2355] = 0;
    exp_48_ram[2356] = 39;
    exp_48_ram[2357] = 7;
    exp_48_ram[2358] = 18;
    exp_48_ram[2359] = 37;
    exp_48_ram[2360] = 240;
    exp_48_ram[2361] = 7;
    exp_48_ram[2362] = 134;
    exp_48_ram[2363] = 7;
    exp_48_ram[2364] = 0;
    exp_48_ram[2365] = 7;
    exp_48_ram[2366] = 0;
    exp_48_ram[2367] = 7;
    exp_48_ram[2368] = 133;
    exp_48_ram[2369] = 32;
    exp_48_ram[2370] = 36;
    exp_48_ram[2371] = 1;
    exp_48_ram[2372] = 128;
    exp_48_ram[2373] = 1;
    exp_48_ram[2374] = 38;
    exp_48_ram[2375] = 36;
    exp_48_ram[2376] = 34;
    exp_48_ram[2377] = 32;
    exp_48_ram[2378] = 46;
    exp_48_ram[2379] = 44;
    exp_48_ram[2380] = 42;
    exp_48_ram[2381] = 40;
    exp_48_ram[2382] = 38;
    exp_48_ram[2383] = 36;
    exp_48_ram[2384] = 34;
    exp_48_ram[2385] = 32;
    exp_48_ram[2386] = 46;
    exp_48_ram[2387] = 4;
    exp_48_ram[2388] = 4;
    exp_48_ram[2389] = 7;
    exp_48_ram[2390] = 8;
    exp_48_ram[2391] = 44;
    exp_48_ram[2392] = 46;
    exp_48_ram[2393] = 7;
    exp_48_ram[2394] = 42;
    exp_48_ram[2395] = 167;
    exp_48_ram[2396] = 38;
    exp_48_ram[2397] = 39;
    exp_48_ram[2398] = 135;
    exp_48_ram[2399] = 39;
    exp_48_ram[2400] = 6;
    exp_48_ram[2401] = 37;
    exp_48_ram[2402] = 240;
    exp_48_ram[2403] = 7;
    exp_48_ram[2404] = 87;
    exp_48_ram[2405] = 135;
    exp_48_ram[2406] = 7;
    exp_48_ram[2407] = 44;
    exp_48_ram[2408] = 46;
    exp_48_ram[2409] = 38;
    exp_48_ram[2410] = 38;
    exp_48_ram[2411] = 40;
    exp_48_ram[2412] = 40;
    exp_48_ram[2413] = 5;
    exp_48_ram[2414] = 7;
    exp_48_ram[2415] = 5;
    exp_48_ram[2416] = 181;
    exp_48_ram[2417] = 133;
    exp_48_ram[2418] = 135;
    exp_48_ram[2419] = 134;
    exp_48_ram[2420] = 135;
    exp_48_ram[2421] = 44;
    exp_48_ram[2422] = 46;
    exp_48_ram[2423] = 39;
    exp_48_ram[2424] = 135;
    exp_48_ram[2425] = 42;
    exp_48_ram[2426] = 240;
    exp_48_ram[2427] = 0;
    exp_48_ram[2428] = 40;
    exp_48_ram[2429] = 167;
    exp_48_ram[2430] = 135;
    exp_48_ram[2431] = 39;
    exp_48_ram[2432] = 128;
    exp_48_ram[2433] = 37;
    exp_48_ram[2434] = 37;
    exp_48_ram[2435] = 240;
    exp_48_ram[2436] = 7;
    exp_48_ram[2437] = 87;
    exp_48_ram[2438] = 135;
    exp_48_ram[2439] = 7;
    exp_48_ram[2440] = 141;
    exp_48_ram[2441] = 13;
    exp_48_ram[2442] = 38;
    exp_48_ram[2443] = 38;
    exp_48_ram[2444] = 7;
    exp_48_ram[2445] = 5;
    exp_48_ram[2446] = 181;
    exp_48_ram[2447] = 135;
    exp_48_ram[2448] = 134;
    exp_48_ram[2449] = 135;
    exp_48_ram[2450] = 44;
    exp_48_ram[2451] = 46;
    exp_48_ram[2452] = 39;
    exp_48_ram[2453] = 135;
    exp_48_ram[2454] = 40;
    exp_48_ram[2455] = 240;
    exp_48_ram[2456] = 0;
    exp_48_ram[2457] = 167;
    exp_48_ram[2458] = 135;
    exp_48_ram[2459] = 87;
    exp_48_ram[2460] = 135;
    exp_48_ram[2461] = 7;
    exp_48_ram[2462] = 140;
    exp_48_ram[2463] = 215;
    exp_48_ram[2464] = 140;
    exp_48_ram[2465] = 38;
    exp_48_ram[2466] = 38;
    exp_48_ram[2467] = 7;
    exp_48_ram[2468] = 5;
    exp_48_ram[2469] = 181;
    exp_48_ram[2470] = 135;
    exp_48_ram[2471] = 134;
    exp_48_ram[2472] = 135;
    exp_48_ram[2473] = 44;
    exp_48_ram[2474] = 46;
    exp_48_ram[2475] = 167;
    exp_48_ram[2476] = 23;
    exp_48_ram[2477] = 135;
    exp_48_ram[2478] = 7;
    exp_48_ram[2479] = 139;
    exp_48_ram[2480] = 215;
    exp_48_ram[2481] = 139;
    exp_48_ram[2482] = 38;
    exp_48_ram[2483] = 38;
    exp_48_ram[2484] = 7;
    exp_48_ram[2485] = 5;
    exp_48_ram[2486] = 181;
    exp_48_ram[2487] = 135;
    exp_48_ram[2488] = 134;
    exp_48_ram[2489] = 135;
    exp_48_ram[2490] = 44;
    exp_48_ram[2491] = 46;
    exp_48_ram[2492] = 167;
    exp_48_ram[2493] = 7;
    exp_48_ram[2494] = 151;
    exp_48_ram[2495] = 135;
    exp_48_ram[2496] = 151;
    exp_48_ram[2497] = 138;
    exp_48_ram[2498] = 215;
    exp_48_ram[2499] = 138;
    exp_48_ram[2500] = 38;
    exp_48_ram[2501] = 38;
    exp_48_ram[2502] = 7;
    exp_48_ram[2503] = 5;
    exp_48_ram[2504] = 181;
    exp_48_ram[2505] = 135;
    exp_48_ram[2506] = 134;
    exp_48_ram[2507] = 135;
    exp_48_ram[2508] = 44;
    exp_48_ram[2509] = 46;
    exp_48_ram[2510] = 167;
    exp_48_ram[2511] = 137;
    exp_48_ram[2512] = 215;
    exp_48_ram[2513] = 137;
    exp_48_ram[2514] = 38;
    exp_48_ram[2515] = 38;
    exp_48_ram[2516] = 7;
    exp_48_ram[2517] = 5;
    exp_48_ram[2518] = 181;
    exp_48_ram[2519] = 135;
    exp_48_ram[2520] = 134;
    exp_48_ram[2521] = 135;
    exp_48_ram[2522] = 44;
    exp_48_ram[2523] = 46;
    exp_48_ram[2524] = 39;
    exp_48_ram[2525] = 39;
    exp_48_ram[2526] = 5;
    exp_48_ram[2527] = 133;
    exp_48_ram[2528] = 32;
    exp_48_ram[2529] = 36;
    exp_48_ram[2530] = 36;
    exp_48_ram[2531] = 41;
    exp_48_ram[2532] = 41;
    exp_48_ram[2533] = 42;
    exp_48_ram[2534] = 42;
    exp_48_ram[2535] = 43;
    exp_48_ram[2536] = 43;
    exp_48_ram[2537] = 44;
    exp_48_ram[2538] = 44;
    exp_48_ram[2539] = 45;
    exp_48_ram[2540] = 45;
    exp_48_ram[2541] = 1;
    exp_48_ram[2542] = 128;
    exp_48_ram[2543] = 1;
    exp_48_ram[2544] = 46;
    exp_48_ram[2545] = 44;
    exp_48_ram[2546] = 42;
    exp_48_ram[2547] = 40;
    exp_48_ram[2548] = 38;
    exp_48_ram[2549] = 4;
    exp_48_ram[2550] = 46;
    exp_48_ram[2551] = 39;
    exp_48_ram[2552] = 163;
    exp_48_ram[2553] = 168;
    exp_48_ram[2554] = 168;
    exp_48_ram[2555] = 165;
    exp_48_ram[2556] = 165;
    exp_48_ram[2557] = 166;
    exp_48_ram[2558] = 166;
    exp_48_ram[2559] = 167;
    exp_48_ram[2560] = 167;
    exp_48_ram[2561] = 38;
    exp_48_ram[2562] = 40;
    exp_48_ram[2563] = 42;
    exp_48_ram[2564] = 44;
    exp_48_ram[2565] = 46;
    exp_48_ram[2566] = 32;
    exp_48_ram[2567] = 34;
    exp_48_ram[2568] = 36;
    exp_48_ram[2569] = 38;
    exp_48_ram[2570] = 35;
    exp_48_ram[2571] = 40;
    exp_48_ram[2572] = 40;
    exp_48_ram[2573] = 37;
    exp_48_ram[2574] = 37;
    exp_48_ram[2575] = 38;
    exp_48_ram[2576] = 38;
    exp_48_ram[2577] = 39;
    exp_48_ram[2578] = 39;
    exp_48_ram[2579] = 32;
    exp_48_ram[2580] = 34;
    exp_48_ram[2581] = 36;
    exp_48_ram[2582] = 38;
    exp_48_ram[2583] = 40;
    exp_48_ram[2584] = 42;
    exp_48_ram[2585] = 44;
    exp_48_ram[2586] = 46;
    exp_48_ram[2587] = 32;
    exp_48_ram[2588] = 7;
    exp_48_ram[2589] = 133;
    exp_48_ram[2590] = 240;
    exp_48_ram[2591] = 40;
    exp_48_ram[2592] = 42;
    exp_48_ram[2593] = 39;
    exp_48_ram[2594] = 94;
    exp_48_ram[2595] = 38;
    exp_48_ram[2596] = 38;
    exp_48_ram[2597] = 245;
    exp_48_ram[2598] = 5;
    exp_48_ram[2599] = 5;
    exp_48_ram[2600] = 7;
    exp_48_ram[2601] = 8;
    exp_48_ram[2602] = 56;
    exp_48_ram[2603] = 135;
    exp_48_ram[2604] = 6;
    exp_48_ram[2605] = 135;
    exp_48_ram[2606] = 44;
    exp_48_ram[2607] = 46;
    exp_48_ram[2608] = 0;
    exp_48_ram[2609] = 39;
    exp_48_ram[2610] = 210;
    exp_48_ram[2611] = 35;
    exp_48_ram[2612] = 40;
    exp_48_ram[2613] = 40;
    exp_48_ram[2614] = 37;
    exp_48_ram[2615] = 37;
    exp_48_ram[2616] = 38;
    exp_48_ram[2617] = 38;
    exp_48_ram[2618] = 39;
    exp_48_ram[2619] = 39;
    exp_48_ram[2620] = 32;
    exp_48_ram[2621] = 34;
    exp_48_ram[2622] = 36;
    exp_48_ram[2623] = 38;
    exp_48_ram[2624] = 40;
    exp_48_ram[2625] = 42;
    exp_48_ram[2626] = 44;
    exp_48_ram[2627] = 46;
    exp_48_ram[2628] = 32;
    exp_48_ram[2629] = 7;
    exp_48_ram[2630] = 133;
    exp_48_ram[2631] = 240;
    exp_48_ram[2632] = 7;
    exp_48_ram[2633] = 138;
    exp_48_ram[2634] = 22;
    exp_48_ram[2635] = 6;
    exp_48_ram[2636] = 6;
    exp_48_ram[2637] = 0;
    exp_48_ram[2638] = 6;
    exp_48_ram[2639] = 6;
    exp_48_ram[2640] = 37;
    exp_48_ram[2641] = 37;
    exp_48_ram[2642] = 7;
    exp_48_ram[2643] = 8;
    exp_48_ram[2644] = 56;
    exp_48_ram[2645] = 135;
    exp_48_ram[2646] = 134;
    exp_48_ram[2647] = 135;
    exp_48_ram[2648] = 44;
    exp_48_ram[2649] = 46;
    exp_48_ram[2650] = 0;
    exp_48_ram[2651] = 39;
    exp_48_ram[2652] = 39;
    exp_48_ram[2653] = 44;
    exp_48_ram[2654] = 46;
    exp_48_ram[2655] = 71;
    exp_48_ram[2656] = 167;
    exp_48_ram[2657] = 137;
    exp_48_ram[2658] = 215;
    exp_48_ram[2659] = 137;
    exp_48_ram[2660] = 38;
    exp_48_ram[2661] = 38;
    exp_48_ram[2662] = 7;
    exp_48_ram[2663] = 5;
    exp_48_ram[2664] = 53;
    exp_48_ram[2665] = 135;
    exp_48_ram[2666] = 134;
    exp_48_ram[2667] = 135;
    exp_48_ram[2668] = 44;
    exp_48_ram[2669] = 46;
    exp_48_ram[2670] = 36;
    exp_48_ram[2671] = 7;
    exp_48_ram[2672] = 37;
    exp_48_ram[2673] = 38;
    exp_48_ram[2674] = 133;
    exp_48_ram[2675] = 0;
    exp_48_ram[2676] = 35;
    exp_48_ram[2677] = 40;
    exp_48_ram[2678] = 40;
    exp_48_ram[2679] = 37;
    exp_48_ram[2680] = 37;
    exp_48_ram[2681] = 38;
    exp_48_ram[2682] = 38;
    exp_48_ram[2683] = 39;
    exp_48_ram[2684] = 39;
    exp_48_ram[2685] = 160;
    exp_48_ram[2686] = 162;
    exp_48_ram[2687] = 164;
    exp_48_ram[2688] = 166;
    exp_48_ram[2689] = 168;
    exp_48_ram[2690] = 170;
    exp_48_ram[2691] = 172;
    exp_48_ram[2692] = 174;
    exp_48_ram[2693] = 160;
    exp_48_ram[2694] = 39;
    exp_48_ram[2695] = 90;
    exp_48_ram[2696] = 39;
    exp_48_ram[2697] = 7;
    exp_48_ram[2698] = 160;
    exp_48_ram[2699] = 0;
    exp_48_ram[2700] = 39;
    exp_48_ram[2701] = 212;
    exp_48_ram[2702] = 35;
    exp_48_ram[2703] = 40;
    exp_48_ram[2704] = 40;
    exp_48_ram[2705] = 37;
    exp_48_ram[2706] = 37;
    exp_48_ram[2707] = 38;
    exp_48_ram[2708] = 38;
    exp_48_ram[2709] = 39;
    exp_48_ram[2710] = 39;
    exp_48_ram[2711] = 32;
    exp_48_ram[2712] = 34;
    exp_48_ram[2713] = 36;
    exp_48_ram[2714] = 38;
    exp_48_ram[2715] = 40;
    exp_48_ram[2716] = 42;
    exp_48_ram[2717] = 44;
    exp_48_ram[2718] = 46;
    exp_48_ram[2719] = 32;
    exp_48_ram[2720] = 7;
    exp_48_ram[2721] = 133;
    exp_48_ram[2722] = 240;
    exp_48_ram[2723] = 7;
    exp_48_ram[2724] = 39;
    exp_48_ram[2725] = 160;
    exp_48_ram[2726] = 0;
    exp_48_ram[2727] = 39;
    exp_48_ram[2728] = 160;
    exp_48_ram[2729] = 39;
    exp_48_ram[2730] = 39;
    exp_48_ram[2731] = 5;
    exp_48_ram[2732] = 133;
    exp_48_ram[2733] = 32;
    exp_48_ram[2734] = 36;
    exp_48_ram[2735] = 36;
    exp_48_ram[2736] = 41;
    exp_48_ram[2737] = 41;
    exp_48_ram[2738] = 1;
    exp_48_ram[2739] = 128;
    exp_48_ram[2740] = 1;
    exp_48_ram[2741] = 46;
    exp_48_ram[2742] = 44;
    exp_48_ram[2743] = 42;
    exp_48_ram[2744] = 40;
    exp_48_ram[2745] = 38;
    exp_48_ram[2746] = 36;
    exp_48_ram[2747] = 34;
    exp_48_ram[2748] = 32;
    exp_48_ram[2749] = 4;
    exp_48_ram[2750] = 38;
    exp_48_ram[2751] = 240;
    exp_48_ram[2752] = 7;
    exp_48_ram[2753] = 135;
    exp_48_ram[2754] = 70;
    exp_48_ram[2755] = 166;
    exp_48_ram[2756] = 138;
    exp_48_ram[2757] = 10;
    exp_48_ram[2758] = 6;
    exp_48_ram[2759] = 134;
    exp_48_ram[2760] = 5;
    exp_48_ram[2761] = 133;
    exp_48_ram[2762] = 208;
    exp_48_ram[2763] = 7;
    exp_48_ram[2764] = 135;
    exp_48_ram[2765] = 46;
    exp_48_ram[2766] = 71;
    exp_48_ram[2767] = 167;
    exp_48_ram[2768] = 167;
    exp_48_ram[2769] = 39;
    exp_48_ram[2770] = 135;
    exp_48_ram[2771] = 46;
    exp_48_ram[2772] = 39;
    exp_48_ram[2773] = 142;
    exp_48_ram[2774] = 39;
    exp_48_ram[2775] = 137;
    exp_48_ram[2776] = 9;
    exp_48_ram[2777] = 39;
    exp_48_ram[2778] = 160;
    exp_48_ram[2779] = 162;
    exp_48_ram[2780] = 39;
    exp_48_ram[2781] = 139;
    exp_48_ram[2782] = 11;
    exp_48_ram[2783] = 7;
    exp_48_ram[2784] = 135;
    exp_48_ram[2785] = 5;
    exp_48_ram[2786] = 133;
    exp_48_ram[2787] = 32;
    exp_48_ram[2788] = 36;
    exp_48_ram[2789] = 41;
    exp_48_ram[2790] = 41;
    exp_48_ram[2791] = 42;
    exp_48_ram[2792] = 42;
    exp_48_ram[2793] = 43;
    exp_48_ram[2794] = 43;
    exp_48_ram[2795] = 1;
    exp_48_ram[2796] = 128;
    exp_48_ram[2797] = 1;
    exp_48_ram[2798] = 38;
    exp_48_ram[2799] = 36;
    exp_48_ram[2800] = 34;
    exp_48_ram[2801] = 32;
    exp_48_ram[2802] = 4;
    exp_48_ram[2803] = 44;
    exp_48_ram[2804] = 46;
    exp_48_ram[2805] = 240;
    exp_48_ram[2806] = 7;
    exp_48_ram[2807] = 135;
    exp_48_ram[2808] = 70;
    exp_48_ram[2809] = 166;
    exp_48_ram[2810] = 137;
    exp_48_ram[2811] = 9;
    exp_48_ram[2812] = 6;
    exp_48_ram[2813] = 134;
    exp_48_ram[2814] = 5;
    exp_48_ram[2815] = 133;
    exp_48_ram[2816] = 208;
    exp_48_ram[2817] = 7;
    exp_48_ram[2818] = 135;
    exp_48_ram[2819] = 36;
    exp_48_ram[2820] = 38;
    exp_48_ram[2821] = 39;
    exp_48_ram[2822] = 39;
    exp_48_ram[2823] = 37;
    exp_48_ram[2824] = 37;
    exp_48_ram[2825] = 6;
    exp_48_ram[2826] = 8;
    exp_48_ram[2827] = 56;
    exp_48_ram[2828] = 134;
    exp_48_ram[2829] = 135;
    exp_48_ram[2830] = 134;
    exp_48_ram[2831] = 7;
    exp_48_ram[2832] = 135;
    exp_48_ram[2833] = 70;
    exp_48_ram[2834] = 164;
    exp_48_ram[2835] = 166;
    exp_48_ram[2836] = 0;
    exp_48_ram[2837] = 32;
    exp_48_ram[2838] = 36;
    exp_48_ram[2839] = 41;
    exp_48_ram[2840] = 41;
    exp_48_ram[2841] = 1;
    exp_48_ram[2842] = 128;
    exp_48_ram[2843] = 1;
    exp_48_ram[2844] = 38;
    exp_48_ram[2845] = 36;
    exp_48_ram[2846] = 4;
    exp_48_ram[2847] = 46;
    exp_48_ram[2848] = 23;
    exp_48_ram[2849] = 135;
    exp_48_ram[2850] = 165;
    exp_48_ram[2851] = 165;
    exp_48_ram[2852] = 166;
    exp_48_ram[2853] = 166;
    exp_48_ram[2854] = 167;
    exp_48_ram[2855] = 42;
    exp_48_ram[2856] = 44;
    exp_48_ram[2857] = 46;
    exp_48_ram[2858] = 32;
    exp_48_ram[2859] = 34;
    exp_48_ram[2860] = 215;
    exp_48_ram[2861] = 20;
    exp_48_ram[2862] = 23;
    exp_48_ram[2863] = 135;
    exp_48_ram[2864] = 174;
    exp_48_ram[2865] = 163;
    exp_48_ram[2866] = 168;
    exp_48_ram[2867] = 168;
    exp_48_ram[2868] = 165;
    exp_48_ram[2869] = 165;
    exp_48_ram[2870] = 166;
    exp_48_ram[2871] = 166;
    exp_48_ram[2872] = 167;
    exp_48_ram[2873] = 38;
    exp_48_ram[2874] = 40;
    exp_48_ram[2875] = 42;
    exp_48_ram[2876] = 44;
    exp_48_ram[2877] = 46;
    exp_48_ram[2878] = 32;
    exp_48_ram[2879] = 34;
    exp_48_ram[2880] = 36;
    exp_48_ram[2881] = 38;
    exp_48_ram[2882] = 199;
    exp_48_ram[2883] = 8;
    exp_48_ram[2884] = 38;
    exp_48_ram[2885] = 0;
    exp_48_ram[2886] = 39;
    exp_48_ram[2887] = 167;
    exp_48_ram[2888] = 7;
    exp_48_ram[2889] = 151;
    exp_48_ram[2890] = 135;
    exp_48_ram[2891] = 39;
    exp_48_ram[2892] = 7;
    exp_48_ram[2893] = 7;
    exp_48_ram[2894] = 7;
    exp_48_ram[2895] = 199;
    exp_48_ram[2896] = 71;
    exp_48_ram[2897] = 134;
    exp_48_ram[2898] = 39;
    exp_48_ram[2899] = 135;
    exp_48_ram[2900] = 128;
    exp_48_ram[2901] = 39;
    exp_48_ram[2902] = 135;
    exp_48_ram[2903] = 38;
    exp_48_ram[2904] = 39;
    exp_48_ram[2905] = 7;
    exp_48_ram[2906] = 216;
    exp_48_ram[2907] = 71;
    exp_48_ram[2908] = 135;
    exp_48_ram[2909] = 7;
    exp_48_ram[2910] = 129;
    exp_48_ram[2911] = 38;
    exp_48_ram[2912] = 0;
    exp_48_ram[2913] = 39;
    exp_48_ram[2914] = 167;
    exp_48_ram[2915] = 7;
    exp_48_ram[2916] = 151;
    exp_48_ram[2917] = 135;
    exp_48_ram[2918] = 39;
    exp_48_ram[2919] = 7;
    exp_48_ram[2920] = 39;
    exp_48_ram[2921] = 135;
    exp_48_ram[2922] = 6;
    exp_48_ram[2923] = 135;
    exp_48_ram[2924] = 71;
    exp_48_ram[2925] = 70;
    exp_48_ram[2926] = 134;
    exp_48_ram[2927] = 135;
    exp_48_ram[2928] = 128;
    exp_48_ram[2929] = 39;
    exp_48_ram[2930] = 135;
    exp_48_ram[2931] = 38;
    exp_48_ram[2932] = 39;
    exp_48_ram[2933] = 7;
    exp_48_ram[2934] = 214;
    exp_48_ram[2935] = 71;
    exp_48_ram[2936] = 135;
    exp_48_ram[2937] = 7;
    exp_48_ram[2938] = 131;
    exp_48_ram[2939] = 39;
    exp_48_ram[2940] = 167;
    exp_48_ram[2941] = 5;
    exp_48_ram[2942] = 133;
    exp_48_ram[2943] = 16;
    exp_48_ram[2944] = 7;
    exp_48_ram[2945] = 135;
    exp_48_ram[2946] = 34;
    exp_48_ram[2947] = 36;
    exp_48_ram[2948] = 39;
    exp_48_ram[2949] = 247;
    exp_48_ram[2950] = 135;
    exp_48_ram[2951] = 247;
    exp_48_ram[2952] = 71;
    exp_48_ram[2953] = 135;
    exp_48_ram[2954] = 132;
    exp_48_ram[2955] = 39;
    exp_48_ram[2956] = 247;
    exp_48_ram[2957] = 135;
    exp_48_ram[2958] = 247;
    exp_48_ram[2959] = 71;
    exp_48_ram[2960] = 135;
    exp_48_ram[2961] = 132;
    exp_48_ram[2962] = 71;
    exp_48_ram[2963] = 135;
    exp_48_ram[2964] = 7;
    exp_48_ram[2965] = 133;
    exp_48_ram[2966] = 39;
    exp_48_ram[2967] = 167;
    exp_48_ram[2968] = 5;
    exp_48_ram[2969] = 133;
    exp_48_ram[2970] = 16;
    exp_48_ram[2971] = 7;
    exp_48_ram[2972] = 135;
    exp_48_ram[2973] = 34;
    exp_48_ram[2974] = 36;
    exp_48_ram[2975] = 39;
    exp_48_ram[2976] = 247;
    exp_48_ram[2977] = 135;
    exp_48_ram[2978] = 247;
    exp_48_ram[2979] = 71;
    exp_48_ram[2980] = 135;
    exp_48_ram[2981] = 133;
    exp_48_ram[2982] = 39;
    exp_48_ram[2983] = 247;
    exp_48_ram[2984] = 135;
    exp_48_ram[2985] = 247;
    exp_48_ram[2986] = 71;
    exp_48_ram[2987] = 135;
    exp_48_ram[2988] = 134;
    exp_48_ram[2989] = 71;
    exp_48_ram[2990] = 135;
    exp_48_ram[2991] = 7;
    exp_48_ram[2992] = 134;
    exp_48_ram[2993] = 39;
    exp_48_ram[2994] = 167;
    exp_48_ram[2995] = 5;
    exp_48_ram[2996] = 133;
    exp_48_ram[2997] = 16;
    exp_48_ram[2998] = 7;
    exp_48_ram[2999] = 135;
    exp_48_ram[3000] = 34;
    exp_48_ram[3001] = 36;
    exp_48_ram[3002] = 39;
    exp_48_ram[3003] = 247;
    exp_48_ram[3004] = 135;
    exp_48_ram[3005] = 247;
    exp_48_ram[3006] = 71;
    exp_48_ram[3007] = 135;
    exp_48_ram[3008] = 135;
    exp_48_ram[3009] = 39;
    exp_48_ram[3010] = 247;
    exp_48_ram[3011] = 135;
    exp_48_ram[3012] = 247;
    exp_48_ram[3013] = 71;
    exp_48_ram[3014] = 135;
    exp_48_ram[3015] = 135;
    exp_48_ram[3016] = 71;
    exp_48_ram[3017] = 135;
    exp_48_ram[3018] = 7;
    exp_48_ram[3019] = 136;
    exp_48_ram[3020] = 39;
    exp_48_ram[3021] = 167;
    exp_48_ram[3022] = 5;
    exp_48_ram[3023] = 133;
    exp_48_ram[3024] = 16;
    exp_48_ram[3025] = 7;
    exp_48_ram[3026] = 135;
    exp_48_ram[3027] = 34;
    exp_48_ram[3028] = 36;
    exp_48_ram[3029] = 39;
    exp_48_ram[3030] = 247;
    exp_48_ram[3031] = 135;
    exp_48_ram[3032] = 247;
    exp_48_ram[3033] = 71;
    exp_48_ram[3034] = 135;
    exp_48_ram[3035] = 136;
    exp_48_ram[3036] = 39;
    exp_48_ram[3037] = 247;
    exp_48_ram[3038] = 135;
    exp_48_ram[3039] = 247;
    exp_48_ram[3040] = 71;
    exp_48_ram[3041] = 135;
    exp_48_ram[3042] = 137;
    exp_48_ram[3043] = 71;
    exp_48_ram[3044] = 135;
    exp_48_ram[3045] = 7;
    exp_48_ram[3046] = 137;
    exp_48_ram[3047] = 39;
    exp_48_ram[3048] = 167;
    exp_48_ram[3049] = 135;
    exp_48_ram[3050] = 5;
    exp_48_ram[3051] = 133;
    exp_48_ram[3052] = 16;
    exp_48_ram[3053] = 7;
    exp_48_ram[3054] = 135;
    exp_48_ram[3055] = 34;
    exp_48_ram[3056] = 36;
    exp_48_ram[3057] = 39;
    exp_48_ram[3058] = 247;
    exp_48_ram[3059] = 135;
    exp_48_ram[3060] = 247;
    exp_48_ram[3061] = 71;
    exp_48_ram[3062] = 135;
    exp_48_ram[3063] = 138;
    exp_48_ram[3064] = 39;
    exp_48_ram[3065] = 5;
    exp_48_ram[3066] = 133;
    exp_48_ram[3067] = 16;
    exp_48_ram[3068] = 7;
    exp_48_ram[3069] = 135;
    exp_48_ram[3070] = 34;
    exp_48_ram[3071] = 36;
    exp_48_ram[3072] = 39;
    exp_48_ram[3073] = 247;
    exp_48_ram[3074] = 135;
    exp_48_ram[3075] = 247;
    exp_48_ram[3076] = 71;
    exp_48_ram[3077] = 135;
    exp_48_ram[3078] = 138;
    exp_48_ram[3079] = 39;
    exp_48_ram[3080] = 5;
    exp_48_ram[3081] = 133;
    exp_48_ram[3082] = 16;
    exp_48_ram[3083] = 7;
    exp_48_ram[3084] = 135;
    exp_48_ram[3085] = 34;
    exp_48_ram[3086] = 36;
    exp_48_ram[3087] = 39;
    exp_48_ram[3088] = 247;
    exp_48_ram[3089] = 135;
    exp_48_ram[3090] = 247;
    exp_48_ram[3091] = 71;
    exp_48_ram[3092] = 135;
    exp_48_ram[3093] = 139;
    exp_48_ram[3094] = 39;
    exp_48_ram[3095] = 247;
    exp_48_ram[3096] = 135;
    exp_48_ram[3097] = 247;
    exp_48_ram[3098] = 71;
    exp_48_ram[3099] = 135;
    exp_48_ram[3100] = 139;
    exp_48_ram[3101] = 71;
    exp_48_ram[3102] = 135;
    exp_48_ram[3103] = 7;
    exp_48_ram[3104] = 140;
    exp_48_ram[3105] = 71;
    exp_48_ram[3106] = 135;
    exp_48_ram[3107] = 140;
    exp_48_ram[3108] = 71;
    exp_48_ram[3109] = 135;
    exp_48_ram[3110] = 133;
    exp_48_ram[3111] = 32;
    exp_48_ram[3112] = 36;
    exp_48_ram[3113] = 1;
    exp_48_ram[3114] = 128;
    exp_48_ram[3115] = 1;
    exp_48_ram[3116] = 46;
    exp_48_ram[3117] = 44;
    exp_48_ram[3118] = 4;
    exp_48_ram[3119] = 38;
    exp_48_ram[3120] = 37;
    exp_48_ram[3121] = 0;
    exp_48_ram[3122] = 7;
    exp_48_ram[3123] = 133;
    exp_48_ram[3124] = 240;
    exp_48_ram[3125] = 7;
    exp_48_ram[3126] = 133;
    exp_48_ram[3127] = 32;
    exp_48_ram[3128] = 36;
    exp_48_ram[3129] = 1;
    exp_48_ram[3130] = 128;
    exp_48_ram[3131] = 1;
    exp_48_ram[3132] = 46;
    exp_48_ram[3133] = 44;
    exp_48_ram[3134] = 42;
    exp_48_ram[3135] = 40;
    exp_48_ram[3136] = 38;
    exp_48_ram[3137] = 36;
    exp_48_ram[3138] = 34;
    exp_48_ram[3139] = 32;
    exp_48_ram[3140] = 46;
    exp_48_ram[3141] = 44;
    exp_48_ram[3142] = 4;
    exp_48_ram[3143] = 38;
    exp_48_ram[3144] = 32;
    exp_48_ram[3145] = 34;
    exp_48_ram[3146] = 7;
    exp_48_ram[3147] = 44;
    exp_48_ram[3148] = 7;
    exp_48_ram[3149] = 46;
    exp_48_ram[3150] = 39;
    exp_48_ram[3151] = 133;
    exp_48_ram[3152] = 240;
    exp_48_ram[3153] = 38;
    exp_48_ram[3154] = 39;
    exp_48_ram[3155] = 87;
    exp_48_ram[3156] = 135;
    exp_48_ram[3157] = 7;
    exp_48_ram[3158] = 36;
    exp_48_ram[3159] = 39;
    exp_48_ram[3160] = 140;
    exp_48_ram[3161] = 12;
    exp_48_ram[3162] = 39;
    exp_48_ram[3163] = 135;
    exp_48_ram[3164] = 234;
    exp_48_ram[3165] = 39;
    exp_48_ram[3166] = 135;
    exp_48_ram[3167] = 152;
    exp_48_ram[3168] = 39;
    exp_48_ram[3169] = 7;
    exp_48_ram[3170] = 238;
    exp_48_ram[3171] = 39;
    exp_48_ram[3172] = 135;
    exp_48_ram[3173] = 44;
    exp_48_ram[3174] = 39;
    exp_48_ram[3175] = 135;
    exp_48_ram[3176] = 39;
    exp_48_ram[3177] = 7;
    exp_48_ram[3178] = 46;
    exp_48_ram[3179] = 39;
    exp_48_ram[3180] = 138;
    exp_48_ram[3181] = 10;
    exp_48_ram[3182] = 38;
    exp_48_ram[3183] = 38;
    exp_48_ram[3184] = 7;
    exp_48_ram[3185] = 5;
    exp_48_ram[3186] = 53;
    exp_48_ram[3187] = 135;
    exp_48_ram[3188] = 134;
    exp_48_ram[3189] = 135;
    exp_48_ram[3190] = 32;
    exp_48_ram[3191] = 34;
    exp_48_ram[3192] = 240;
    exp_48_ram[3193] = 0;
    exp_48_ram[3194] = 42;
    exp_48_ram[3195] = 32;
    exp_48_ram[3196] = 39;
    exp_48_ram[3197] = 135;
    exp_48_ram[3198] = 39;
    exp_48_ram[3199] = 133;
    exp_48_ram[3200] = 5;
    exp_48_ram[3201] = 240;
    exp_48_ram[3202] = 38;
    exp_48_ram[3203] = 39;
    exp_48_ram[3204] = 87;
    exp_48_ram[3205] = 135;
    exp_48_ram[3206] = 7;
    exp_48_ram[3207] = 36;
    exp_48_ram[3208] = 39;
    exp_48_ram[3209] = 139;
    exp_48_ram[3210] = 11;
    exp_48_ram[3211] = 39;
    exp_48_ram[3212] = 135;
    exp_48_ram[3213] = 228;
    exp_48_ram[3214] = 39;
    exp_48_ram[3215] = 135;
    exp_48_ram[3216] = 152;
    exp_48_ram[3217] = 39;
    exp_48_ram[3218] = 7;
    exp_48_ram[3219] = 232;
    exp_48_ram[3220] = 39;
    exp_48_ram[3221] = 135;
    exp_48_ram[3222] = 42;
    exp_48_ram[3223] = 39;
    exp_48_ram[3224] = 135;
    exp_48_ram[3225] = 39;
    exp_48_ram[3226] = 7;
    exp_48_ram[3227] = 46;
    exp_48_ram[3228] = 39;
    exp_48_ram[3229] = 135;
    exp_48_ram[3230] = 39;
    exp_48_ram[3231] = 7;
    exp_48_ram[3232] = 32;
    exp_48_ram[3233] = 39;
    exp_48_ram[3234] = 137;
    exp_48_ram[3235] = 9;
    exp_48_ram[3236] = 38;
    exp_48_ram[3237] = 38;
    exp_48_ram[3238] = 7;
    exp_48_ram[3239] = 5;
    exp_48_ram[3240] = 53;
    exp_48_ram[3241] = 135;
    exp_48_ram[3242] = 134;
    exp_48_ram[3243] = 135;
    exp_48_ram[3244] = 32;
    exp_48_ram[3245] = 34;
    exp_48_ram[3246] = 240;
    exp_48_ram[3247] = 0;
    exp_48_ram[3248] = 39;
    exp_48_ram[3249] = 135;
    exp_48_ram[3250] = 44;
    exp_48_ram[3251] = 39;
    exp_48_ram[3252] = 87;
    exp_48_ram[3253] = 133;
    exp_48_ram[3254] = 5;
    exp_48_ram[3255] = 0;
    exp_48_ram[3256] = 7;
    exp_48_ram[3257] = 135;
    exp_48_ram[3258] = 46;
    exp_48_ram[3259] = 32;
    exp_48_ram[3260] = 39;
    exp_48_ram[3261] = 135;
    exp_48_ram[3262] = 40;
    exp_48_ram[3263] = 39;
    exp_48_ram[3264] = 39;
    exp_48_ram[3265] = 7;
    exp_48_ram[3266] = 46;
    exp_48_ram[3267] = 39;
    exp_48_ram[3268] = 7;
    exp_48_ram[3269] = 103;
    exp_48_ram[3270] = 46;
    exp_48_ram[3271] = 39;
    exp_48_ram[3272] = 39;
    exp_48_ram[3273] = 7;
    exp_48_ram[3274] = 32;
    exp_48_ram[3275] = 39;
    exp_48_ram[3276] = 32;
    exp_48_ram[3277] = 215;
    exp_48_ram[3278] = 34;
    exp_48_ram[3279] = 39;
    exp_48_ram[3280] = 23;
    exp_48_ram[3281] = 133;
    exp_48_ram[3282] = 5;
    exp_48_ram[3283] = 0;
    exp_48_ram[3284] = 7;
    exp_48_ram[3285] = 135;
    exp_48_ram[3286] = 46;
    exp_48_ram[3287] = 32;
    exp_48_ram[3288] = 39;
    exp_48_ram[3289] = 38;
    exp_48_ram[3290] = 39;
    exp_48_ram[3291] = 32;
    exp_48_ram[3292] = 215;
    exp_48_ram[3293] = 34;
    exp_48_ram[3294] = 39;
    exp_48_ram[3295] = 5;
    exp_48_ram[3296] = 133;
    exp_48_ram[3297] = 0;
    exp_48_ram[3298] = 7;
    exp_48_ram[3299] = 135;
    exp_48_ram[3300] = 46;
    exp_48_ram[3301] = 32;
    exp_48_ram[3302] = 39;
    exp_48_ram[3303] = 36;
    exp_48_ram[3304] = 39;
    exp_48_ram[3305] = 32;
    exp_48_ram[3306] = 215;
    exp_48_ram[3307] = 34;
    exp_48_ram[3308] = 39;
    exp_48_ram[3309] = 34;
    exp_48_ram[3310] = 39;
    exp_48_ram[3311] = 46;
    exp_48_ram[3312] = 35;
    exp_48_ram[3313] = 40;
    exp_48_ram[3314] = 40;
    exp_48_ram[3315] = 37;
    exp_48_ram[3316] = 37;
    exp_48_ram[3317] = 38;
    exp_48_ram[3318] = 38;
    exp_48_ram[3319] = 39;
    exp_48_ram[3320] = 160;
    exp_48_ram[3321] = 162;
    exp_48_ram[3322] = 164;
    exp_48_ram[3323] = 166;
    exp_48_ram[3324] = 168;
    exp_48_ram[3325] = 170;
    exp_48_ram[3326] = 172;
    exp_48_ram[3327] = 174;
    exp_48_ram[3328] = 160;
    exp_48_ram[3329] = 37;
    exp_48_ram[3330] = 32;
    exp_48_ram[3331] = 36;
    exp_48_ram[3332] = 41;
    exp_48_ram[3333] = 41;
    exp_48_ram[3334] = 42;
    exp_48_ram[3335] = 42;
    exp_48_ram[3336] = 43;
    exp_48_ram[3337] = 43;
    exp_48_ram[3338] = 44;
    exp_48_ram[3339] = 44;
    exp_48_ram[3340] = 1;
    exp_48_ram[3341] = 128;
    exp_48_ram[3342] = 1;
    exp_48_ram[3343] = 46;
    exp_48_ram[3344] = 44;
    exp_48_ram[3345] = 42;
    exp_48_ram[3346] = 40;
    exp_48_ram[3347] = 38;
    exp_48_ram[3348] = 4;
    exp_48_ram[3349] = 46;
    exp_48_ram[3350] = 7;
    exp_48_ram[3351] = 8;
    exp_48_ram[3352] = 44;
    exp_48_ram[3353] = 46;
    exp_48_ram[3354] = 39;
    exp_48_ram[3355] = 167;
    exp_48_ram[3356] = 167;
    exp_48_ram[3357] = 40;
    exp_48_ram[3358] = 42;
    exp_48_ram[3359] = 37;
    exp_48_ram[3360] = 37;
    exp_48_ram[3361] = 224;
    exp_48_ram[3362] = 7;
    exp_48_ram[3363] = 140;
    exp_48_ram[3364] = 23;
    exp_48_ram[3365] = 7;
    exp_48_ram[3366] = 7;
    exp_48_ram[3367] = 44;
    exp_48_ram[3368] = 46;
    exp_48_ram[3369] = 71;
    exp_48_ram[3370] = 167;
    exp_48_ram[3371] = 137;
    exp_48_ram[3372] = 215;
    exp_48_ram[3373] = 137;
    exp_48_ram[3374] = 38;
    exp_48_ram[3375] = 38;
    exp_48_ram[3376] = 7;
    exp_48_ram[3377] = 5;
    exp_48_ram[3378] = 181;
    exp_48_ram[3379] = 135;
    exp_48_ram[3380] = 134;
    exp_48_ram[3381] = 135;
    exp_48_ram[3382] = 5;
    exp_48_ram[3383] = 133;
    exp_48_ram[3384] = 38;
    exp_48_ram[3385] = 38;
    exp_48_ram[3386] = 7;
    exp_48_ram[3387] = 8;
    exp_48_ram[3388] = 56;
    exp_48_ram[3389] = 135;
    exp_48_ram[3390] = 6;
    exp_48_ram[3391] = 135;
    exp_48_ram[3392] = 36;
    exp_48_ram[3393] = 38;
    exp_48_ram[3394] = 71;
    exp_48_ram[3395] = 132;
    exp_48_ram[3396] = 7;
    exp_48_ram[3397] = 37;
    exp_48_ram[3398] = 38;
    exp_48_ram[3399] = 133;
    exp_48_ram[3400] = 240;
    exp_48_ram[3401] = 35;
    exp_48_ram[3402] = 40;
    exp_48_ram[3403] = 40;
    exp_48_ram[3404] = 37;
    exp_48_ram[3405] = 37;
    exp_48_ram[3406] = 38;
    exp_48_ram[3407] = 38;
    exp_48_ram[3408] = 39;
    exp_48_ram[3409] = 39;
    exp_48_ram[3410] = 160;
    exp_48_ram[3411] = 162;
    exp_48_ram[3412] = 164;
    exp_48_ram[3413] = 166;
    exp_48_ram[3414] = 168;
    exp_48_ram[3415] = 170;
    exp_48_ram[3416] = 172;
    exp_48_ram[3417] = 174;
    exp_48_ram[3418] = 160;
    exp_48_ram[3419] = 37;
    exp_48_ram[3420] = 37;
    exp_48_ram[3421] = 224;
    exp_48_ram[3422] = 7;
    exp_48_ram[3423] = 71;
    exp_48_ram[3424] = 135;
    exp_48_ram[3425] = 160;
    exp_48_ram[3426] = 71;
    exp_48_ram[3427] = 135;
    exp_48_ram[3428] = 133;
    exp_48_ram[3429] = 32;
    exp_48_ram[3430] = 36;
    exp_48_ram[3431] = 36;
    exp_48_ram[3432] = 41;
    exp_48_ram[3433] = 41;
    exp_48_ram[3434] = 1;
    exp_48_ram[3435] = 128;
    exp_48_ram[3436] = 1;
    exp_48_ram[3437] = 38;
    exp_48_ram[3438] = 36;
    exp_48_ram[3439] = 4;
    exp_48_ram[3440] = 46;
    exp_48_ram[3441] = 38;
    exp_48_ram[3442] = 37;
    exp_48_ram[3443] = 208;
    exp_48_ram[3444] = 7;
    exp_48_ram[3445] = 5;
    exp_48_ram[3446] = 71;
    exp_48_ram[3447] = 135;
    exp_48_ram[3448] = 7;
    exp_48_ram[3449] = 234;
    exp_48_ram[3450] = 39;
    exp_48_ram[3451] = 7;
    exp_48_ram[3452] = 151;
    exp_48_ram[3453] = 135;
    exp_48_ram[3454] = 151;
    exp_48_ram[3455] = 38;
    exp_48_ram[3456] = 71;
    exp_48_ram[3457] = 39;
    exp_48_ram[3458] = 7;
    exp_48_ram[3459] = 135;
    exp_48_ram[3460] = 38;
    exp_48_ram[3461] = 240;
    exp_48_ram[3462] = 0;
    exp_48_ram[3463] = 39;
    exp_48_ram[3464] = 133;
    exp_48_ram[3465] = 32;
    exp_48_ram[3466] = 36;
    exp_48_ram[3467] = 1;
    exp_48_ram[3468] = 128;
    exp_48_ram[3469] = 1;
    exp_48_ram[3470] = 38;
    exp_48_ram[3471] = 36;
    exp_48_ram[3472] = 4;
    exp_48_ram[3473] = 71;
    exp_48_ram[3474] = 167;
    exp_48_ram[3475] = 133;
    exp_48_ram[3476] = 240;
    exp_48_ram[3477] = 7;
    exp_48_ram[3478] = 133;
    exp_48_ram[3479] = 32;
    exp_48_ram[3480] = 36;
    exp_48_ram[3481] = 1;
    exp_48_ram[3482] = 128;
    exp_48_ram[3483] = 1;
    exp_48_ram[3484] = 38;
    exp_48_ram[3485] = 36;
    exp_48_ram[3486] = 34;
    exp_48_ram[3487] = 32;
    exp_48_ram[3488] = 4;
    exp_48_ram[3489] = 46;
    exp_48_ram[3490] = 224;
    exp_48_ram[3491] = 36;
    exp_48_ram[3492] = 38;
    exp_48_ram[3493] = 0;
    exp_48_ram[3494] = 224;
    exp_48_ram[3495] = 6;
    exp_48_ram[3496] = 134;
    exp_48_ram[3497] = 37;
    exp_48_ram[3498] = 37;
    exp_48_ram[3499] = 7;
    exp_48_ram[3500] = 8;
    exp_48_ram[3501] = 56;
    exp_48_ram[3502] = 135;
    exp_48_ram[3503] = 134;
    exp_48_ram[3504] = 135;
    exp_48_ram[3505] = 38;
    exp_48_ram[3506] = 137;
    exp_48_ram[3507] = 9;
    exp_48_ram[3508] = 134;
    exp_48_ram[3509] = 134;
    exp_48_ram[3510] = 224;
    exp_48_ram[3511] = 134;
    exp_48_ram[3512] = 134;
    exp_48_ram[3513] = 24;
    exp_48_ram[3514] = 6;
    exp_48_ram[3515] = 7;
    exp_48_ram[3516] = 228;
    exp_48_ram[3517] = 0;
    exp_48_ram[3518] = 133;
    exp_48_ram[3519] = 32;
    exp_48_ram[3520] = 36;
    exp_48_ram[3521] = 41;
    exp_48_ram[3522] = 41;
    exp_48_ram[3523] = 1;
    exp_48_ram[3524] = 128;
    exp_48_ram[3525] = 1;
    exp_48_ram[3526] = 38;
    exp_48_ram[3527] = 36;
    exp_48_ram[3528] = 4;
    exp_48_ram[3529] = 23;
    exp_48_ram[3530] = 133;
    exp_48_ram[3531] = 224;
    exp_48_ram[3532] = 0;
    exp_48_ram[3533] = 32;
    exp_48_ram[3534] = 36;
    exp_48_ram[3535] = 1;
    exp_48_ram[3536] = 128;
    exp_48_ram[3537] = 1;
    exp_48_ram[3538] = 46;
    exp_48_ram[3539] = 44;
    exp_48_ram[3540] = 4;
    exp_48_ram[3541] = 23;
    exp_48_ram[3542] = 133;
    exp_48_ram[3543] = 224;
    exp_48_ram[3544] = 7;
    exp_48_ram[3545] = 38;
    exp_48_ram[3546] = 36;
    exp_48_ram[3547] = 0;
    exp_48_ram[3548] = 37;
    exp_48_ram[3549] = 23;
    exp_48_ram[3550] = 133;
    exp_48_ram[3551] = 224;
    exp_48_ram[3552] = 0;
    exp_48_ram[3553] = 39;
    exp_48_ram[3554] = 151;
    exp_48_ram[3555] = 38;
    exp_48_ram[3556] = 71;
    exp_48_ram[3557] = 167;
    exp_48_ram[3558] = 133;
    exp_48_ram[3559] = 37;
    exp_48_ram[3560] = 208;
    exp_48_ram[3561] = 71;
    exp_48_ram[3562] = 167;
    exp_48_ram[3563] = 7;
    exp_48_ram[3564] = 87;
    exp_48_ram[3565] = 133;
    exp_48_ram[3566] = 240;
    exp_48_ram[3567] = 39;
    exp_48_ram[3568] = 7;
    exp_48_ram[3569] = 208;
    exp_48_ram[3570] = 0;
    exp_48_ram[3571] = 39;
    exp_48_ram[3572] = 215;
    exp_48_ram[3573] = 38;
    exp_48_ram[3574] = 71;
    exp_48_ram[3575] = 167;
    exp_48_ram[3576] = 133;
    exp_48_ram[3577] = 37;
    exp_48_ram[3578] = 208;
    exp_48_ram[3579] = 71;
    exp_48_ram[3580] = 167;
    exp_48_ram[3581] = 7;
    exp_48_ram[3582] = 87;
    exp_48_ram[3583] = 133;
    exp_48_ram[3584] = 240;
    exp_48_ram[3585] = 39;
    exp_48_ram[3586] = 7;
    exp_48_ram[3587] = 192;
    exp_48_ram[3588] = 39;
    exp_48_ram[3589] = 135;
    exp_48_ram[3590] = 36;
    exp_48_ram[3591] = 39;
    exp_48_ram[3592] = 7;
    exp_48_ram[3593] = 214;
    exp_48_ram[3594] = 71;
    exp_48_ram[3595] = 167;
    exp_48_ram[3596] = 133;
    exp_48_ram[3597] = 5;
    exp_48_ram[3598] = 208;
    exp_48_ram[3599] = 0;
    exp_48_ram[3600] = 32;
    exp_48_ram[3601] = 36;
    exp_48_ram[3602] = 1;
    exp_48_ram[3603] = 128;
    exp_48_ram[3604] = 1;
    exp_48_ram[3605] = 38;
    exp_48_ram[3606] = 36;
    exp_48_ram[3607] = 34;
    exp_48_ram[3608] = 32;
    exp_48_ram[3609] = 46;
    exp_48_ram[3610] = 44;
    exp_48_ram[3611] = 42;
    exp_48_ram[3612] = 40;
    exp_48_ram[3613] = 38;
    exp_48_ram[3614] = 36;
    exp_48_ram[3615] = 34;
    exp_48_ram[3616] = 32;
    exp_48_ram[3617] = 4;
    exp_48_ram[3618] = 7;
    exp_48_ram[3619] = 46;
    exp_48_ram[3620] = 7;
    exp_48_ram[3621] = 7;
    exp_48_ram[3622] = 40;
    exp_48_ram[3623] = 42;
    exp_48_ram[3624] = 224;
    exp_48_ram[3625] = 32;
    exp_48_ram[3626] = 34;
    exp_48_ram[3627] = 38;
    exp_48_ram[3628] = 0;
    exp_48_ram[3629] = 39;
    exp_48_ram[3630] = 87;
    exp_48_ram[3631] = 135;
    exp_48_ram[3632] = 7;
    exp_48_ram[3633] = 46;
    exp_48_ram[3634] = 39;
    exp_48_ram[3635] = 87;
    exp_48_ram[3636] = 135;
    exp_48_ram[3637] = 7;
    exp_48_ram[3638] = 46;
    exp_48_ram[3639] = 39;
    exp_48_ram[3640] = 87;
    exp_48_ram[3641] = 135;
    exp_48_ram[3642] = 7;
    exp_48_ram[3643] = 46;
    exp_48_ram[3644] = 39;
    exp_48_ram[3645] = 87;
    exp_48_ram[3646] = 135;
    exp_48_ram[3647] = 7;
    exp_48_ram[3648] = 46;
    exp_48_ram[3649] = 39;
    exp_48_ram[3650] = 135;
    exp_48_ram[3651] = 38;
    exp_48_ram[3652] = 224;
    exp_48_ram[3653] = 6;
    exp_48_ram[3654] = 134;
    exp_48_ram[3655] = 37;
    exp_48_ram[3656] = 37;
    exp_48_ram[3657] = 7;
    exp_48_ram[3658] = 8;
    exp_48_ram[3659] = 56;
    exp_48_ram[3660] = 135;
    exp_48_ram[3661] = 134;
    exp_48_ram[3662] = 135;
    exp_48_ram[3663] = 70;
    exp_48_ram[3664] = 166;
    exp_48_ram[3665] = 36;
    exp_48_ram[3666] = 38;
    exp_48_ram[3667] = 37;
    exp_48_ram[3668] = 37;
    exp_48_ram[3669] = 134;
    exp_48_ram[3670] = 134;
    exp_48_ram[3671] = 236;
    exp_48_ram[3672] = 134;
    exp_48_ram[3673] = 134;
    exp_48_ram[3674] = 24;
    exp_48_ram[3675] = 6;
    exp_48_ram[3676] = 7;
    exp_48_ram[3677] = 224;
    exp_48_ram[3678] = 37;
    exp_48_ram[3679] = 23;
    exp_48_ram[3680] = 133;
    exp_48_ram[3681] = 224;
    exp_48_ram[3682] = 224;
    exp_48_ram[3683] = 32;
    exp_48_ram[3684] = 34;
    exp_48_ram[3685] = 38;
    exp_48_ram[3686] = 0;
    exp_48_ram[3687] = 39;
    exp_48_ram[3688] = 39;
    exp_48_ram[3689] = 86;
    exp_48_ram[3690] = 134;
    exp_48_ram[3691] = 134;
    exp_48_ram[3692] = 6;
    exp_48_ram[3693] = 6;
    exp_48_ram[3694] = 6;
    exp_48_ram[3695] = 86;
    exp_48_ram[3696] = 134;
    exp_48_ram[3697] = 5;
    exp_48_ram[3698] = 57;
    exp_48_ram[3699] = 137;
    exp_48_ram[3700] = 7;
    exp_48_ram[3701] = 137;
    exp_48_ram[3702] = 40;
    exp_48_ram[3703] = 42;
    exp_48_ram[3704] = 39;
    exp_48_ram[3705] = 39;
    exp_48_ram[3706] = 86;
    exp_48_ram[3707] = 134;
    exp_48_ram[3708] = 134;
    exp_48_ram[3709] = 6;
    exp_48_ram[3710] = 6;
    exp_48_ram[3711] = 6;
    exp_48_ram[3712] = 86;
    exp_48_ram[3713] = 134;
    exp_48_ram[3714] = 5;
    exp_48_ram[3715] = 58;
    exp_48_ram[3716] = 138;
    exp_48_ram[3717] = 7;
    exp_48_ram[3718] = 138;
    exp_48_ram[3719] = 40;
    exp_48_ram[3720] = 42;
    exp_48_ram[3721] = 39;
    exp_48_ram[3722] = 39;
    exp_48_ram[3723] = 86;
    exp_48_ram[3724] = 134;
    exp_48_ram[3725] = 134;
    exp_48_ram[3726] = 6;
    exp_48_ram[3727] = 6;
    exp_48_ram[3728] = 6;
    exp_48_ram[3729] = 86;
    exp_48_ram[3730] = 134;
    exp_48_ram[3731] = 5;
    exp_48_ram[3732] = 59;
    exp_48_ram[3733] = 139;
    exp_48_ram[3734] = 7;
    exp_48_ram[3735] = 139;
    exp_48_ram[3736] = 40;
    exp_48_ram[3737] = 42;
    exp_48_ram[3738] = 39;
    exp_48_ram[3739] = 39;
    exp_48_ram[3740] = 86;
    exp_48_ram[3741] = 134;
    exp_48_ram[3742] = 134;
    exp_48_ram[3743] = 6;
    exp_48_ram[3744] = 6;
    exp_48_ram[3745] = 6;
    exp_48_ram[3746] = 86;
    exp_48_ram[3747] = 134;
    exp_48_ram[3748] = 5;
    exp_48_ram[3749] = 60;
    exp_48_ram[3750] = 140;
    exp_48_ram[3751] = 7;
    exp_48_ram[3752] = 140;
    exp_48_ram[3753] = 40;
    exp_48_ram[3754] = 42;
    exp_48_ram[3755] = 39;
    exp_48_ram[3756] = 135;
    exp_48_ram[3757] = 38;
    exp_48_ram[3758] = 224;
    exp_48_ram[3759] = 6;
    exp_48_ram[3760] = 134;
    exp_48_ram[3761] = 37;
    exp_48_ram[3762] = 37;
    exp_48_ram[3763] = 7;
    exp_48_ram[3764] = 8;
    exp_48_ram[3765] = 56;
    exp_48_ram[3766] = 135;
    exp_48_ram[3767] = 134;
    exp_48_ram[3768] = 135;
    exp_48_ram[3769] = 70;
    exp_48_ram[3770] = 166;
    exp_48_ram[3771] = 32;
    exp_48_ram[3772] = 34;
    exp_48_ram[3773] = 37;
    exp_48_ram[3774] = 37;
    exp_48_ram[3775] = 134;
    exp_48_ram[3776] = 134;
    exp_48_ram[3777] = 236;
    exp_48_ram[3778] = 134;
    exp_48_ram[3779] = 134;
    exp_48_ram[3780] = 24;
    exp_48_ram[3781] = 6;
    exp_48_ram[3782] = 7;
    exp_48_ram[3783] = 224;
    exp_48_ram[3784] = 37;
    exp_48_ram[3785] = 23;
    exp_48_ram[3786] = 133;
    exp_48_ram[3787] = 224;
    exp_48_ram[3788] = 224;
    exp_48_ram[3789] = 32;
    exp_48_ram[3790] = 34;
    exp_48_ram[3791] = 38;
    exp_48_ram[3792] = 0;
    exp_48_ram[3793] = 39;
    exp_48_ram[3794] = 87;
    exp_48_ram[3795] = 135;
    exp_48_ram[3796] = 87;
    exp_48_ram[3797] = 46;
    exp_48_ram[3798] = 39;
    exp_48_ram[3799] = 87;
    exp_48_ram[3800] = 135;
    exp_48_ram[3801] = 87;
    exp_48_ram[3802] = 46;
    exp_48_ram[3803] = 39;
    exp_48_ram[3804] = 87;
    exp_48_ram[3805] = 135;
    exp_48_ram[3806] = 87;
    exp_48_ram[3807] = 46;
    exp_48_ram[3808] = 39;
    exp_48_ram[3809] = 87;
    exp_48_ram[3810] = 135;
    exp_48_ram[3811] = 87;
    exp_48_ram[3812] = 46;
    exp_48_ram[3813] = 39;
    exp_48_ram[3814] = 135;
    exp_48_ram[3815] = 38;
    exp_48_ram[3816] = 224;
    exp_48_ram[3817] = 6;
    exp_48_ram[3818] = 134;
    exp_48_ram[3819] = 37;
    exp_48_ram[3820] = 37;
    exp_48_ram[3821] = 7;
    exp_48_ram[3822] = 8;
    exp_48_ram[3823] = 56;
    exp_48_ram[3824] = 135;
    exp_48_ram[3825] = 134;
    exp_48_ram[3826] = 135;
    exp_48_ram[3827] = 70;
    exp_48_ram[3828] = 166;
    exp_48_ram[3829] = 44;
    exp_48_ram[3830] = 46;
    exp_48_ram[3831] = 37;
    exp_48_ram[3832] = 37;
    exp_48_ram[3833] = 134;
    exp_48_ram[3834] = 134;
    exp_48_ram[3835] = 236;
    exp_48_ram[3836] = 134;
    exp_48_ram[3837] = 134;
    exp_48_ram[3838] = 24;
    exp_48_ram[3839] = 6;
    exp_48_ram[3840] = 7;
    exp_48_ram[3841] = 224;
    exp_48_ram[3842] = 37;
    exp_48_ram[3843] = 23;
    exp_48_ram[3844] = 133;
    exp_48_ram[3845] = 224;
    exp_48_ram[3846] = 224;
    exp_48_ram[3847] = 32;
    exp_48_ram[3848] = 34;
    exp_48_ram[3849] = 38;
    exp_48_ram[3850] = 0;
    exp_48_ram[3851] = 39;
    exp_48_ram[3852] = 39;
    exp_48_ram[3853] = 86;
    exp_48_ram[3854] = 6;
    exp_48_ram[3855] = 6;
    exp_48_ram[3856] = 5;
    exp_48_ram[3857] = 133;
    exp_48_ram[3858] = 192;
    exp_48_ram[3859] = 7;
    exp_48_ram[3860] = 135;
    exp_48_ram[3861] = 40;
    exp_48_ram[3862] = 42;
    exp_48_ram[3863] = 39;
    exp_48_ram[3864] = 39;
    exp_48_ram[3865] = 86;
    exp_48_ram[3866] = 6;
    exp_48_ram[3867] = 6;
    exp_48_ram[3868] = 5;
    exp_48_ram[3869] = 133;
    exp_48_ram[3870] = 192;
    exp_48_ram[3871] = 7;
    exp_48_ram[3872] = 135;
    exp_48_ram[3873] = 40;
    exp_48_ram[3874] = 42;
    exp_48_ram[3875] = 39;
    exp_48_ram[3876] = 39;
    exp_48_ram[3877] = 86;
    exp_48_ram[3878] = 6;
    exp_48_ram[3879] = 6;
    exp_48_ram[3880] = 5;
    exp_48_ram[3881] = 133;
    exp_48_ram[3882] = 192;
    exp_48_ram[3883] = 7;
    exp_48_ram[3884] = 135;
    exp_48_ram[3885] = 40;
    exp_48_ram[3886] = 42;
    exp_48_ram[3887] = 39;
    exp_48_ram[3888] = 39;
    exp_48_ram[3889] = 86;
    exp_48_ram[3890] = 6;
    exp_48_ram[3891] = 6;
    exp_48_ram[3892] = 5;
    exp_48_ram[3893] = 133;
    exp_48_ram[3894] = 192;
    exp_48_ram[3895] = 7;
    exp_48_ram[3896] = 135;
    exp_48_ram[3897] = 40;
    exp_48_ram[3898] = 42;
    exp_48_ram[3899] = 39;
    exp_48_ram[3900] = 135;
    exp_48_ram[3901] = 38;
    exp_48_ram[3902] = 224;
    exp_48_ram[3903] = 6;
    exp_48_ram[3904] = 134;
    exp_48_ram[3905] = 37;
    exp_48_ram[3906] = 37;
    exp_48_ram[3907] = 7;
    exp_48_ram[3908] = 8;
    exp_48_ram[3909] = 56;
    exp_48_ram[3910] = 135;
    exp_48_ram[3911] = 134;
    exp_48_ram[3912] = 135;
    exp_48_ram[3913] = 70;
    exp_48_ram[3914] = 166;
    exp_48_ram[3915] = 141;
    exp_48_ram[3916] = 13;
    exp_48_ram[3917] = 134;
    exp_48_ram[3918] = 134;
    exp_48_ram[3919] = 232;
    exp_48_ram[3920] = 134;
    exp_48_ram[3921] = 134;
    exp_48_ram[3922] = 24;
    exp_48_ram[3923] = 6;
    exp_48_ram[3924] = 7;
    exp_48_ram[3925] = 236;
    exp_48_ram[3926] = 37;
    exp_48_ram[3927] = 23;
    exp_48_ram[3928] = 133;
    exp_48_ram[3929] = 224;
    exp_48_ram[3930] = 0;
    exp_48_ram[3931] = 32;
    exp_48_ram[3932] = 36;
    exp_48_ram[3933] = 41;
    exp_48_ram[3934] = 41;
    exp_48_ram[3935] = 42;
    exp_48_ram[3936] = 42;
    exp_48_ram[3937] = 43;
    exp_48_ram[3938] = 43;
    exp_48_ram[3939] = 44;
    exp_48_ram[3940] = 44;
    exp_48_ram[3941] = 45;
    exp_48_ram[3942] = 45;
    exp_48_ram[3943] = 1;
    exp_48_ram[3944] = 128;
    exp_48_ram[3945] = 1;
    exp_48_ram[3946] = 46;
    exp_48_ram[3947] = 44;
    exp_48_ram[3948] = 42;
    exp_48_ram[3949] = 40;
    exp_48_ram[3950] = 38;
    exp_48_ram[3951] = 36;
    exp_48_ram[3952] = 4;
    exp_48_ram[3953] = 23;
    exp_48_ram[3954] = 133;
    exp_48_ram[3955] = 224;
    exp_48_ram[3956] = 240;
    exp_48_ram[3957] = 7;
    exp_48_ram[3958] = 135;
    exp_48_ram[3959] = 34;
    exp_48_ram[3960] = 23;
    exp_48_ram[3961] = 133;
    exp_48_ram[3962] = 224;
    exp_48_ram[3963] = 240;
    exp_48_ram[3964] = 7;
    exp_48_ram[3965] = 135;
    exp_48_ram[3966] = 32;
    exp_48_ram[3967] = 23;
    exp_48_ram[3968] = 133;
    exp_48_ram[3969] = 224;
    exp_48_ram[3970] = 240;
    exp_48_ram[3971] = 7;
    exp_48_ram[3972] = 46;
    exp_48_ram[3973] = 23;
    exp_48_ram[3974] = 133;
    exp_48_ram[3975] = 224;
    exp_48_ram[3976] = 240;
    exp_48_ram[3977] = 7;
    exp_48_ram[3978] = 44;
    exp_48_ram[3979] = 23;
    exp_48_ram[3980] = 133;
    exp_48_ram[3981] = 224;
    exp_48_ram[3982] = 240;
    exp_48_ram[3983] = 7;
    exp_48_ram[3984] = 42;
    exp_48_ram[3985] = 7;
    exp_48_ram[3986] = 40;
    exp_48_ram[3987] = 7;
    exp_48_ram[3988] = 40;
    exp_48_ram[3989] = 7;
    exp_48_ram[3990] = 133;
    exp_48_ram[3991] = 224;
    exp_48_ram[3992] = 7;
    exp_48_ram[3993] = 135;
    exp_48_ram[3994] = 36;
    exp_48_ram[3995] = 38;
    exp_48_ram[3996] = 39;
    exp_48_ram[3997] = 39;
    exp_48_ram[3998] = 5;
    exp_48_ram[3999] = 133;
    exp_48_ram[4000] = 224;
    exp_48_ram[4001] = 224;
    exp_48_ram[4002] = 44;
    exp_48_ram[4003] = 46;
    exp_48_ram[4004] = 42;
    exp_48_ram[4005] = 0;
    exp_48_ram[4006] = 0;
    exp_48_ram[4007] = 224;
    exp_48_ram[4008] = 7;
    exp_48_ram[4009] = 135;
    exp_48_ram[4010] = 38;
    exp_48_ram[4011] = 38;
    exp_48_ram[4012] = 5;
    exp_48_ram[4013] = 133;
    exp_48_ram[4014] = 224;
    exp_48_ram[4015] = 10;
    exp_48_ram[4016] = 138;
    exp_48_ram[4017] = 71;
    exp_48_ram[4018] = 167;
    exp_48_ram[4019] = 133;
    exp_48_ram[4020] = 192;
    exp_48_ram[4021] = 7;
    exp_48_ram[4022] = 135;
    exp_48_ram[4023] = 6;
    exp_48_ram[4024] = 134;
    exp_48_ram[4025] = 5;
    exp_48_ram[4026] = 133;
    exp_48_ram[4027] = 192;
    exp_48_ram[4028] = 7;
    exp_48_ram[4029] = 196;
    exp_48_ram[4030] = 71;
    exp_48_ram[4031] = 167;
    exp_48_ram[4032] = 137;
    exp_48_ram[4033] = 9;
    exp_48_ram[4034] = 38;
    exp_48_ram[4035] = 38;
    exp_48_ram[4036] = 7;
    exp_48_ram[4037] = 5;
    exp_48_ram[4038] = 181;
    exp_48_ram[4039] = 135;
    exp_48_ram[4040] = 134;
    exp_48_ram[4041] = 135;
    exp_48_ram[4042] = 44;
    exp_48_ram[4043] = 46;
    exp_48_ram[4044] = 5;
    exp_48_ram[4045] = 224;
    exp_48_ram[4046] = 7;
    exp_48_ram[4047] = 135;
    exp_48_ram[4048] = 36;
    exp_48_ram[4049] = 38;
    exp_48_ram[4050] = 7;
    exp_48_ram[4051] = 133;
    exp_48_ram[4052] = 240;
    exp_48_ram[4053] = 7;
    exp_48_ram[4054] = 133;
    exp_48_ram[4055] = 192;
    exp_48_ram[4056] = 39;
    exp_48_ram[4057] = 135;
    exp_48_ram[4058] = 42;
    exp_48_ram[4059] = 39;
    exp_48_ram[4060] = 7;
    exp_48_ram[4061] = 210;
    exp_48_ram[4062] = 0;
    exp_48_ram[4063] = 0;
    exp_48_ram[4064] = 32;
    exp_48_ram[4065] = 36;
    exp_48_ram[4066] = 41;
    exp_48_ram[4067] = 41;
    exp_48_ram[4068] = 42;
    exp_48_ram[4069] = 42;
    exp_48_ram[4070] = 1;
    exp_48_ram[4071] = 128;
    exp_48_ram[4072] = 1;
    exp_48_ram[4073] = 46;
    exp_48_ram[4074] = 44;
    exp_48_ram[4075] = 4;
    exp_48_ram[4076] = 23;
    exp_48_ram[4077] = 133;
    exp_48_ram[4078] = 208;
    exp_48_ram[4079] = 23;
    exp_48_ram[4080] = 133;
    exp_48_ram[4081] = 208;
    exp_48_ram[4082] = 23;
    exp_48_ram[4083] = 133;
    exp_48_ram[4084] = 208;
    exp_48_ram[4085] = 23;
    exp_48_ram[4086] = 133;
    exp_48_ram[4087] = 208;
    exp_48_ram[4088] = 23;
    exp_48_ram[4089] = 133;
    exp_48_ram[4090] = 208;
    exp_48_ram[4091] = 192;
    exp_48_ram[4092] = 7;
    exp_48_ram[4093] = 7;
    exp_48_ram[4094] = 71;
    exp_48_ram[4095] = 7;
    exp_48_ram[4096] = 132;
    exp_48_ram[4097] = 7;
    exp_48_ram[4098] = 68;
    exp_48_ram[4099] = 7;
    exp_48_ram[4100] = 136;
    exp_48_ram[4101] = 7;
    exp_48_ram[4102] = 76;
    exp_48_ram[4103] = 7;
    exp_48_ram[4104] = 136;
    exp_48_ram[4105] = 7;
    exp_48_ram[4106] = 136;
    exp_48_ram[4107] = 0;
    exp_48_ram[4108] = 240;
    exp_48_ram[4109] = 0;
    exp_48_ram[4110] = 240;
    exp_48_ram[4111] = 0;
    exp_48_ram[4112] = 240;
    exp_48_ram[4113] = 0;
    exp_48_ram[4114] = 240;
    exp_48_ram[4115] = 0;
    exp_48_ram[4116] = 240;
    exp_48_ram[4117] = 7;
    exp_48_ram[4118] = 135;
    exp_48_ram[4119] = 69;
    exp_48_ram[4120] = 1;
    exp_48_ram[4121] = 101;
    exp_48_ram[4122] = 76;
    exp_48_ram[4123] = 214;
    exp_48_ram[4124] = 5;
    exp_48_ram[4125] = 133;
    exp_48_ram[4126] = 1;
    exp_48_ram[4127] = 128;
    exp_48_ram[4128] = 92;
    exp_48_ram[4129] = 5;
    exp_48_ram[4130] = 133;
    exp_48_ram[4131] = 240;
    exp_48_ram[4132] = 240;
    exp_48_ram[4133] = 0;
    exp_48_ram[4134] = 0;
    exp_48_ram[4135] = 0;
    exp_48_ram[4136] = 21;
    exp_48_ram[4137] = 21;
    exp_48_ram[4138] = 21;
    exp_48_ram[4139] = 21;
    exp_48_ram[4140] = 21;
    exp_48_ram[4141] = 21;
    exp_48_ram[4142] = 21;
    exp_48_ram[4143] = 21;
    exp_48_ram[4144] = 21;
    exp_48_ram[4145] = 21;
    exp_48_ram[4146] = 21;
    exp_48_ram[4147] = 21;
    exp_48_ram[4148] = 21;
    exp_48_ram[4149] = 20;
    exp_48_ram[4150] = 21;
    exp_48_ram[4151] = 21;
    exp_48_ram[4152] = 20;
    exp_48_ram[4153] = 23;
    exp_48_ram[4154] = 23;
    exp_48_ram[4155] = 23;
    exp_48_ram[4156] = 23;
    exp_48_ram[4157] = 22;
    exp_48_ram[4158] = 23;
    exp_48_ram[4159] = 23;
    exp_48_ram[4160] = 23;
    exp_48_ram[4161] = 23;
    exp_48_ram[4162] = 23;
    exp_48_ram[4163] = 23;
    exp_48_ram[4164] = 23;
    exp_48_ram[4165] = 23;
    exp_48_ram[4166] = 23;
    exp_48_ram[4167] = 23;
    exp_48_ram[4168] = 23;
    exp_48_ram[4169] = 23;
    exp_48_ram[4170] = 23;
    exp_48_ram[4171] = 23;
    exp_48_ram[4172] = 29;
    exp_48_ram[4173] = 30;
    exp_48_ram[4174] = 30;
    exp_48_ram[4175] = 30;
    exp_48_ram[4176] = 30;
    exp_48_ram[4177] = 30;
    exp_48_ram[4178] = 30;
    exp_48_ram[4179] = 30;
    exp_48_ram[4180] = 30;
    exp_48_ram[4181] = 30;
    exp_48_ram[4182] = 30;
    exp_48_ram[4183] = 30;
    exp_48_ram[4184] = 30;
    exp_48_ram[4185] = 30;
    exp_48_ram[4186] = 30;
    exp_48_ram[4187] = 30;
    exp_48_ram[4188] = 30;
    exp_48_ram[4189] = 30;
    exp_48_ram[4190] = 30;
    exp_48_ram[4191] = 30;
    exp_48_ram[4192] = 30;
    exp_48_ram[4193] = 30;
    exp_48_ram[4194] = 30;
    exp_48_ram[4195] = 30;
    exp_48_ram[4196] = 30;
    exp_48_ram[4197] = 30;
    exp_48_ram[4198] = 30;
    exp_48_ram[4199] = 30;
    exp_48_ram[4200] = 30;
    exp_48_ram[4201] = 30;
    exp_48_ram[4202] = 30;
    exp_48_ram[4203] = 30;
    exp_48_ram[4204] = 30;
    exp_48_ram[4205] = 30;
    exp_48_ram[4206] = 30;
    exp_48_ram[4207] = 30;
    exp_48_ram[4208] = 30;
    exp_48_ram[4209] = 30;
    exp_48_ram[4210] = 30;
    exp_48_ram[4211] = 30;
    exp_48_ram[4212] = 30;
    exp_48_ram[4213] = 30;
    exp_48_ram[4214] = 30;
    exp_48_ram[4215] = 30;
    exp_48_ram[4216] = 30;
    exp_48_ram[4217] = 30;
    exp_48_ram[4218] = 30;
    exp_48_ram[4219] = 30;
    exp_48_ram[4220] = 30;
    exp_48_ram[4221] = 30;
    exp_48_ram[4222] = 30;
    exp_48_ram[4223] = 23;
    exp_48_ram[4224] = 30;
    exp_48_ram[4225] = 30;
    exp_48_ram[4226] = 30;
    exp_48_ram[4227] = 30;
    exp_48_ram[4228] = 30;
    exp_48_ram[4229] = 30;
    exp_48_ram[4230] = 30;
    exp_48_ram[4231] = 30;
    exp_48_ram[4232] = 30;
    exp_48_ram[4233] = 23;
    exp_48_ram[4234] = 27;
    exp_48_ram[4235] = 23;
    exp_48_ram[4236] = 30;
    exp_48_ram[4237] = 30;
    exp_48_ram[4238] = 30;
    exp_48_ram[4239] = 30;
    exp_48_ram[4240] = 23;
    exp_48_ram[4241] = 30;
    exp_48_ram[4242] = 30;
    exp_48_ram[4243] = 30;
    exp_48_ram[4244] = 30;
    exp_48_ram[4245] = 30;
    exp_48_ram[4246] = 23;
    exp_48_ram[4247] = 29;
    exp_48_ram[4248] = 30;
    exp_48_ram[4249] = 30;
    exp_48_ram[4250] = 28;
    exp_48_ram[4251] = 30;
    exp_48_ram[4252] = 23;
    exp_48_ram[4253] = 30;
    exp_48_ram[4254] = 30;
    exp_48_ram[4255] = 23;
    exp_48_ram[4256] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_46) begin
      exp_48_ram[exp_42] <= exp_44;
    end
  end
  assign exp_48 = exp_48_ram[exp_43];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_74) begin
        exp_48_ram[exp_70] <= exp_72;
    end
  end
  assign exp_76 = exp_48_ram[exp_71];
  assign exp_75 = exp_98;
  assign exp_98 = 1;
  assign exp_71 = exp_97;
  assign exp_97 = exp_16[31:2];
  assign exp_74 = exp_92;
  assign exp_70 = exp_91;
  assign exp_72 = exp_91;
  assign exp_47 = exp_133;
  assign exp_133 = 1;
  assign exp_43 = exp_132;
  assign exp_132 = exp_18[31:2];
  assign exp_46 = exp_114;
  assign exp_114 = exp_112 & exp_113;
  assign exp_112 = exp_22 & exp_23;
  assign exp_113 = exp_24[1:1];
  assign exp_42 = exp_110;
  assign exp_110 = exp_18[31:2];
  assign exp_44 = exp_111;
  assign exp_111 = exp_19[15:8];

  //Create RAM
  reg [7:0] exp_41_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_41_ram[0] = 147;
    exp_41_ram[1] = 19;
    exp_41_ram[2] = 147;
    exp_41_ram[3] = 19;
    exp_41_ram[4] = 147;
    exp_41_ram[5] = 19;
    exp_41_ram[6] = 147;
    exp_41_ram[7] = 19;
    exp_41_ram[8] = 147;
    exp_41_ram[9] = 19;
    exp_41_ram[10] = 147;
    exp_41_ram[11] = 19;
    exp_41_ram[12] = 147;
    exp_41_ram[13] = 19;
    exp_41_ram[14] = 147;
    exp_41_ram[15] = 19;
    exp_41_ram[16] = 147;
    exp_41_ram[17] = 19;
    exp_41_ram[18] = 147;
    exp_41_ram[19] = 19;
    exp_41_ram[20] = 147;
    exp_41_ram[21] = 19;
    exp_41_ram[22] = 147;
    exp_41_ram[23] = 19;
    exp_41_ram[24] = 147;
    exp_41_ram[25] = 19;
    exp_41_ram[26] = 147;
    exp_41_ram[27] = 19;
    exp_41_ram[28] = 147;
    exp_41_ram[29] = 19;
    exp_41_ram[30] = 147;
    exp_41_ram[31] = 55;
    exp_41_ram[32] = 19;
    exp_41_ram[33] = 239;
    exp_41_ram[34] = 111;
    exp_41_ram[35] = 147;
    exp_41_ram[36] = 147;
    exp_41_ram[37] = 19;
    exp_41_ram[38] = 19;
    exp_41_ram[39] = 19;
    exp_41_ram[40] = 99;
    exp_41_ram[41] = 183;
    exp_41_ram[42] = 147;
    exp_41_ram[43] = 99;
    exp_41_ram[44] = 55;
    exp_41_ram[45] = 99;
    exp_41_ram[46] = 19;
    exp_41_ram[47] = 51;
    exp_41_ram[48] = 19;
    exp_41_ram[49] = 51;
    exp_41_ram[50] = 179;
    exp_41_ram[51] = 131;
    exp_41_ram[52] = 19;
    exp_41_ram[53] = 51;
    exp_41_ram[54] = 179;
    exp_41_ram[55] = 99;
    exp_41_ram[56] = 179;
    exp_41_ram[57] = 51;
    exp_41_ram[58] = 51;
    exp_41_ram[59] = 179;
    exp_41_ram[60] = 51;
    exp_41_ram[61] = 147;
    exp_41_ram[62] = 179;
    exp_41_ram[63] = 19;
    exp_41_ram[64] = 19;
    exp_41_ram[65] = 147;
    exp_41_ram[66] = 51;
    exp_41_ram[67] = 19;
    exp_41_ram[68] = 179;
    exp_41_ram[69] = 19;
    exp_41_ram[70] = 179;
    exp_41_ram[71] = 99;
    exp_41_ram[72] = 179;
    exp_41_ram[73] = 19;
    exp_41_ram[74] = 99;
    exp_41_ram[75] = 99;
    exp_41_ram[76] = 19;
    exp_41_ram[77] = 179;
    exp_41_ram[78] = 179;
    exp_41_ram[79] = 51;
    exp_41_ram[80] = 19;
    exp_41_ram[81] = 19;
    exp_41_ram[82] = 179;
    exp_41_ram[83] = 19;
    exp_41_ram[84] = 51;
    exp_41_ram[85] = 179;
    exp_41_ram[86] = 19;
    exp_41_ram[87] = 99;
    exp_41_ram[88] = 51;
    exp_41_ram[89] = 19;
    exp_41_ram[90] = 99;
    exp_41_ram[91] = 99;
    exp_41_ram[92] = 19;
    exp_41_ram[93] = 19;
    exp_41_ram[94] = 51;
    exp_41_ram[95] = 147;
    exp_41_ram[96] = 111;
    exp_41_ram[97] = 55;
    exp_41_ram[98] = 19;
    exp_41_ram[99] = 227;
    exp_41_ram[100] = 19;
    exp_41_ram[101] = 111;
    exp_41_ram[102] = 99;
    exp_41_ram[103] = 19;
    exp_41_ram[104] = 51;
    exp_41_ram[105] = 55;
    exp_41_ram[106] = 99;
    exp_41_ram[107] = 19;
    exp_41_ram[108] = 99;
    exp_41_ram[109] = 19;
    exp_41_ram[110] = 51;
    exp_41_ram[111] = 179;
    exp_41_ram[112] = 3;
    exp_41_ram[113] = 19;
    exp_41_ram[114] = 51;
    exp_41_ram[115] = 179;
    exp_41_ram[116] = 99;
    exp_41_ram[117] = 179;
    exp_41_ram[118] = 147;
    exp_41_ram[119] = 147;
    exp_41_ram[120] = 19;
    exp_41_ram[121] = 19;
    exp_41_ram[122] = 19;
    exp_41_ram[123] = 179;
    exp_41_ram[124] = 179;
    exp_41_ram[125] = 147;
    exp_41_ram[126] = 51;
    exp_41_ram[127] = 51;
    exp_41_ram[128] = 19;
    exp_41_ram[129] = 99;
    exp_41_ram[130] = 51;
    exp_41_ram[131] = 19;
    exp_41_ram[132] = 99;
    exp_41_ram[133] = 99;
    exp_41_ram[134] = 19;
    exp_41_ram[135] = 51;
    exp_41_ram[136] = 51;
    exp_41_ram[137] = 179;
    exp_41_ram[138] = 19;
    exp_41_ram[139] = 19;
    exp_41_ram[140] = 51;
    exp_41_ram[141] = 147;
    exp_41_ram[142] = 51;
    exp_41_ram[143] = 179;
    exp_41_ram[144] = 19;
    exp_41_ram[145] = 99;
    exp_41_ram[146] = 51;
    exp_41_ram[147] = 19;
    exp_41_ram[148] = 99;
    exp_41_ram[149] = 99;
    exp_41_ram[150] = 19;
    exp_41_ram[151] = 19;
    exp_41_ram[152] = 51;
    exp_41_ram[153] = 103;
    exp_41_ram[154] = 55;
    exp_41_ram[155] = 19;
    exp_41_ram[156] = 227;
    exp_41_ram[157] = 19;
    exp_41_ram[158] = 111;
    exp_41_ram[159] = 51;
    exp_41_ram[160] = 51;
    exp_41_ram[161] = 51;
    exp_41_ram[162] = 179;
    exp_41_ram[163] = 51;
    exp_41_ram[164] = 147;
    exp_41_ram[165] = 51;
    exp_41_ram[166] = 51;
    exp_41_ram[167] = 147;
    exp_41_ram[168] = 147;
    exp_41_ram[169] = 147;
    exp_41_ram[170] = 51;
    exp_41_ram[171] = 19;
    exp_41_ram[172] = 51;
    exp_41_ram[173] = 179;
    exp_41_ram[174] = 147;
    exp_41_ram[175] = 99;
    exp_41_ram[176] = 51;
    exp_41_ram[177] = 147;
    exp_41_ram[178] = 99;
    exp_41_ram[179] = 99;
    exp_41_ram[180] = 147;
    exp_41_ram[181] = 51;
    exp_41_ram[182] = 179;
    exp_41_ram[183] = 51;
    exp_41_ram[184] = 19;
    exp_41_ram[185] = 19;
    exp_41_ram[186] = 179;
    exp_41_ram[187] = 19;
    exp_41_ram[188] = 51;
    exp_41_ram[189] = 179;
    exp_41_ram[190] = 19;
    exp_41_ram[191] = 99;
    exp_41_ram[192] = 179;
    exp_41_ram[193] = 19;
    exp_41_ram[194] = 99;
    exp_41_ram[195] = 99;
    exp_41_ram[196] = 19;
    exp_41_ram[197] = 179;
    exp_41_ram[198] = 147;
    exp_41_ram[199] = 179;
    exp_41_ram[200] = 179;
    exp_41_ram[201] = 111;
    exp_41_ram[202] = 99;
    exp_41_ram[203] = 55;
    exp_41_ram[204] = 99;
    exp_41_ram[205] = 19;
    exp_41_ram[206] = 179;
    exp_41_ram[207] = 147;
    exp_41_ram[208] = 55;
    exp_41_ram[209] = 51;
    exp_41_ram[210] = 19;
    exp_41_ram[211] = 51;
    exp_41_ram[212] = 3;
    exp_41_ram[213] = 19;
    exp_41_ram[214] = 51;
    exp_41_ram[215] = 179;
    exp_41_ram[216] = 99;
    exp_41_ram[217] = 19;
    exp_41_ram[218] = 227;
    exp_41_ram[219] = 51;
    exp_41_ram[220] = 19;
    exp_41_ram[221] = 111;
    exp_41_ram[222] = 55;
    exp_41_ram[223] = 147;
    exp_41_ram[224] = 227;
    exp_41_ram[225] = 147;
    exp_41_ram[226] = 111;
    exp_41_ram[227] = 51;
    exp_41_ram[228] = 179;
    exp_41_ram[229] = 51;
    exp_41_ram[230] = 51;
    exp_41_ram[231] = 147;
    exp_41_ram[232] = 179;
    exp_41_ram[233] = 179;
    exp_41_ram[234] = 51;
    exp_41_ram[235] = 51;
    exp_41_ram[236] = 51;
    exp_41_ram[237] = 147;
    exp_41_ram[238] = 147;
    exp_41_ram[239] = 19;
    exp_41_ram[240] = 51;
    exp_41_ram[241] = 147;
    exp_41_ram[242] = 51;
    exp_41_ram[243] = 51;
    exp_41_ram[244] = 19;
    exp_41_ram[245] = 99;
    exp_41_ram[246] = 51;
    exp_41_ram[247] = 19;
    exp_41_ram[248] = 99;
    exp_41_ram[249] = 99;
    exp_41_ram[250] = 19;
    exp_41_ram[251] = 51;
    exp_41_ram[252] = 51;
    exp_41_ram[253] = 179;
    exp_41_ram[254] = 51;
    exp_41_ram[255] = 147;
    exp_41_ram[256] = 51;
    exp_41_ram[257] = 147;
    exp_41_ram[258] = 147;
    exp_41_ram[259] = 179;
    exp_41_ram[260] = 19;
    exp_41_ram[261] = 99;
    exp_41_ram[262] = 179;
    exp_41_ram[263] = 19;
    exp_41_ram[264] = 99;
    exp_41_ram[265] = 99;
    exp_41_ram[266] = 19;
    exp_41_ram[267] = 179;
    exp_41_ram[268] = 19;
    exp_41_ram[269] = 183;
    exp_41_ram[270] = 51;
    exp_41_ram[271] = 147;
    exp_41_ram[272] = 51;
    exp_41_ram[273] = 19;
    exp_41_ram[274] = 179;
    exp_41_ram[275] = 19;
    exp_41_ram[276] = 179;
    exp_41_ram[277] = 51;
    exp_41_ram[278] = 179;
    exp_41_ram[279] = 19;
    exp_41_ram[280] = 51;
    exp_41_ram[281] = 51;
    exp_41_ram[282] = 51;
    exp_41_ram[283] = 51;
    exp_41_ram[284] = 99;
    exp_41_ram[285] = 51;
    exp_41_ram[286] = 147;
    exp_41_ram[287] = 51;
    exp_41_ram[288] = 99;
    exp_41_ram[289] = 227;
    exp_41_ram[290] = 183;
    exp_41_ram[291] = 147;
    exp_41_ram[292] = 51;
    exp_41_ram[293] = 19;
    exp_41_ram[294] = 51;
    exp_41_ram[295] = 179;
    exp_41_ram[296] = 51;
    exp_41_ram[297] = 147;
    exp_41_ram[298] = 227;
    exp_41_ram[299] = 19;
    exp_41_ram[300] = 111;
    exp_41_ram[301] = 147;
    exp_41_ram[302] = 19;
    exp_41_ram[303] = 111;
    exp_41_ram[304] = 55;
    exp_41_ram[305] = 19;
    exp_41_ram[306] = 19;
    exp_41_ram[307] = 179;
    exp_41_ram[308] = 147;
    exp_41_ram[309] = 19;
    exp_41_ram[310] = 19;
    exp_41_ram[311] = 19;
    exp_41_ram[312] = 147;
    exp_41_ram[313] = 147;
    exp_41_ram[314] = 51;
    exp_41_ram[315] = 19;
    exp_41_ram[316] = 147;
    exp_41_ram[317] = 147;
    exp_41_ram[318] = 99;
    exp_41_ram[319] = 179;
    exp_41_ram[320] = 99;
    exp_41_ram[321] = 19;
    exp_41_ram[322] = 103;
    exp_41_ram[323] = 99;
    exp_41_ram[324] = 179;
    exp_41_ram[325] = 227;
    exp_41_ram[326] = 99;
    exp_41_ram[327] = 179;
    exp_41_ram[328] = 147;
    exp_41_ram[329] = 99;
    exp_41_ram[330] = 51;
    exp_41_ram[331] = 99;
    exp_41_ram[332] = 99;
    exp_41_ram[333] = 99;
    exp_41_ram[334] = 99;
    exp_41_ram[335] = 99;
    exp_41_ram[336] = 19;
    exp_41_ram[337] = 103;
    exp_41_ram[338] = 19;
    exp_41_ram[339] = 99;
    exp_41_ram[340] = 19;
    exp_41_ram[341] = 103;
    exp_41_ram[342] = 99;
    exp_41_ram[343] = 227;
    exp_41_ram[344] = 103;
    exp_41_ram[345] = 227;
    exp_41_ram[346] = 99;
    exp_41_ram[347] = 227;
    exp_41_ram[348] = 227;
    exp_41_ram[349] = 19;
    exp_41_ram[350] = 103;
    exp_41_ram[351] = 19;
    exp_41_ram[352] = 103;
    exp_41_ram[353] = 227;
    exp_41_ram[354] = 111;
    exp_41_ram[355] = 227;
    exp_41_ram[356] = 111;
    exp_41_ram[357] = 227;
    exp_41_ram[358] = 227;
    exp_41_ram[359] = 147;
    exp_41_ram[360] = 111;
    exp_41_ram[361] = 19;
    exp_41_ram[362] = 35;
    exp_41_ram[363] = 35;
    exp_41_ram[364] = 19;
    exp_41_ram[365] = 99;
    exp_41_ram[366] = 239;
    exp_41_ram[367] = 19;
    exp_41_ram[368] = 147;
    exp_41_ram[369] = 51;
    exp_41_ram[370] = 99;
    exp_41_ram[371] = 147;
    exp_41_ram[372] = 179;
    exp_41_ram[373] = 19;
    exp_41_ram[374] = 179;
    exp_41_ram[375] = 51;
    exp_41_ram[376] = 131;
    exp_41_ram[377] = 19;
    exp_41_ram[378] = 147;
    exp_41_ram[379] = 3;
    exp_41_ram[380] = 19;
    exp_41_ram[381] = 147;
    exp_41_ram[382] = 179;
    exp_41_ram[383] = 147;
    exp_41_ram[384] = 19;
    exp_41_ram[385] = 103;
    exp_41_ram[386] = 147;
    exp_41_ram[387] = 179;
    exp_41_ram[388] = 19;
    exp_41_ram[389] = 111;
    exp_41_ram[390] = 147;
    exp_41_ram[391] = 19;
    exp_41_ram[392] = 111;
    exp_41_ram[393] = 19;
    exp_41_ram[394] = 35;
    exp_41_ram[395] = 35;
    exp_41_ram[396] = 35;
    exp_41_ram[397] = 35;
    exp_41_ram[398] = 35;
    exp_41_ram[399] = 35;
    exp_41_ram[400] = 179;
    exp_41_ram[401] = 99;
    exp_41_ram[402] = 19;
    exp_41_ram[403] = 19;
    exp_41_ram[404] = 147;
    exp_41_ram[405] = 99;
    exp_41_ram[406] = 19;
    exp_41_ram[407] = 239;
    exp_41_ram[408] = 147;
    exp_41_ram[409] = 19;
    exp_41_ram[410] = 51;
    exp_41_ram[411] = 147;
    exp_41_ram[412] = 99;
    exp_41_ram[413] = 19;
    exp_41_ram[414] = 147;
    exp_41_ram[415] = 99;
    exp_41_ram[416] = 19;
    exp_41_ram[417] = 99;
    exp_41_ram[418] = 147;
    exp_41_ram[419] = 19;
    exp_41_ram[420] = 179;
    exp_41_ram[421] = 179;
    exp_41_ram[422] = 179;
    exp_41_ram[423] = 179;
    exp_41_ram[424] = 179;
    exp_41_ram[425] = 131;
    exp_41_ram[426] = 3;
    exp_41_ram[427] = 147;
    exp_41_ram[428] = 19;
    exp_41_ram[429] = 147;
    exp_41_ram[430] = 51;
    exp_41_ram[431] = 131;
    exp_41_ram[432] = 3;
    exp_41_ram[433] = 131;
    exp_41_ram[434] = 3;
    exp_41_ram[435] = 19;
    exp_41_ram[436] = 147;
    exp_41_ram[437] = 19;
    exp_41_ram[438] = 103;
    exp_41_ram[439] = 239;
    exp_41_ram[440] = 147;
    exp_41_ram[441] = 111;
    exp_41_ram[442] = 147;
    exp_41_ram[443] = 179;
    exp_41_ram[444] = 147;
    exp_41_ram[445] = 111;
    exp_41_ram[446] = 147;
    exp_41_ram[447] = 99;
    exp_41_ram[448] = 19;
    exp_41_ram[449] = 19;
    exp_41_ram[450] = 147;
    exp_41_ram[451] = 239;
    exp_41_ram[452] = 51;
    exp_41_ram[453] = 19;
    exp_41_ram[454] = 179;
    exp_41_ram[455] = 147;
    exp_41_ram[456] = 19;
    exp_41_ram[457] = 51;
    exp_41_ram[458] = 239;
    exp_41_ram[459] = 51;
    exp_41_ram[460] = 19;
    exp_41_ram[461] = 19;
    exp_41_ram[462] = 147;
    exp_41_ram[463] = 147;
    exp_41_ram[464] = 99;
    exp_41_ram[465] = 19;
    exp_41_ram[466] = 99;
    exp_41_ram[467] = 19;
    exp_41_ram[468] = 179;
    exp_41_ram[469] = 19;
    exp_41_ram[470] = 51;
    exp_41_ram[471] = 51;
    exp_41_ram[472] = 179;
    exp_41_ram[473] = 179;
    exp_41_ram[474] = 55;
    exp_41_ram[475] = 19;
    exp_41_ram[476] = 179;
    exp_41_ram[477] = 19;
    exp_41_ram[478] = 99;
    exp_41_ram[479] = 19;
    exp_41_ram[480] = 147;
    exp_41_ram[481] = 99;
    exp_41_ram[482] = 19;
    exp_41_ram[483] = 179;
    exp_41_ram[484] = 179;
    exp_41_ram[485] = 147;
    exp_41_ram[486] = 55;
    exp_41_ram[487] = 51;
    exp_41_ram[488] = 99;
    exp_41_ram[489] = 55;
    exp_41_ram[490] = 19;
    exp_41_ram[491] = 19;
    exp_41_ram[492] = 179;
    exp_41_ram[493] = 51;
    exp_41_ram[494] = 147;
    exp_41_ram[495] = 19;
    exp_41_ram[496] = 179;
    exp_41_ram[497] = 147;
    exp_41_ram[498] = 111;
    exp_41_ram[499] = 147;
    exp_41_ram[500] = 179;
    exp_41_ram[501] = 147;
    exp_41_ram[502] = 111;
    exp_41_ram[503] = 147;
    exp_41_ram[504] = 147;
    exp_41_ram[505] = 19;
    exp_41_ram[506] = 111;
    exp_41_ram[507] = 99;
    exp_41_ram[508] = 147;
    exp_41_ram[509] = 179;
    exp_41_ram[510] = 99;
    exp_41_ram[511] = 19;
    exp_41_ram[512] = 19;
    exp_41_ram[513] = 51;
    exp_41_ram[514] = 147;
    exp_41_ram[515] = 103;
    exp_41_ram[516] = 51;
    exp_41_ram[517] = 51;
    exp_41_ram[518] = 179;
    exp_41_ram[519] = 51;
    exp_41_ram[520] = 111;
    exp_41_ram[521] = 99;
    exp_41_ram[522] = 147;
    exp_41_ram[523] = 179;
    exp_41_ram[524] = 99;
    exp_41_ram[525] = 147;
    exp_41_ram[526] = 19;
    exp_41_ram[527] = 179;
    exp_41_ram[528] = 19;
    exp_41_ram[529] = 103;
    exp_41_ram[530] = 51;
    exp_41_ram[531] = 179;
    exp_41_ram[532] = 51;
    exp_41_ram[533] = 179;
    exp_41_ram[534] = 111;
    exp_41_ram[535] = 183;
    exp_41_ram[536] = 99;
    exp_41_ram[537] = 147;
    exp_41_ram[538] = 179;
    exp_41_ram[539] = 147;
    exp_41_ram[540] = 55;
    exp_41_ram[541] = 147;
    exp_41_ram[542] = 179;
    exp_41_ram[543] = 51;
    exp_41_ram[544] = 147;
    exp_41_ram[545] = 51;
    exp_41_ram[546] = 3;
    exp_41_ram[547] = 51;
    exp_41_ram[548] = 103;
    exp_41_ram[549] = 55;
    exp_41_ram[550] = 147;
    exp_41_ram[551] = 227;
    exp_41_ram[552] = 147;
    exp_41_ram[553] = 111;
    exp_41_ram[554] = 83;
    exp_41_ram[555] = 111;
    exp_41_ram[556] = 101;
    exp_41_ram[557] = 84;
    exp_41_ram[558] = 114;
    exp_41_ram[559] = 116;
    exp_41_ram[560] = 74;
    exp_41_ram[561] = 101;
    exp_41_ram[562] = 114;
    exp_41_ram[563] = 77;
    exp_41_ram[564] = 117;
    exp_41_ram[565] = 108;
    exp_41_ram[566] = 83;
    exp_41_ram[567] = 99;
    exp_41_ram[568] = 118;
    exp_41_ram[569] = 0;
    exp_41_ram[570] = 72;
    exp_41_ram[571] = 111;
    exp_41_ram[572] = 114;
    exp_41_ram[573] = 10;
    exp_41_ram[574] = 114;
    exp_41_ram[575] = 105;
    exp_41_ram[576] = 107;
    exp_41_ram[577] = 104;
    exp_41_ram[578] = 105;
    exp_41_ram[579] = 32;
    exp_41_ram[580] = 111;
    exp_41_ram[581] = 10;
    exp_41_ram[582] = 37;
    exp_41_ram[583] = 37;
    exp_41_ram[584] = 50;
    exp_41_ram[585] = 116;
    exp_41_ram[586] = 116;
    exp_41_ram[587] = 114;
    exp_41_ram[588] = 108;
    exp_41_ram[589] = 108;
    exp_41_ram[590] = 32;
    exp_41_ram[591] = 49;
    exp_41_ram[592] = 99;
    exp_41_ram[593] = 10;
    exp_41_ram[594] = 37;
    exp_41_ram[595] = 52;
    exp_41_ram[596] = 116;
    exp_41_ram[597] = 116;
    exp_41_ram[598] = 114;
    exp_41_ram[599] = 108;
    exp_41_ram[600] = 108;
    exp_41_ram[601] = 32;
    exp_41_ram[602] = 49;
    exp_41_ram[603] = 99;
    exp_41_ram[604] = 10;
    exp_41_ram[605] = 37;
    exp_41_ram[606] = 50;
    exp_41_ram[607] = 116;
    exp_41_ram[608] = 116;
    exp_41_ram[609] = 114;
    exp_41_ram[610] = 118;
    exp_41_ram[611] = 115;
    exp_41_ram[612] = 32;
    exp_41_ram[613] = 101;
    exp_41_ram[614] = 100;
    exp_41_ram[615] = 37;
    exp_41_ram[616] = 52;
    exp_41_ram[617] = 116;
    exp_41_ram[618] = 116;
    exp_41_ram[619] = 114;
    exp_41_ram[620] = 118;
    exp_41_ram[621] = 115;
    exp_41_ram[622] = 32;
    exp_41_ram[623] = 101;
    exp_41_ram[624] = 100;
    exp_41_ram[625] = 89;
    exp_41_ram[626] = 58;
    exp_41_ram[627] = 77;
    exp_41_ram[628] = 104;
    exp_41_ram[629] = 68;
    exp_41_ram[630] = 10;
    exp_41_ram[631] = 72;
    exp_41_ram[632] = 58;
    exp_41_ram[633] = 77;
    exp_41_ram[634] = 116;
    exp_41_ram[635] = 0;
    exp_41_ram[636] = 10;
    exp_41_ram[637] = 112;
    exp_41_ram[638] = 32;
    exp_41_ram[639] = 111;
    exp_41_ram[640] = 10;
    exp_41_ram[641] = 72;
    exp_41_ram[642] = 111;
    exp_41_ram[643] = 114;
    exp_41_ram[644] = 0;
    exp_41_ram[645] = 98;
    exp_41_ram[646] = 110;
    exp_41_ram[647] = 116;
    exp_41_ram[648] = 100;
    exp_41_ram[649] = 0;
    exp_41_ram[650] = 99;
    exp_41_ram[651] = 101;
    exp_41_ram[652] = 77;
    exp_41_ram[653] = 105;
    exp_41_ram[654] = 99;
    exp_41_ram[655] = 111;
    exp_41_ram[656] = 100;
    exp_41_ram[657] = 97;
    exp_41_ram[658] = 67;
    exp_41_ram[659] = 107;
    exp_41_ram[660] = 0;
    exp_41_ram[661] = 3;
    exp_41_ram[662] = 4;
    exp_41_ram[663] = 4;
    exp_41_ram[664] = 5;
    exp_41_ram[665] = 5;
    exp_41_ram[666] = 5;
    exp_41_ram[667] = 5;
    exp_41_ram[668] = 6;
    exp_41_ram[669] = 6;
    exp_41_ram[670] = 6;
    exp_41_ram[671] = 6;
    exp_41_ram[672] = 6;
    exp_41_ram[673] = 6;
    exp_41_ram[674] = 6;
    exp_41_ram[675] = 6;
    exp_41_ram[676] = 7;
    exp_41_ram[677] = 7;
    exp_41_ram[678] = 7;
    exp_41_ram[679] = 7;
    exp_41_ram[680] = 7;
    exp_41_ram[681] = 7;
    exp_41_ram[682] = 7;
    exp_41_ram[683] = 7;
    exp_41_ram[684] = 7;
    exp_41_ram[685] = 7;
    exp_41_ram[686] = 7;
    exp_41_ram[687] = 7;
    exp_41_ram[688] = 7;
    exp_41_ram[689] = 7;
    exp_41_ram[690] = 7;
    exp_41_ram[691] = 7;
    exp_41_ram[692] = 8;
    exp_41_ram[693] = 8;
    exp_41_ram[694] = 8;
    exp_41_ram[695] = 8;
    exp_41_ram[696] = 8;
    exp_41_ram[697] = 8;
    exp_41_ram[698] = 8;
    exp_41_ram[699] = 8;
    exp_41_ram[700] = 8;
    exp_41_ram[701] = 8;
    exp_41_ram[702] = 8;
    exp_41_ram[703] = 8;
    exp_41_ram[704] = 8;
    exp_41_ram[705] = 8;
    exp_41_ram[706] = 8;
    exp_41_ram[707] = 8;
    exp_41_ram[708] = 8;
    exp_41_ram[709] = 8;
    exp_41_ram[710] = 8;
    exp_41_ram[711] = 8;
    exp_41_ram[712] = 8;
    exp_41_ram[713] = 8;
    exp_41_ram[714] = 8;
    exp_41_ram[715] = 8;
    exp_41_ram[716] = 8;
    exp_41_ram[717] = 8;
    exp_41_ram[718] = 8;
    exp_41_ram[719] = 8;
    exp_41_ram[720] = 8;
    exp_41_ram[721] = 8;
    exp_41_ram[722] = 8;
    exp_41_ram[723] = 8;
    exp_41_ram[724] = 19;
    exp_41_ram[725] = 35;
    exp_41_ram[726] = 19;
    exp_41_ram[727] = 35;
    exp_41_ram[728] = 131;
    exp_41_ram[729] = 35;
    exp_41_ram[730] = 131;
    exp_41_ram[731] = 131;
    exp_41_ram[732] = 19;
    exp_41_ram[733] = 3;
    exp_41_ram[734] = 19;
    exp_41_ram[735] = 103;
    exp_41_ram[736] = 19;
    exp_41_ram[737] = 35;
    exp_41_ram[738] = 19;
    exp_41_ram[739] = 35;
    exp_41_ram[740] = 35;
    exp_41_ram[741] = 131;
    exp_41_ram[742] = 35;
    exp_41_ram[743] = 3;
    exp_41_ram[744] = 131;
    exp_41_ram[745] = 35;
    exp_41_ram[746] = 131;
    exp_41_ram[747] = 19;
    exp_41_ram[748] = 3;
    exp_41_ram[749] = 19;
    exp_41_ram[750] = 103;
    exp_41_ram[751] = 19;
    exp_41_ram[752] = 35;
    exp_41_ram[753] = 35;
    exp_41_ram[754] = 19;
    exp_41_ram[755] = 183;
    exp_41_ram[756] = 131;
    exp_41_ram[757] = 19;
    exp_41_ram[758] = 239;
    exp_41_ram[759] = 147;
    exp_41_ram[760] = 19;
    exp_41_ram[761] = 131;
    exp_41_ram[762] = 3;
    exp_41_ram[763] = 19;
    exp_41_ram[764] = 103;
    exp_41_ram[765] = 19;
    exp_41_ram[766] = 35;
    exp_41_ram[767] = 35;
    exp_41_ram[768] = 19;
    exp_41_ram[769] = 35;
    exp_41_ram[770] = 35;
    exp_41_ram[771] = 35;
    exp_41_ram[772] = 111;
    exp_41_ram[773] = 131;
    exp_41_ram[774] = 19;
    exp_41_ram[775] = 35;
    exp_41_ram[776] = 3;
    exp_41_ram[777] = 179;
    exp_41_ram[778] = 131;
    exp_41_ram[779] = 131;
    exp_41_ram[780] = 19;
    exp_41_ram[781] = 239;
    exp_41_ram[782] = 3;
    exp_41_ram[783] = 131;
    exp_41_ram[784] = 179;
    exp_41_ram[785] = 131;
    exp_41_ram[786] = 227;
    exp_41_ram[787] = 131;
    exp_41_ram[788] = 19;
    exp_41_ram[789] = 131;
    exp_41_ram[790] = 3;
    exp_41_ram[791] = 19;
    exp_41_ram[792] = 103;
    exp_41_ram[793] = 19;
    exp_41_ram[794] = 35;
    exp_41_ram[795] = 35;
    exp_41_ram[796] = 19;
    exp_41_ram[797] = 35;
    exp_41_ram[798] = 183;
    exp_41_ram[799] = 131;
    exp_41_ram[800] = 147;
    exp_41_ram[801] = 3;
    exp_41_ram[802] = 239;
    exp_41_ram[803] = 183;
    exp_41_ram[804] = 131;
    exp_41_ram[805] = 147;
    exp_41_ram[806] = 19;
    exp_41_ram[807] = 239;
    exp_41_ram[808] = 147;
    exp_41_ram[809] = 19;
    exp_41_ram[810] = 131;
    exp_41_ram[811] = 3;
    exp_41_ram[812] = 19;
    exp_41_ram[813] = 103;
    exp_41_ram[814] = 19;
    exp_41_ram[815] = 35;
    exp_41_ram[816] = 19;
    exp_41_ram[817] = 147;
    exp_41_ram[818] = 35;
    exp_41_ram[819] = 35;
    exp_41_ram[820] = 35;
    exp_41_ram[821] = 163;
    exp_41_ram[822] = 19;
    exp_41_ram[823] = 3;
    exp_41_ram[824] = 19;
    exp_41_ram[825] = 103;
    exp_41_ram[826] = 19;
    exp_41_ram[827] = 35;
    exp_41_ram[828] = 35;
    exp_41_ram[829] = 19;
    exp_41_ram[830] = 147;
    exp_41_ram[831] = 35;
    exp_41_ram[832] = 35;
    exp_41_ram[833] = 35;
    exp_41_ram[834] = 163;
    exp_41_ram[835] = 131;
    exp_41_ram[836] = 99;
    exp_41_ram[837] = 131;
    exp_41_ram[838] = 19;
    exp_41_ram[839] = 239;
    exp_41_ram[840] = 19;
    exp_41_ram[841] = 131;
    exp_41_ram[842] = 3;
    exp_41_ram[843] = 19;
    exp_41_ram[844] = 103;
    exp_41_ram[845] = 19;
    exp_41_ram[846] = 35;
    exp_41_ram[847] = 19;
    exp_41_ram[848] = 35;
    exp_41_ram[849] = 35;
    exp_41_ram[850] = 131;
    exp_41_ram[851] = 35;
    exp_41_ram[852] = 111;
    exp_41_ram[853] = 131;
    exp_41_ram[854] = 147;
    exp_41_ram[855] = 35;
    exp_41_ram[856] = 131;
    exp_41_ram[857] = 131;
    exp_41_ram[858] = 99;
    exp_41_ram[859] = 131;
    exp_41_ram[860] = 19;
    exp_41_ram[861] = 35;
    exp_41_ram[862] = 227;
    exp_41_ram[863] = 3;
    exp_41_ram[864] = 131;
    exp_41_ram[865] = 179;
    exp_41_ram[866] = 19;
    exp_41_ram[867] = 3;
    exp_41_ram[868] = 19;
    exp_41_ram[869] = 103;
    exp_41_ram[870] = 19;
    exp_41_ram[871] = 35;
    exp_41_ram[872] = 19;
    exp_41_ram[873] = 147;
    exp_41_ram[874] = 163;
    exp_41_ram[875] = 3;
    exp_41_ram[876] = 147;
    exp_41_ram[877] = 99;
    exp_41_ram[878] = 3;
    exp_41_ram[879] = 147;
    exp_41_ram[880] = 99;
    exp_41_ram[881] = 147;
    exp_41_ram[882] = 111;
    exp_41_ram[883] = 147;
    exp_41_ram[884] = 147;
    exp_41_ram[885] = 147;
    exp_41_ram[886] = 19;
    exp_41_ram[887] = 3;
    exp_41_ram[888] = 19;
    exp_41_ram[889] = 103;
    exp_41_ram[890] = 19;
    exp_41_ram[891] = 35;
    exp_41_ram[892] = 35;
    exp_41_ram[893] = 19;
    exp_41_ram[894] = 35;
    exp_41_ram[895] = 35;
    exp_41_ram[896] = 111;
    exp_41_ram[897] = 3;
    exp_41_ram[898] = 147;
    exp_41_ram[899] = 147;
    exp_41_ram[900] = 179;
    exp_41_ram[901] = 147;
    exp_41_ram[902] = 19;
    exp_41_ram[903] = 131;
    exp_41_ram[904] = 131;
    exp_41_ram[905] = 147;
    exp_41_ram[906] = 3;
    exp_41_ram[907] = 35;
    exp_41_ram[908] = 131;
    exp_41_ram[909] = 179;
    exp_41_ram[910] = 147;
    exp_41_ram[911] = 35;
    exp_41_ram[912] = 131;
    exp_41_ram[913] = 131;
    exp_41_ram[914] = 131;
    exp_41_ram[915] = 19;
    exp_41_ram[916] = 239;
    exp_41_ram[917] = 147;
    exp_41_ram[918] = 227;
    exp_41_ram[919] = 131;
    exp_41_ram[920] = 19;
    exp_41_ram[921] = 131;
    exp_41_ram[922] = 3;
    exp_41_ram[923] = 19;
    exp_41_ram[924] = 103;
    exp_41_ram[925] = 19;
    exp_41_ram[926] = 35;
    exp_41_ram[927] = 35;
    exp_41_ram[928] = 19;
    exp_41_ram[929] = 35;
    exp_41_ram[930] = 35;
    exp_41_ram[931] = 35;
    exp_41_ram[932] = 35;
    exp_41_ram[933] = 35;
    exp_41_ram[934] = 35;
    exp_41_ram[935] = 35;
    exp_41_ram[936] = 35;
    exp_41_ram[937] = 131;
    exp_41_ram[938] = 35;
    exp_41_ram[939] = 131;
    exp_41_ram[940] = 147;
    exp_41_ram[941] = 99;
    exp_41_ram[942] = 131;
    exp_41_ram[943] = 147;
    exp_41_ram[944] = 99;
    exp_41_ram[945] = 131;
    exp_41_ram[946] = 35;
    exp_41_ram[947] = 111;
    exp_41_ram[948] = 131;
    exp_41_ram[949] = 19;
    exp_41_ram[950] = 35;
    exp_41_ram[951] = 3;
    exp_41_ram[952] = 131;
    exp_41_ram[953] = 19;
    exp_41_ram[954] = 131;
    exp_41_ram[955] = 19;
    exp_41_ram[956] = 231;
    exp_41_ram[957] = 131;
    exp_41_ram[958] = 147;
    exp_41_ram[959] = 35;
    exp_41_ram[960] = 3;
    exp_41_ram[961] = 131;
    exp_41_ram[962] = 227;
    exp_41_ram[963] = 111;
    exp_41_ram[964] = 131;
    exp_41_ram[965] = 147;
    exp_41_ram[966] = 35;
    exp_41_ram[967] = 3;
    exp_41_ram[968] = 131;
    exp_41_ram[969] = 179;
    exp_41_ram[970] = 3;
    exp_41_ram[971] = 131;
    exp_41_ram[972] = 19;
    exp_41_ram[973] = 35;
    exp_41_ram[974] = 3;
    exp_41_ram[975] = 131;
    exp_41_ram[976] = 19;
    exp_41_ram[977] = 131;
    exp_41_ram[978] = 231;
    exp_41_ram[979] = 131;
    exp_41_ram[980] = 227;
    exp_41_ram[981] = 131;
    exp_41_ram[982] = 147;
    exp_41_ram[983] = 99;
    exp_41_ram[984] = 111;
    exp_41_ram[985] = 131;
    exp_41_ram[986] = 19;
    exp_41_ram[987] = 35;
    exp_41_ram[988] = 3;
    exp_41_ram[989] = 131;
    exp_41_ram[990] = 19;
    exp_41_ram[991] = 131;
    exp_41_ram[992] = 19;
    exp_41_ram[993] = 231;
    exp_41_ram[994] = 3;
    exp_41_ram[995] = 131;
    exp_41_ram[996] = 179;
    exp_41_ram[997] = 3;
    exp_41_ram[998] = 227;
    exp_41_ram[999] = 131;
    exp_41_ram[1000] = 19;
    exp_41_ram[1001] = 131;
    exp_41_ram[1002] = 3;
    exp_41_ram[1003] = 19;
    exp_41_ram[1004] = 103;
    exp_41_ram[1005] = 19;
    exp_41_ram[1006] = 35;
    exp_41_ram[1007] = 35;
    exp_41_ram[1008] = 19;
    exp_41_ram[1009] = 35;
    exp_41_ram[1010] = 35;
    exp_41_ram[1011] = 35;
    exp_41_ram[1012] = 35;
    exp_41_ram[1013] = 35;
    exp_41_ram[1014] = 35;
    exp_41_ram[1015] = 147;
    exp_41_ram[1016] = 35;
    exp_41_ram[1017] = 163;
    exp_41_ram[1018] = 131;
    exp_41_ram[1019] = 147;
    exp_41_ram[1020] = 99;
    exp_41_ram[1021] = 131;
    exp_41_ram[1022] = 99;
    exp_41_ram[1023] = 131;
    exp_41_ram[1024] = 147;
    exp_41_ram[1025] = 99;
    exp_41_ram[1026] = 131;
    exp_41_ram[1027] = 99;
    exp_41_ram[1028] = 131;
    exp_41_ram[1029] = 147;
    exp_41_ram[1030] = 99;
    exp_41_ram[1031] = 131;
    exp_41_ram[1032] = 147;
    exp_41_ram[1033] = 35;
    exp_41_ram[1034] = 111;
    exp_41_ram[1035] = 131;
    exp_41_ram[1036] = 19;
    exp_41_ram[1037] = 35;
    exp_41_ram[1038] = 3;
    exp_41_ram[1039] = 179;
    exp_41_ram[1040] = 19;
    exp_41_ram[1041] = 35;
    exp_41_ram[1042] = 3;
    exp_41_ram[1043] = 131;
    exp_41_ram[1044] = 99;
    exp_41_ram[1045] = 3;
    exp_41_ram[1046] = 147;
    exp_41_ram[1047] = 227;
    exp_41_ram[1048] = 111;
    exp_41_ram[1049] = 131;
    exp_41_ram[1050] = 19;
    exp_41_ram[1051] = 35;
    exp_41_ram[1052] = 3;
    exp_41_ram[1053] = 179;
    exp_41_ram[1054] = 19;
    exp_41_ram[1055] = 35;
    exp_41_ram[1056] = 131;
    exp_41_ram[1057] = 147;
    exp_41_ram[1058] = 99;
    exp_41_ram[1059] = 3;
    exp_41_ram[1060] = 131;
    exp_41_ram[1061] = 99;
    exp_41_ram[1062] = 3;
    exp_41_ram[1063] = 147;
    exp_41_ram[1064] = 227;
    exp_41_ram[1065] = 131;
    exp_41_ram[1066] = 147;
    exp_41_ram[1067] = 99;
    exp_41_ram[1068] = 131;
    exp_41_ram[1069] = 147;
    exp_41_ram[1070] = 99;
    exp_41_ram[1071] = 131;
    exp_41_ram[1072] = 99;
    exp_41_ram[1073] = 3;
    exp_41_ram[1074] = 131;
    exp_41_ram[1075] = 99;
    exp_41_ram[1076] = 3;
    exp_41_ram[1077] = 131;
    exp_41_ram[1078] = 99;
    exp_41_ram[1079] = 131;
    exp_41_ram[1080] = 147;
    exp_41_ram[1081] = 35;
    exp_41_ram[1082] = 131;
    exp_41_ram[1083] = 99;
    exp_41_ram[1084] = 3;
    exp_41_ram[1085] = 147;
    exp_41_ram[1086] = 99;
    exp_41_ram[1087] = 131;
    exp_41_ram[1088] = 147;
    exp_41_ram[1089] = 35;
    exp_41_ram[1090] = 3;
    exp_41_ram[1091] = 147;
    exp_41_ram[1092] = 99;
    exp_41_ram[1093] = 131;
    exp_41_ram[1094] = 147;
    exp_41_ram[1095] = 99;
    exp_41_ram[1096] = 3;
    exp_41_ram[1097] = 147;
    exp_41_ram[1098] = 99;
    exp_41_ram[1099] = 131;
    exp_41_ram[1100] = 19;
    exp_41_ram[1101] = 35;
    exp_41_ram[1102] = 3;
    exp_41_ram[1103] = 179;
    exp_41_ram[1104] = 19;
    exp_41_ram[1105] = 35;
    exp_41_ram[1106] = 111;
    exp_41_ram[1107] = 3;
    exp_41_ram[1108] = 147;
    exp_41_ram[1109] = 99;
    exp_41_ram[1110] = 131;
    exp_41_ram[1111] = 147;
    exp_41_ram[1112] = 99;
    exp_41_ram[1113] = 3;
    exp_41_ram[1114] = 147;
    exp_41_ram[1115] = 99;
    exp_41_ram[1116] = 131;
    exp_41_ram[1117] = 19;
    exp_41_ram[1118] = 35;
    exp_41_ram[1119] = 3;
    exp_41_ram[1120] = 179;
    exp_41_ram[1121] = 19;
    exp_41_ram[1122] = 35;
    exp_41_ram[1123] = 111;
    exp_41_ram[1124] = 3;
    exp_41_ram[1125] = 147;
    exp_41_ram[1126] = 99;
    exp_41_ram[1127] = 3;
    exp_41_ram[1128] = 147;
    exp_41_ram[1129] = 99;
    exp_41_ram[1130] = 131;
    exp_41_ram[1131] = 19;
    exp_41_ram[1132] = 35;
    exp_41_ram[1133] = 3;
    exp_41_ram[1134] = 179;
    exp_41_ram[1135] = 19;
    exp_41_ram[1136] = 35;
    exp_41_ram[1137] = 3;
    exp_41_ram[1138] = 147;
    exp_41_ram[1139] = 99;
    exp_41_ram[1140] = 131;
    exp_41_ram[1141] = 19;
    exp_41_ram[1142] = 35;
    exp_41_ram[1143] = 3;
    exp_41_ram[1144] = 179;
    exp_41_ram[1145] = 19;
    exp_41_ram[1146] = 35;
    exp_41_ram[1147] = 3;
    exp_41_ram[1148] = 147;
    exp_41_ram[1149] = 99;
    exp_41_ram[1150] = 131;
    exp_41_ram[1151] = 99;
    exp_41_ram[1152] = 131;
    exp_41_ram[1153] = 19;
    exp_41_ram[1154] = 35;
    exp_41_ram[1155] = 3;
    exp_41_ram[1156] = 179;
    exp_41_ram[1157] = 19;
    exp_41_ram[1158] = 35;
    exp_41_ram[1159] = 111;
    exp_41_ram[1160] = 131;
    exp_41_ram[1161] = 147;
    exp_41_ram[1162] = 99;
    exp_41_ram[1163] = 131;
    exp_41_ram[1164] = 19;
    exp_41_ram[1165] = 35;
    exp_41_ram[1166] = 3;
    exp_41_ram[1167] = 179;
    exp_41_ram[1168] = 19;
    exp_41_ram[1169] = 35;
    exp_41_ram[1170] = 111;
    exp_41_ram[1171] = 131;
    exp_41_ram[1172] = 147;
    exp_41_ram[1173] = 99;
    exp_41_ram[1174] = 131;
    exp_41_ram[1175] = 19;
    exp_41_ram[1176] = 35;
    exp_41_ram[1177] = 3;
    exp_41_ram[1178] = 179;
    exp_41_ram[1179] = 19;
    exp_41_ram[1180] = 35;
    exp_41_ram[1181] = 131;
    exp_41_ram[1182] = 3;
    exp_41_ram[1183] = 131;
    exp_41_ram[1184] = 3;
    exp_41_ram[1185] = 131;
    exp_41_ram[1186] = 3;
    exp_41_ram[1187] = 131;
    exp_41_ram[1188] = 3;
    exp_41_ram[1189] = 239;
    exp_41_ram[1190] = 147;
    exp_41_ram[1191] = 19;
    exp_41_ram[1192] = 131;
    exp_41_ram[1193] = 3;
    exp_41_ram[1194] = 19;
    exp_41_ram[1195] = 103;
    exp_41_ram[1196] = 19;
    exp_41_ram[1197] = 35;
    exp_41_ram[1198] = 35;
    exp_41_ram[1199] = 19;
    exp_41_ram[1200] = 35;
    exp_41_ram[1201] = 35;
    exp_41_ram[1202] = 35;
    exp_41_ram[1203] = 35;
    exp_41_ram[1204] = 35;
    exp_41_ram[1205] = 35;
    exp_41_ram[1206] = 35;
    exp_41_ram[1207] = 163;
    exp_41_ram[1208] = 35;
    exp_41_ram[1209] = 131;
    exp_41_ram[1210] = 99;
    exp_41_ram[1211] = 131;
    exp_41_ram[1212] = 147;
    exp_41_ram[1213] = 35;
    exp_41_ram[1214] = 131;
    exp_41_ram[1215] = 147;
    exp_41_ram[1216] = 99;
    exp_41_ram[1217] = 131;
    exp_41_ram[1218] = 99;
    exp_41_ram[1219] = 3;
    exp_41_ram[1220] = 131;
    exp_41_ram[1221] = 179;
    exp_41_ram[1222] = 163;
    exp_41_ram[1223] = 3;
    exp_41_ram[1224] = 147;
    exp_41_ram[1225] = 99;
    exp_41_ram[1226] = 131;
    exp_41_ram[1227] = 147;
    exp_41_ram[1228] = 147;
    exp_41_ram[1229] = 111;
    exp_41_ram[1230] = 131;
    exp_41_ram[1231] = 147;
    exp_41_ram[1232] = 99;
    exp_41_ram[1233] = 147;
    exp_41_ram[1234] = 111;
    exp_41_ram[1235] = 147;
    exp_41_ram[1236] = 3;
    exp_41_ram[1237] = 179;
    exp_41_ram[1238] = 147;
    exp_41_ram[1239] = 147;
    exp_41_ram[1240] = 147;
    exp_41_ram[1241] = 3;
    exp_41_ram[1242] = 147;
    exp_41_ram[1243] = 35;
    exp_41_ram[1244] = 147;
    exp_41_ram[1245] = 51;
    exp_41_ram[1246] = 35;
    exp_41_ram[1247] = 3;
    exp_41_ram[1248] = 131;
    exp_41_ram[1249] = 179;
    exp_41_ram[1250] = 35;
    exp_41_ram[1251] = 131;
    exp_41_ram[1252] = 99;
    exp_41_ram[1253] = 3;
    exp_41_ram[1254] = 147;
    exp_41_ram[1255] = 227;
    exp_41_ram[1256] = 131;
    exp_41_ram[1257] = 19;
    exp_41_ram[1258] = 131;
    exp_41_ram[1259] = 35;
    exp_41_ram[1260] = 131;
    exp_41_ram[1261] = 35;
    exp_41_ram[1262] = 131;
    exp_41_ram[1263] = 35;
    exp_41_ram[1264] = 131;
    exp_41_ram[1265] = 19;
    exp_41_ram[1266] = 131;
    exp_41_ram[1267] = 131;
    exp_41_ram[1268] = 3;
    exp_41_ram[1269] = 131;
    exp_41_ram[1270] = 3;
    exp_41_ram[1271] = 239;
    exp_41_ram[1272] = 147;
    exp_41_ram[1273] = 19;
    exp_41_ram[1274] = 131;
    exp_41_ram[1275] = 3;
    exp_41_ram[1276] = 19;
    exp_41_ram[1277] = 103;
    exp_41_ram[1278] = 19;
    exp_41_ram[1279] = 35;
    exp_41_ram[1280] = 35;
    exp_41_ram[1281] = 19;
    exp_41_ram[1282] = 35;
    exp_41_ram[1283] = 35;
    exp_41_ram[1284] = 35;
    exp_41_ram[1285] = 35;
    exp_41_ram[1286] = 35;
    exp_41_ram[1287] = 35;
    exp_41_ram[1288] = 131;
    exp_41_ram[1289] = 227;
    exp_41_ram[1290] = 183;
    exp_41_ram[1291] = 147;
    exp_41_ram[1292] = 35;
    exp_41_ram[1293] = 111;
    exp_41_ram[1294] = 131;
    exp_41_ram[1295] = 3;
    exp_41_ram[1296] = 147;
    exp_41_ram[1297] = 99;
    exp_41_ram[1298] = 131;
    exp_41_ram[1299] = 3;
    exp_41_ram[1300] = 131;
    exp_41_ram[1301] = 19;
    exp_41_ram[1302] = 35;
    exp_41_ram[1303] = 3;
    exp_41_ram[1304] = 131;
    exp_41_ram[1305] = 19;
    exp_41_ram[1306] = 131;
    exp_41_ram[1307] = 231;
    exp_41_ram[1308] = 131;
    exp_41_ram[1309] = 147;
    exp_41_ram[1310] = 35;
    exp_41_ram[1311] = 111;
    exp_41_ram[1312] = 131;
    exp_41_ram[1313] = 147;
    exp_41_ram[1314] = 35;
    exp_41_ram[1315] = 35;
    exp_41_ram[1316] = 131;
    exp_41_ram[1317] = 131;
    exp_41_ram[1318] = 147;
    exp_41_ram[1319] = 19;
    exp_41_ram[1320] = 99;
    exp_41_ram[1321] = 19;
    exp_41_ram[1322] = 183;
    exp_41_ram[1323] = 147;
    exp_41_ram[1324] = 179;
    exp_41_ram[1325] = 131;
    exp_41_ram[1326] = 103;
    exp_41_ram[1327] = 131;
    exp_41_ram[1328] = 147;
    exp_41_ram[1329] = 35;
    exp_41_ram[1330] = 131;
    exp_41_ram[1331] = 147;
    exp_41_ram[1332] = 35;
    exp_41_ram[1333] = 147;
    exp_41_ram[1334] = 35;
    exp_41_ram[1335] = 111;
    exp_41_ram[1336] = 131;
    exp_41_ram[1337] = 147;
    exp_41_ram[1338] = 35;
    exp_41_ram[1339] = 131;
    exp_41_ram[1340] = 147;
    exp_41_ram[1341] = 35;
    exp_41_ram[1342] = 147;
    exp_41_ram[1343] = 35;
    exp_41_ram[1344] = 111;
    exp_41_ram[1345] = 131;
    exp_41_ram[1346] = 147;
    exp_41_ram[1347] = 35;
    exp_41_ram[1348] = 131;
    exp_41_ram[1349] = 147;
    exp_41_ram[1350] = 35;
    exp_41_ram[1351] = 147;
    exp_41_ram[1352] = 35;
    exp_41_ram[1353] = 111;
    exp_41_ram[1354] = 131;
    exp_41_ram[1355] = 147;
    exp_41_ram[1356] = 35;
    exp_41_ram[1357] = 131;
    exp_41_ram[1358] = 147;
    exp_41_ram[1359] = 35;
    exp_41_ram[1360] = 147;
    exp_41_ram[1361] = 35;
    exp_41_ram[1362] = 111;
    exp_41_ram[1363] = 131;
    exp_41_ram[1364] = 147;
    exp_41_ram[1365] = 35;
    exp_41_ram[1366] = 131;
    exp_41_ram[1367] = 147;
    exp_41_ram[1368] = 35;
    exp_41_ram[1369] = 147;
    exp_41_ram[1370] = 35;
    exp_41_ram[1371] = 111;
    exp_41_ram[1372] = 35;
    exp_41_ram[1373] = 19;
    exp_41_ram[1374] = 131;
    exp_41_ram[1375] = 227;
    exp_41_ram[1376] = 35;
    exp_41_ram[1377] = 131;
    exp_41_ram[1378] = 131;
    exp_41_ram[1379] = 19;
    exp_41_ram[1380] = 239;
    exp_41_ram[1381] = 147;
    exp_41_ram[1382] = 99;
    exp_41_ram[1383] = 147;
    exp_41_ram[1384] = 19;
    exp_41_ram[1385] = 239;
    exp_41_ram[1386] = 35;
    exp_41_ram[1387] = 111;
    exp_41_ram[1388] = 131;
    exp_41_ram[1389] = 3;
    exp_41_ram[1390] = 147;
    exp_41_ram[1391] = 99;
    exp_41_ram[1392] = 131;
    exp_41_ram[1393] = 19;
    exp_41_ram[1394] = 35;
    exp_41_ram[1395] = 131;
    exp_41_ram[1396] = 35;
    exp_41_ram[1397] = 131;
    exp_41_ram[1398] = 99;
    exp_41_ram[1399] = 131;
    exp_41_ram[1400] = 147;
    exp_41_ram[1401] = 35;
    exp_41_ram[1402] = 131;
    exp_41_ram[1403] = 179;
    exp_41_ram[1404] = 35;
    exp_41_ram[1405] = 111;
    exp_41_ram[1406] = 131;
    exp_41_ram[1407] = 35;
    exp_41_ram[1408] = 131;
    exp_41_ram[1409] = 147;
    exp_41_ram[1410] = 35;
    exp_41_ram[1411] = 35;
    exp_41_ram[1412] = 131;
    exp_41_ram[1413] = 3;
    exp_41_ram[1414] = 147;
    exp_41_ram[1415] = 99;
    exp_41_ram[1416] = 131;
    exp_41_ram[1417] = 147;
    exp_41_ram[1418] = 35;
    exp_41_ram[1419] = 131;
    exp_41_ram[1420] = 147;
    exp_41_ram[1421] = 35;
    exp_41_ram[1422] = 131;
    exp_41_ram[1423] = 131;
    exp_41_ram[1424] = 19;
    exp_41_ram[1425] = 239;
    exp_41_ram[1426] = 147;
    exp_41_ram[1427] = 99;
    exp_41_ram[1428] = 147;
    exp_41_ram[1429] = 19;
    exp_41_ram[1430] = 239;
    exp_41_ram[1431] = 35;
    exp_41_ram[1432] = 111;
    exp_41_ram[1433] = 131;
    exp_41_ram[1434] = 3;
    exp_41_ram[1435] = 147;
    exp_41_ram[1436] = 99;
    exp_41_ram[1437] = 131;
    exp_41_ram[1438] = 19;
    exp_41_ram[1439] = 35;
    exp_41_ram[1440] = 131;
    exp_41_ram[1441] = 35;
    exp_41_ram[1442] = 131;
    exp_41_ram[1443] = 99;
    exp_41_ram[1444] = 147;
    exp_41_ram[1445] = 35;
    exp_41_ram[1446] = 131;
    exp_41_ram[1447] = 147;
    exp_41_ram[1448] = 35;
    exp_41_ram[1449] = 131;
    exp_41_ram[1450] = 131;
    exp_41_ram[1451] = 147;
    exp_41_ram[1452] = 19;
    exp_41_ram[1453] = 99;
    exp_41_ram[1454] = 19;
    exp_41_ram[1455] = 183;
    exp_41_ram[1456] = 147;
    exp_41_ram[1457] = 179;
    exp_41_ram[1458] = 131;
    exp_41_ram[1459] = 103;
    exp_41_ram[1460] = 131;
    exp_41_ram[1461] = 147;
    exp_41_ram[1462] = 35;
    exp_41_ram[1463] = 131;
    exp_41_ram[1464] = 147;
    exp_41_ram[1465] = 35;
    exp_41_ram[1466] = 131;
    exp_41_ram[1467] = 3;
    exp_41_ram[1468] = 147;
    exp_41_ram[1469] = 99;
    exp_41_ram[1470] = 131;
    exp_41_ram[1471] = 147;
    exp_41_ram[1472] = 35;
    exp_41_ram[1473] = 131;
    exp_41_ram[1474] = 147;
    exp_41_ram[1475] = 35;
    exp_41_ram[1476] = 111;
    exp_41_ram[1477] = 131;
    exp_41_ram[1478] = 147;
    exp_41_ram[1479] = 35;
    exp_41_ram[1480] = 131;
    exp_41_ram[1481] = 147;
    exp_41_ram[1482] = 35;
    exp_41_ram[1483] = 131;
    exp_41_ram[1484] = 3;
    exp_41_ram[1485] = 147;
    exp_41_ram[1486] = 99;
    exp_41_ram[1487] = 131;
    exp_41_ram[1488] = 147;
    exp_41_ram[1489] = 35;
    exp_41_ram[1490] = 131;
    exp_41_ram[1491] = 147;
    exp_41_ram[1492] = 35;
    exp_41_ram[1493] = 111;
    exp_41_ram[1494] = 131;
    exp_41_ram[1495] = 147;
    exp_41_ram[1496] = 35;
    exp_41_ram[1497] = 131;
    exp_41_ram[1498] = 147;
    exp_41_ram[1499] = 35;
    exp_41_ram[1500] = 111;
    exp_41_ram[1501] = 131;
    exp_41_ram[1502] = 147;
    exp_41_ram[1503] = 35;
    exp_41_ram[1504] = 131;
    exp_41_ram[1505] = 147;
    exp_41_ram[1506] = 35;
    exp_41_ram[1507] = 111;
    exp_41_ram[1508] = 131;
    exp_41_ram[1509] = 147;
    exp_41_ram[1510] = 35;
    exp_41_ram[1511] = 131;
    exp_41_ram[1512] = 147;
    exp_41_ram[1513] = 35;
    exp_41_ram[1514] = 111;
    exp_41_ram[1515] = 19;
    exp_41_ram[1516] = 111;
    exp_41_ram[1517] = 19;
    exp_41_ram[1518] = 111;
    exp_41_ram[1519] = 19;
    exp_41_ram[1520] = 131;
    exp_41_ram[1521] = 131;
    exp_41_ram[1522] = 147;
    exp_41_ram[1523] = 19;
    exp_41_ram[1524] = 99;
    exp_41_ram[1525] = 19;
    exp_41_ram[1526] = 183;
    exp_41_ram[1527] = 147;
    exp_41_ram[1528] = 179;
    exp_41_ram[1529] = 131;
    exp_41_ram[1530] = 103;
    exp_41_ram[1531] = 131;
    exp_41_ram[1532] = 3;
    exp_41_ram[1533] = 147;
    exp_41_ram[1534] = 99;
    exp_41_ram[1535] = 131;
    exp_41_ram[1536] = 3;
    exp_41_ram[1537] = 147;
    exp_41_ram[1538] = 99;
    exp_41_ram[1539] = 147;
    exp_41_ram[1540] = 35;
    exp_41_ram[1541] = 111;
    exp_41_ram[1542] = 131;
    exp_41_ram[1543] = 3;
    exp_41_ram[1544] = 147;
    exp_41_ram[1545] = 99;
    exp_41_ram[1546] = 147;
    exp_41_ram[1547] = 35;
    exp_41_ram[1548] = 111;
    exp_41_ram[1549] = 131;
    exp_41_ram[1550] = 3;
    exp_41_ram[1551] = 147;
    exp_41_ram[1552] = 99;
    exp_41_ram[1553] = 147;
    exp_41_ram[1554] = 35;
    exp_41_ram[1555] = 111;
    exp_41_ram[1556] = 147;
    exp_41_ram[1557] = 35;
    exp_41_ram[1558] = 131;
    exp_41_ram[1559] = 147;
    exp_41_ram[1560] = 35;
    exp_41_ram[1561] = 131;
    exp_41_ram[1562] = 3;
    exp_41_ram[1563] = 147;
    exp_41_ram[1564] = 99;
    exp_41_ram[1565] = 131;
    exp_41_ram[1566] = 147;
    exp_41_ram[1567] = 35;
    exp_41_ram[1568] = 131;
    exp_41_ram[1569] = 3;
    exp_41_ram[1570] = 147;
    exp_41_ram[1571] = 99;
    exp_41_ram[1572] = 131;
    exp_41_ram[1573] = 3;
    exp_41_ram[1574] = 147;
    exp_41_ram[1575] = 99;
    exp_41_ram[1576] = 131;
    exp_41_ram[1577] = 147;
    exp_41_ram[1578] = 35;
    exp_41_ram[1579] = 131;
    exp_41_ram[1580] = 147;
    exp_41_ram[1581] = 99;
    exp_41_ram[1582] = 131;
    exp_41_ram[1583] = 147;
    exp_41_ram[1584] = 35;
    exp_41_ram[1585] = 131;
    exp_41_ram[1586] = 3;
    exp_41_ram[1587] = 147;
    exp_41_ram[1588] = 99;
    exp_41_ram[1589] = 131;
    exp_41_ram[1590] = 3;
    exp_41_ram[1591] = 147;
    exp_41_ram[1592] = 99;
    exp_41_ram[1593] = 131;
    exp_41_ram[1594] = 147;
    exp_41_ram[1595] = 99;
    exp_41_ram[1596] = 131;
    exp_41_ram[1597] = 147;
    exp_41_ram[1598] = 99;
    exp_41_ram[1599] = 131;
    exp_41_ram[1600] = 19;
    exp_41_ram[1601] = 35;
    exp_41_ram[1602] = 131;
    exp_41_ram[1603] = 35;
    exp_41_ram[1604] = 131;
    exp_41_ram[1605] = 19;
    exp_41_ram[1606] = 131;
    exp_41_ram[1607] = 179;
    exp_41_ram[1608] = 179;
    exp_41_ram[1609] = 147;
    exp_41_ram[1610] = 131;
    exp_41_ram[1611] = 147;
    exp_41_ram[1612] = 19;
    exp_41_ram[1613] = 131;
    exp_41_ram[1614] = 35;
    exp_41_ram[1615] = 131;
    exp_41_ram[1616] = 35;
    exp_41_ram[1617] = 131;
    exp_41_ram[1618] = 3;
    exp_41_ram[1619] = 147;
    exp_41_ram[1620] = 19;
    exp_41_ram[1621] = 131;
    exp_41_ram[1622] = 3;
    exp_41_ram[1623] = 131;
    exp_41_ram[1624] = 3;
    exp_41_ram[1625] = 239;
    exp_41_ram[1626] = 35;
    exp_41_ram[1627] = 111;
    exp_41_ram[1628] = 131;
    exp_41_ram[1629] = 147;
    exp_41_ram[1630] = 99;
    exp_41_ram[1631] = 131;
    exp_41_ram[1632] = 19;
    exp_41_ram[1633] = 35;
    exp_41_ram[1634] = 131;
    exp_41_ram[1635] = 147;
    exp_41_ram[1636] = 111;
    exp_41_ram[1637] = 131;
    exp_41_ram[1638] = 147;
    exp_41_ram[1639] = 99;
    exp_41_ram[1640] = 131;
    exp_41_ram[1641] = 19;
    exp_41_ram[1642] = 35;
    exp_41_ram[1643] = 131;
    exp_41_ram[1644] = 147;
    exp_41_ram[1645] = 147;
    exp_41_ram[1646] = 111;
    exp_41_ram[1647] = 131;
    exp_41_ram[1648] = 19;
    exp_41_ram[1649] = 35;
    exp_41_ram[1650] = 131;
    exp_41_ram[1651] = 35;
    exp_41_ram[1652] = 131;
    exp_41_ram[1653] = 19;
    exp_41_ram[1654] = 131;
    exp_41_ram[1655] = 179;
    exp_41_ram[1656] = 179;
    exp_41_ram[1657] = 147;
    exp_41_ram[1658] = 131;
    exp_41_ram[1659] = 147;
    exp_41_ram[1660] = 19;
    exp_41_ram[1661] = 131;
    exp_41_ram[1662] = 35;
    exp_41_ram[1663] = 131;
    exp_41_ram[1664] = 35;
    exp_41_ram[1665] = 131;
    exp_41_ram[1666] = 3;
    exp_41_ram[1667] = 147;
    exp_41_ram[1668] = 19;
    exp_41_ram[1669] = 131;
    exp_41_ram[1670] = 3;
    exp_41_ram[1671] = 131;
    exp_41_ram[1672] = 3;
    exp_41_ram[1673] = 239;
    exp_41_ram[1674] = 35;
    exp_41_ram[1675] = 111;
    exp_41_ram[1676] = 131;
    exp_41_ram[1677] = 147;
    exp_41_ram[1678] = 99;
    exp_41_ram[1679] = 131;
    exp_41_ram[1680] = 147;
    exp_41_ram[1681] = 99;
    exp_41_ram[1682] = 131;
    exp_41_ram[1683] = 19;
    exp_41_ram[1684] = 35;
    exp_41_ram[1685] = 3;
    exp_41_ram[1686] = 131;
    exp_41_ram[1687] = 35;
    exp_41_ram[1688] = 131;
    exp_41_ram[1689] = 35;
    exp_41_ram[1690] = 131;
    exp_41_ram[1691] = 3;
    exp_41_ram[1692] = 147;
    exp_41_ram[1693] = 131;
    exp_41_ram[1694] = 3;
    exp_41_ram[1695] = 131;
    exp_41_ram[1696] = 3;
    exp_41_ram[1697] = 239;
    exp_41_ram[1698] = 35;
    exp_41_ram[1699] = 111;
    exp_41_ram[1700] = 131;
    exp_41_ram[1701] = 147;
    exp_41_ram[1702] = 99;
    exp_41_ram[1703] = 131;
    exp_41_ram[1704] = 19;
    exp_41_ram[1705] = 35;
    exp_41_ram[1706] = 131;
    exp_41_ram[1707] = 147;
    exp_41_ram[1708] = 111;
    exp_41_ram[1709] = 131;
    exp_41_ram[1710] = 147;
    exp_41_ram[1711] = 99;
    exp_41_ram[1712] = 131;
    exp_41_ram[1713] = 19;
    exp_41_ram[1714] = 35;
    exp_41_ram[1715] = 131;
    exp_41_ram[1716] = 147;
    exp_41_ram[1717] = 147;
    exp_41_ram[1718] = 111;
    exp_41_ram[1719] = 131;
    exp_41_ram[1720] = 19;
    exp_41_ram[1721] = 35;
    exp_41_ram[1722] = 131;
    exp_41_ram[1723] = 35;
    exp_41_ram[1724] = 131;
    exp_41_ram[1725] = 35;
    exp_41_ram[1726] = 131;
    exp_41_ram[1727] = 35;
    exp_41_ram[1728] = 131;
    exp_41_ram[1729] = 3;
    exp_41_ram[1730] = 147;
    exp_41_ram[1731] = 3;
    exp_41_ram[1732] = 131;
    exp_41_ram[1733] = 3;
    exp_41_ram[1734] = 131;
    exp_41_ram[1735] = 3;
    exp_41_ram[1736] = 239;
    exp_41_ram[1737] = 35;
    exp_41_ram[1738] = 131;
    exp_41_ram[1739] = 147;
    exp_41_ram[1740] = 35;
    exp_41_ram[1741] = 111;
    exp_41_ram[1742] = 147;
    exp_41_ram[1743] = 35;
    exp_41_ram[1744] = 131;
    exp_41_ram[1745] = 147;
    exp_41_ram[1746] = 99;
    exp_41_ram[1747] = 111;
    exp_41_ram[1748] = 131;
    exp_41_ram[1749] = 19;
    exp_41_ram[1750] = 35;
    exp_41_ram[1751] = 3;
    exp_41_ram[1752] = 131;
    exp_41_ram[1753] = 19;
    exp_41_ram[1754] = 131;
    exp_41_ram[1755] = 19;
    exp_41_ram[1756] = 231;
    exp_41_ram[1757] = 131;
    exp_41_ram[1758] = 19;
    exp_41_ram[1759] = 35;
    exp_41_ram[1760] = 3;
    exp_41_ram[1761] = 227;
    exp_41_ram[1762] = 131;
    exp_41_ram[1763] = 19;
    exp_41_ram[1764] = 35;
    exp_41_ram[1765] = 131;
    exp_41_ram[1766] = 19;
    exp_41_ram[1767] = 131;
    exp_41_ram[1768] = 19;
    exp_41_ram[1769] = 35;
    exp_41_ram[1770] = 3;
    exp_41_ram[1771] = 131;
    exp_41_ram[1772] = 19;
    exp_41_ram[1773] = 131;
    exp_41_ram[1774] = 231;
    exp_41_ram[1775] = 131;
    exp_41_ram[1776] = 147;
    exp_41_ram[1777] = 99;
    exp_41_ram[1778] = 111;
    exp_41_ram[1779] = 131;
    exp_41_ram[1780] = 19;
    exp_41_ram[1781] = 35;
    exp_41_ram[1782] = 3;
    exp_41_ram[1783] = 131;
    exp_41_ram[1784] = 19;
    exp_41_ram[1785] = 131;
    exp_41_ram[1786] = 19;
    exp_41_ram[1787] = 231;
    exp_41_ram[1788] = 131;
    exp_41_ram[1789] = 19;
    exp_41_ram[1790] = 35;
    exp_41_ram[1791] = 3;
    exp_41_ram[1792] = 227;
    exp_41_ram[1793] = 131;
    exp_41_ram[1794] = 147;
    exp_41_ram[1795] = 35;
    exp_41_ram[1796] = 111;
    exp_41_ram[1797] = 131;
    exp_41_ram[1798] = 19;
    exp_41_ram[1799] = 35;
    exp_41_ram[1800] = 131;
    exp_41_ram[1801] = 35;
    exp_41_ram[1802] = 131;
    exp_41_ram[1803] = 99;
    exp_41_ram[1804] = 131;
    exp_41_ram[1805] = 111;
    exp_41_ram[1806] = 147;
    exp_41_ram[1807] = 147;
    exp_41_ram[1808] = 3;
    exp_41_ram[1809] = 239;
    exp_41_ram[1810] = 35;
    exp_41_ram[1811] = 131;
    exp_41_ram[1812] = 147;
    exp_41_ram[1813] = 99;
    exp_41_ram[1814] = 3;
    exp_41_ram[1815] = 131;
    exp_41_ram[1816] = 99;
    exp_41_ram[1817] = 147;
    exp_41_ram[1818] = 35;
    exp_41_ram[1819] = 131;
    exp_41_ram[1820] = 147;
    exp_41_ram[1821] = 99;
    exp_41_ram[1822] = 111;
    exp_41_ram[1823] = 131;
    exp_41_ram[1824] = 19;
    exp_41_ram[1825] = 35;
    exp_41_ram[1826] = 3;
    exp_41_ram[1827] = 131;
    exp_41_ram[1828] = 19;
    exp_41_ram[1829] = 131;
    exp_41_ram[1830] = 19;
    exp_41_ram[1831] = 231;
    exp_41_ram[1832] = 131;
    exp_41_ram[1833] = 19;
    exp_41_ram[1834] = 35;
    exp_41_ram[1835] = 3;
    exp_41_ram[1836] = 227;
    exp_41_ram[1837] = 111;
    exp_41_ram[1838] = 131;
    exp_41_ram[1839] = 19;
    exp_41_ram[1840] = 35;
    exp_41_ram[1841] = 3;
    exp_41_ram[1842] = 131;
    exp_41_ram[1843] = 19;
    exp_41_ram[1844] = 35;
    exp_41_ram[1845] = 3;
    exp_41_ram[1846] = 131;
    exp_41_ram[1847] = 19;
    exp_41_ram[1848] = 131;
    exp_41_ram[1849] = 231;
    exp_41_ram[1850] = 131;
    exp_41_ram[1851] = 131;
    exp_41_ram[1852] = 99;
    exp_41_ram[1853] = 131;
    exp_41_ram[1854] = 147;
    exp_41_ram[1855] = 227;
    exp_41_ram[1856] = 131;
    exp_41_ram[1857] = 19;
    exp_41_ram[1858] = 35;
    exp_41_ram[1859] = 227;
    exp_41_ram[1860] = 131;
    exp_41_ram[1861] = 147;
    exp_41_ram[1862] = 99;
    exp_41_ram[1863] = 111;
    exp_41_ram[1864] = 131;
    exp_41_ram[1865] = 19;
    exp_41_ram[1866] = 35;
    exp_41_ram[1867] = 3;
    exp_41_ram[1868] = 131;
    exp_41_ram[1869] = 19;
    exp_41_ram[1870] = 131;
    exp_41_ram[1871] = 19;
    exp_41_ram[1872] = 231;
    exp_41_ram[1873] = 131;
    exp_41_ram[1874] = 19;
    exp_41_ram[1875] = 35;
    exp_41_ram[1876] = 3;
    exp_41_ram[1877] = 227;
    exp_41_ram[1878] = 131;
    exp_41_ram[1879] = 147;
    exp_41_ram[1880] = 35;
    exp_41_ram[1881] = 111;
    exp_41_ram[1882] = 147;
    exp_41_ram[1883] = 35;
    exp_41_ram[1884] = 131;
    exp_41_ram[1885] = 147;
    exp_41_ram[1886] = 35;
    exp_41_ram[1887] = 131;
    exp_41_ram[1888] = 19;
    exp_41_ram[1889] = 35;
    exp_41_ram[1890] = 131;
    exp_41_ram[1891] = 19;
    exp_41_ram[1892] = 131;
    exp_41_ram[1893] = 35;
    exp_41_ram[1894] = 131;
    exp_41_ram[1895] = 35;
    exp_41_ram[1896] = 131;
    exp_41_ram[1897] = 19;
    exp_41_ram[1898] = 147;
    exp_41_ram[1899] = 131;
    exp_41_ram[1900] = 3;
    exp_41_ram[1901] = 131;
    exp_41_ram[1902] = 3;
    exp_41_ram[1903] = 239;
    exp_41_ram[1904] = 35;
    exp_41_ram[1905] = 131;
    exp_41_ram[1906] = 147;
    exp_41_ram[1907] = 35;
    exp_41_ram[1908] = 111;
    exp_41_ram[1909] = 131;
    exp_41_ram[1910] = 19;
    exp_41_ram[1911] = 35;
    exp_41_ram[1912] = 3;
    exp_41_ram[1913] = 131;
    exp_41_ram[1914] = 19;
    exp_41_ram[1915] = 131;
    exp_41_ram[1916] = 19;
    exp_41_ram[1917] = 231;
    exp_41_ram[1918] = 131;
    exp_41_ram[1919] = 147;
    exp_41_ram[1920] = 35;
    exp_41_ram[1921] = 111;
    exp_41_ram[1922] = 131;
    exp_41_ram[1923] = 3;
    exp_41_ram[1924] = 131;
    exp_41_ram[1925] = 19;
    exp_41_ram[1926] = 35;
    exp_41_ram[1927] = 3;
    exp_41_ram[1928] = 131;
    exp_41_ram[1929] = 19;
    exp_41_ram[1930] = 131;
    exp_41_ram[1931] = 231;
    exp_41_ram[1932] = 131;
    exp_41_ram[1933] = 147;
    exp_41_ram[1934] = 35;
    exp_41_ram[1935] = 19;
    exp_41_ram[1936] = 131;
    exp_41_ram[1937] = 131;
    exp_41_ram[1938] = 99;
    exp_41_ram[1939] = 3;
    exp_41_ram[1940] = 131;
    exp_41_ram[1941] = 99;
    exp_41_ram[1942] = 131;
    exp_41_ram[1943] = 147;
    exp_41_ram[1944] = 111;
    exp_41_ram[1945] = 131;
    exp_41_ram[1946] = 3;
    exp_41_ram[1947] = 131;
    exp_41_ram[1948] = 19;
    exp_41_ram[1949] = 131;
    exp_41_ram[1950] = 19;
    exp_41_ram[1951] = 231;
    exp_41_ram[1952] = 131;
    exp_41_ram[1953] = 19;
    exp_41_ram[1954] = 131;
    exp_41_ram[1955] = 3;
    exp_41_ram[1956] = 19;
    exp_41_ram[1957] = 103;
    exp_41_ram[1958] = 19;
    exp_41_ram[1959] = 35;
    exp_41_ram[1960] = 35;
    exp_41_ram[1961] = 19;
    exp_41_ram[1962] = 35;
    exp_41_ram[1963] = 35;
    exp_41_ram[1964] = 35;
    exp_41_ram[1965] = 35;
    exp_41_ram[1966] = 35;
    exp_41_ram[1967] = 35;
    exp_41_ram[1968] = 35;
    exp_41_ram[1969] = 35;
    exp_41_ram[1970] = 147;
    exp_41_ram[1971] = 35;
    exp_41_ram[1972] = 131;
    exp_41_ram[1973] = 147;
    exp_41_ram[1974] = 35;
    exp_41_ram[1975] = 3;
    exp_41_ram[1976] = 147;
    exp_41_ram[1977] = 131;
    exp_41_ram[1978] = 19;
    exp_41_ram[1979] = 147;
    exp_41_ram[1980] = 183;
    exp_41_ram[1981] = 19;
    exp_41_ram[1982] = 239;
    exp_41_ram[1983] = 35;
    exp_41_ram[1984] = 131;
    exp_41_ram[1985] = 19;
    exp_41_ram[1986] = 131;
    exp_41_ram[1987] = 3;
    exp_41_ram[1988] = 19;
    exp_41_ram[1989] = 103;
    exp_41_ram[1990] = 19;
    exp_41_ram[1991] = 35;
    exp_41_ram[1992] = 35;
    exp_41_ram[1993] = 19;
    exp_41_ram[1994] = 147;
    exp_41_ram[1995] = 163;
    exp_41_ram[1996] = 3;
    exp_41_ram[1997] = 183;
    exp_41_ram[1998] = 131;
    exp_41_ram[1999] = 147;
    exp_41_ram[2000] = 19;
    exp_41_ram[2001] = 239;
    exp_41_ram[2002] = 19;
    exp_41_ram[2003] = 131;
    exp_41_ram[2004] = 3;
    exp_41_ram[2005] = 19;
    exp_41_ram[2006] = 103;
    exp_41_ram[2007] = 19;
    exp_41_ram[2008] = 35;
    exp_41_ram[2009] = 35;
    exp_41_ram[2010] = 35;
    exp_41_ram[2011] = 19;
    exp_41_ram[2012] = 147;
    exp_41_ram[2013] = 131;
    exp_41_ram[2014] = 35;
    exp_41_ram[2015] = 147;
    exp_41_ram[2016] = 35;
    exp_41_ram[2017] = 147;
    exp_41_ram[2018] = 35;
    exp_41_ram[2019] = 147;
    exp_41_ram[2020] = 35;
    exp_41_ram[2021] = 35;
    exp_41_ram[2022] = 35;
    exp_41_ram[2023] = 35;
    exp_41_ram[2024] = 3;
    exp_41_ram[2025] = 131;
    exp_41_ram[2026] = 3;
    exp_41_ram[2027] = 3;
    exp_41_ram[2028] = 131;
    exp_41_ram[2029] = 3;
    exp_41_ram[2030] = 131;
    exp_41_ram[2031] = 3;
    exp_41_ram[2032] = 131;
    exp_41_ram[2033] = 35;
    exp_41_ram[2034] = 35;
    exp_41_ram[2035] = 35;
    exp_41_ram[2036] = 35;
    exp_41_ram[2037] = 35;
    exp_41_ram[2038] = 35;
    exp_41_ram[2039] = 35;
    exp_41_ram[2040] = 35;
    exp_41_ram[2041] = 35;
    exp_41_ram[2042] = 147;
    exp_41_ram[2043] = 19;
    exp_41_ram[2044] = 239;
    exp_41_ram[2045] = 35;
    exp_41_ram[2046] = 35;
    exp_41_ram[2047] = 147;
    exp_41_ram[2048] = 131;
    exp_41_ram[2049] = 3;
    exp_41_ram[2050] = 19;
    exp_41_ram[2051] = 239;
    exp_41_ram[2052] = 3;
    exp_41_ram[2053] = 131;
    exp_41_ram[2054] = 179;
    exp_41_ram[2055] = 35;
    exp_41_ram[2056] = 3;
    exp_41_ram[2057] = 131;
    exp_41_ram[2058] = 3;
    exp_41_ram[2059] = 3;
    exp_41_ram[2060] = 131;
    exp_41_ram[2061] = 3;
    exp_41_ram[2062] = 131;
    exp_41_ram[2063] = 3;
    exp_41_ram[2064] = 131;
    exp_41_ram[2065] = 35;
    exp_41_ram[2066] = 35;
    exp_41_ram[2067] = 35;
    exp_41_ram[2068] = 35;
    exp_41_ram[2069] = 35;
    exp_41_ram[2070] = 35;
    exp_41_ram[2071] = 35;
    exp_41_ram[2072] = 35;
    exp_41_ram[2073] = 35;
    exp_41_ram[2074] = 147;
    exp_41_ram[2075] = 19;
    exp_41_ram[2076] = 239;
    exp_41_ram[2077] = 35;
    exp_41_ram[2078] = 35;
    exp_41_ram[2079] = 131;
    exp_41_ram[2080] = 35;
    exp_41_ram[2081] = 147;
    exp_41_ram[2082] = 35;
    exp_41_ram[2083] = 147;
    exp_41_ram[2084] = 35;
    exp_41_ram[2085] = 147;
    exp_41_ram[2086] = 35;
    exp_41_ram[2087] = 35;
    exp_41_ram[2088] = 35;
    exp_41_ram[2089] = 35;
    exp_41_ram[2090] = 3;
    exp_41_ram[2091] = 131;
    exp_41_ram[2092] = 3;
    exp_41_ram[2093] = 3;
    exp_41_ram[2094] = 131;
    exp_41_ram[2095] = 3;
    exp_41_ram[2096] = 131;
    exp_41_ram[2097] = 3;
    exp_41_ram[2098] = 131;
    exp_41_ram[2099] = 35;
    exp_41_ram[2100] = 35;
    exp_41_ram[2101] = 35;
    exp_41_ram[2102] = 35;
    exp_41_ram[2103] = 35;
    exp_41_ram[2104] = 35;
    exp_41_ram[2105] = 35;
    exp_41_ram[2106] = 35;
    exp_41_ram[2107] = 35;
    exp_41_ram[2108] = 147;
    exp_41_ram[2109] = 19;
    exp_41_ram[2110] = 239;
    exp_41_ram[2111] = 35;
    exp_41_ram[2112] = 35;
    exp_41_ram[2113] = 147;
    exp_41_ram[2114] = 131;
    exp_41_ram[2115] = 3;
    exp_41_ram[2116] = 19;
    exp_41_ram[2117] = 239;
    exp_41_ram[2118] = 3;
    exp_41_ram[2119] = 131;
    exp_41_ram[2120] = 179;
    exp_41_ram[2121] = 35;
    exp_41_ram[2122] = 3;
    exp_41_ram[2123] = 131;
    exp_41_ram[2124] = 3;
    exp_41_ram[2125] = 3;
    exp_41_ram[2126] = 131;
    exp_41_ram[2127] = 3;
    exp_41_ram[2128] = 131;
    exp_41_ram[2129] = 3;
    exp_41_ram[2130] = 131;
    exp_41_ram[2131] = 35;
    exp_41_ram[2132] = 35;
    exp_41_ram[2133] = 35;
    exp_41_ram[2134] = 35;
    exp_41_ram[2135] = 35;
    exp_41_ram[2136] = 35;
    exp_41_ram[2137] = 35;
    exp_41_ram[2138] = 35;
    exp_41_ram[2139] = 35;
    exp_41_ram[2140] = 147;
    exp_41_ram[2141] = 19;
    exp_41_ram[2142] = 239;
    exp_41_ram[2143] = 35;
    exp_41_ram[2144] = 35;
    exp_41_ram[2145] = 3;
    exp_41_ram[2146] = 131;
    exp_41_ram[2147] = 3;
    exp_41_ram[2148] = 3;
    exp_41_ram[2149] = 131;
    exp_41_ram[2150] = 3;
    exp_41_ram[2151] = 131;
    exp_41_ram[2152] = 3;
    exp_41_ram[2153] = 131;
    exp_41_ram[2154] = 35;
    exp_41_ram[2155] = 35;
    exp_41_ram[2156] = 35;
    exp_41_ram[2157] = 35;
    exp_41_ram[2158] = 35;
    exp_41_ram[2159] = 35;
    exp_41_ram[2160] = 35;
    exp_41_ram[2161] = 35;
    exp_41_ram[2162] = 35;
    exp_41_ram[2163] = 147;
    exp_41_ram[2164] = 19;
    exp_41_ram[2165] = 239;
    exp_41_ram[2166] = 35;
    exp_41_ram[2167] = 35;
    exp_41_ram[2168] = 3;
    exp_41_ram[2169] = 131;
    exp_41_ram[2170] = 99;
    exp_41_ram[2171] = 3;
    exp_41_ram[2172] = 131;
    exp_41_ram[2173] = 99;
    exp_41_ram[2174] = 3;
    exp_41_ram[2175] = 131;
    exp_41_ram[2176] = 99;
    exp_41_ram[2177] = 3;
    exp_41_ram[2178] = 131;
    exp_41_ram[2179] = 99;
    exp_41_ram[2180] = 3;
    exp_41_ram[2181] = 131;
    exp_41_ram[2182] = 99;
    exp_41_ram[2183] = 3;
    exp_41_ram[2184] = 131;
    exp_41_ram[2185] = 99;
    exp_41_ram[2186] = 147;
    exp_41_ram[2187] = 111;
    exp_41_ram[2188] = 147;
    exp_41_ram[2189] = 19;
    exp_41_ram[2190] = 131;
    exp_41_ram[2191] = 3;
    exp_41_ram[2192] = 131;
    exp_41_ram[2193] = 19;
    exp_41_ram[2194] = 103;
    exp_41_ram[2195] = 19;
    exp_41_ram[2196] = 35;
    exp_41_ram[2197] = 35;
    exp_41_ram[2198] = 19;
    exp_41_ram[2199] = 35;
    exp_41_ram[2200] = 35;
    exp_41_ram[2201] = 147;
    exp_41_ram[2202] = 131;
    exp_41_ram[2203] = 3;
    exp_41_ram[2204] = 19;
    exp_41_ram[2205] = 239;
    exp_41_ram[2206] = 3;
    exp_41_ram[2207] = 131;
    exp_41_ram[2208] = 3;
    exp_41_ram[2209] = 3;
    exp_41_ram[2210] = 131;
    exp_41_ram[2211] = 3;
    exp_41_ram[2212] = 131;
    exp_41_ram[2213] = 3;
    exp_41_ram[2214] = 131;
    exp_41_ram[2215] = 35;
    exp_41_ram[2216] = 35;
    exp_41_ram[2217] = 35;
    exp_41_ram[2218] = 35;
    exp_41_ram[2219] = 35;
    exp_41_ram[2220] = 35;
    exp_41_ram[2221] = 35;
    exp_41_ram[2222] = 35;
    exp_41_ram[2223] = 35;
    exp_41_ram[2224] = 147;
    exp_41_ram[2225] = 19;
    exp_41_ram[2226] = 239;
    exp_41_ram[2227] = 147;
    exp_41_ram[2228] = 19;
    exp_41_ram[2229] = 131;
    exp_41_ram[2230] = 3;
    exp_41_ram[2231] = 19;
    exp_41_ram[2232] = 103;
    exp_41_ram[2233] = 19;
    exp_41_ram[2234] = 35;
    exp_41_ram[2235] = 19;
    exp_41_ram[2236] = 183;
    exp_41_ram[2237] = 35;
    exp_41_ram[2238] = 183;
    exp_41_ram[2239] = 147;
    exp_41_ram[2240] = 35;
    exp_41_ram[2241] = 131;
    exp_41_ram[2242] = 131;
    exp_41_ram[2243] = 35;
    exp_41_ram[2244] = 35;
    exp_41_ram[2245] = 131;
    exp_41_ram[2246] = 147;
    exp_41_ram[2247] = 35;
    exp_41_ram[2248] = 35;
    exp_41_ram[2249] = 131;
    exp_41_ram[2250] = 131;
    exp_41_ram[2251] = 19;
    exp_41_ram[2252] = 147;
    exp_41_ram[2253] = 131;
    exp_41_ram[2254] = 179;
    exp_41_ram[2255] = 35;
    exp_41_ram[2256] = 131;
    exp_41_ram[2257] = 179;
    exp_41_ram[2258] = 35;
    exp_41_ram[2259] = 3;
    exp_41_ram[2260] = 131;
    exp_41_ram[2261] = 19;
    exp_41_ram[2262] = 147;
    exp_41_ram[2263] = 3;
    exp_41_ram[2264] = 19;
    exp_41_ram[2265] = 103;
    exp_41_ram[2266] = 19;
    exp_41_ram[2267] = 35;
    exp_41_ram[2268] = 35;
    exp_41_ram[2269] = 19;
    exp_41_ram[2270] = 35;
    exp_41_ram[2271] = 35;
    exp_41_ram[2272] = 35;
    exp_41_ram[2273] = 35;
    exp_41_ram[2274] = 3;
    exp_41_ram[2275] = 131;
    exp_41_ram[2276] = 3;
    exp_41_ram[2277] = 131;
    exp_41_ram[2278] = 51;
    exp_41_ram[2279] = 19;
    exp_41_ram[2280] = 51;
    exp_41_ram[2281] = 179;
    exp_41_ram[2282] = 179;
    exp_41_ram[2283] = 147;
    exp_41_ram[2284] = 19;
    exp_41_ram[2285] = 147;
    exp_41_ram[2286] = 19;
    exp_41_ram[2287] = 147;
    exp_41_ram[2288] = 239;
    exp_41_ram[2289] = 19;
    exp_41_ram[2290] = 147;
    exp_41_ram[2291] = 19;
    exp_41_ram[2292] = 147;
    exp_41_ram[2293] = 131;
    exp_41_ram[2294] = 3;
    exp_41_ram[2295] = 19;
    exp_41_ram[2296] = 103;
    exp_41_ram[2297] = 19;
    exp_41_ram[2298] = 35;
    exp_41_ram[2299] = 19;
    exp_41_ram[2300] = 35;
    exp_41_ram[2301] = 131;
    exp_41_ram[2302] = 147;
    exp_41_ram[2303] = 99;
    exp_41_ram[2304] = 3;
    exp_41_ram[2305] = 147;
    exp_41_ram[2306] = 179;
    exp_41_ram[2307] = 99;
    exp_41_ram[2308] = 3;
    exp_41_ram[2309] = 147;
    exp_41_ram[2310] = 179;
    exp_41_ram[2311] = 99;
    exp_41_ram[2312] = 147;
    exp_41_ram[2313] = 111;
    exp_41_ram[2314] = 147;
    exp_41_ram[2315] = 19;
    exp_41_ram[2316] = 3;
    exp_41_ram[2317] = 19;
    exp_41_ram[2318] = 103;
    exp_41_ram[2319] = 19;
    exp_41_ram[2320] = 35;
    exp_41_ram[2321] = 35;
    exp_41_ram[2322] = 19;
    exp_41_ram[2323] = 35;
    exp_41_ram[2324] = 3;
    exp_41_ram[2325] = 239;
    exp_41_ram[2326] = 147;
    exp_41_ram[2327] = 99;
    exp_41_ram[2328] = 147;
    exp_41_ram[2329] = 111;
    exp_41_ram[2330] = 147;
    exp_41_ram[2331] = 19;
    exp_41_ram[2332] = 131;
    exp_41_ram[2333] = 3;
    exp_41_ram[2334] = 19;
    exp_41_ram[2335] = 103;
    exp_41_ram[2336] = 19;
    exp_41_ram[2337] = 35;
    exp_41_ram[2338] = 35;
    exp_41_ram[2339] = 19;
    exp_41_ram[2340] = 35;
    exp_41_ram[2341] = 35;
    exp_41_ram[2342] = 3;
    exp_41_ram[2343] = 147;
    exp_41_ram[2344] = 99;
    exp_41_ram[2345] = 3;
    exp_41_ram[2346] = 147;
    exp_41_ram[2347] = 99;
    exp_41_ram[2348] = 3;
    exp_41_ram[2349] = 147;
    exp_41_ram[2350] = 99;
    exp_41_ram[2351] = 3;
    exp_41_ram[2352] = 147;
    exp_41_ram[2353] = 99;
    exp_41_ram[2354] = 147;
    exp_41_ram[2355] = 111;
    exp_41_ram[2356] = 3;
    exp_41_ram[2357] = 147;
    exp_41_ram[2358] = 99;
    exp_41_ram[2359] = 3;
    exp_41_ram[2360] = 239;
    exp_41_ram[2361] = 147;
    exp_41_ram[2362] = 99;
    exp_41_ram[2363] = 147;
    exp_41_ram[2364] = 111;
    exp_41_ram[2365] = 147;
    exp_41_ram[2366] = 111;
    exp_41_ram[2367] = 147;
    exp_41_ram[2368] = 19;
    exp_41_ram[2369] = 131;
    exp_41_ram[2370] = 3;
    exp_41_ram[2371] = 19;
    exp_41_ram[2372] = 103;
    exp_41_ram[2373] = 19;
    exp_41_ram[2374] = 35;
    exp_41_ram[2375] = 35;
    exp_41_ram[2376] = 35;
    exp_41_ram[2377] = 35;
    exp_41_ram[2378] = 35;
    exp_41_ram[2379] = 35;
    exp_41_ram[2380] = 35;
    exp_41_ram[2381] = 35;
    exp_41_ram[2382] = 35;
    exp_41_ram[2383] = 35;
    exp_41_ram[2384] = 35;
    exp_41_ram[2385] = 35;
    exp_41_ram[2386] = 35;
    exp_41_ram[2387] = 19;
    exp_41_ram[2388] = 147;
    exp_41_ram[2389] = 147;
    exp_41_ram[2390] = 19;
    exp_41_ram[2391] = 35;
    exp_41_ram[2392] = 35;
    exp_41_ram[2393] = 147;
    exp_41_ram[2394] = 35;
    exp_41_ram[2395] = 131;
    exp_41_ram[2396] = 35;
    exp_41_ram[2397] = 131;
    exp_41_ram[2398] = 147;
    exp_41_ram[2399] = 3;
    exp_41_ram[2400] = 99;
    exp_41_ram[2401] = 3;
    exp_41_ram[2402] = 239;
    exp_41_ram[2403] = 19;
    exp_41_ram[2404] = 183;
    exp_41_ram[2405] = 147;
    exp_41_ram[2406] = 179;
    exp_41_ram[2407] = 35;
    exp_41_ram[2408] = 35;
    exp_41_ram[2409] = 3;
    exp_41_ram[2410] = 131;
    exp_41_ram[2411] = 3;
    exp_41_ram[2412] = 131;
    exp_41_ram[2413] = 147;
    exp_41_ram[2414] = 51;
    exp_41_ram[2415] = 147;
    exp_41_ram[2416] = 179;
    exp_41_ram[2417] = 19;
    exp_41_ram[2418] = 179;
    exp_41_ram[2419] = 179;
    exp_41_ram[2420] = 147;
    exp_41_ram[2421] = 35;
    exp_41_ram[2422] = 35;
    exp_41_ram[2423] = 131;
    exp_41_ram[2424] = 147;
    exp_41_ram[2425] = 35;
    exp_41_ram[2426] = 111;
    exp_41_ram[2427] = 19;
    exp_41_ram[2428] = 35;
    exp_41_ram[2429] = 131;
    exp_41_ram[2430] = 19;
    exp_41_ram[2431] = 131;
    exp_41_ram[2432] = 99;
    exp_41_ram[2433] = 131;
    exp_41_ram[2434] = 3;
    exp_41_ram[2435] = 239;
    exp_41_ram[2436] = 19;
    exp_41_ram[2437] = 183;
    exp_41_ram[2438] = 147;
    exp_41_ram[2439] = 179;
    exp_41_ram[2440] = 19;
    exp_41_ram[2441] = 147;
    exp_41_ram[2442] = 3;
    exp_41_ram[2443] = 131;
    exp_41_ram[2444] = 51;
    exp_41_ram[2445] = 147;
    exp_41_ram[2446] = 179;
    exp_41_ram[2447] = 179;
    exp_41_ram[2448] = 179;
    exp_41_ram[2449] = 147;
    exp_41_ram[2450] = 35;
    exp_41_ram[2451] = 35;
    exp_41_ram[2452] = 131;
    exp_41_ram[2453] = 147;
    exp_41_ram[2454] = 35;
    exp_41_ram[2455] = 111;
    exp_41_ram[2456] = 19;
    exp_41_ram[2457] = 131;
    exp_41_ram[2458] = 19;
    exp_41_ram[2459] = 183;
    exp_41_ram[2460] = 147;
    exp_41_ram[2461] = 179;
    exp_41_ram[2462] = 19;
    exp_41_ram[2463] = 147;
    exp_41_ram[2464] = 147;
    exp_41_ram[2465] = 3;
    exp_41_ram[2466] = 131;
    exp_41_ram[2467] = 51;
    exp_41_ram[2468] = 147;
    exp_41_ram[2469] = 179;
    exp_41_ram[2470] = 179;
    exp_41_ram[2471] = 179;
    exp_41_ram[2472] = 147;
    exp_41_ram[2473] = 35;
    exp_41_ram[2474] = 35;
    exp_41_ram[2475] = 3;
    exp_41_ram[2476] = 183;
    exp_41_ram[2477] = 147;
    exp_41_ram[2478] = 179;
    exp_41_ram[2479] = 19;
    exp_41_ram[2480] = 147;
    exp_41_ram[2481] = 147;
    exp_41_ram[2482] = 3;
    exp_41_ram[2483] = 131;
    exp_41_ram[2484] = 51;
    exp_41_ram[2485] = 147;
    exp_41_ram[2486] = 179;
    exp_41_ram[2487] = 179;
    exp_41_ram[2488] = 179;
    exp_41_ram[2489] = 147;
    exp_41_ram[2490] = 35;
    exp_41_ram[2491] = 35;
    exp_41_ram[2492] = 3;
    exp_41_ram[2493] = 147;
    exp_41_ram[2494] = 147;
    exp_41_ram[2495] = 179;
    exp_41_ram[2496] = 147;
    exp_41_ram[2497] = 19;
    exp_41_ram[2498] = 147;
    exp_41_ram[2499] = 147;
    exp_41_ram[2500] = 3;
    exp_41_ram[2501] = 131;
    exp_41_ram[2502] = 51;
    exp_41_ram[2503] = 147;
    exp_41_ram[2504] = 179;
    exp_41_ram[2505] = 179;
    exp_41_ram[2506] = 179;
    exp_41_ram[2507] = 147;
    exp_41_ram[2508] = 35;
    exp_41_ram[2509] = 35;
    exp_41_ram[2510] = 131;
    exp_41_ram[2511] = 19;
    exp_41_ram[2512] = 147;
    exp_41_ram[2513] = 147;
    exp_41_ram[2514] = 3;
    exp_41_ram[2515] = 131;
    exp_41_ram[2516] = 51;
    exp_41_ram[2517] = 147;
    exp_41_ram[2518] = 179;
    exp_41_ram[2519] = 179;
    exp_41_ram[2520] = 179;
    exp_41_ram[2521] = 147;
    exp_41_ram[2522] = 35;
    exp_41_ram[2523] = 35;
    exp_41_ram[2524] = 3;
    exp_41_ram[2525] = 131;
    exp_41_ram[2526] = 19;
    exp_41_ram[2527] = 147;
    exp_41_ram[2528] = 131;
    exp_41_ram[2529] = 3;
    exp_41_ram[2530] = 131;
    exp_41_ram[2531] = 3;
    exp_41_ram[2532] = 131;
    exp_41_ram[2533] = 3;
    exp_41_ram[2534] = 131;
    exp_41_ram[2535] = 3;
    exp_41_ram[2536] = 131;
    exp_41_ram[2537] = 3;
    exp_41_ram[2538] = 131;
    exp_41_ram[2539] = 3;
    exp_41_ram[2540] = 131;
    exp_41_ram[2541] = 19;
    exp_41_ram[2542] = 103;
    exp_41_ram[2543] = 19;
    exp_41_ram[2544] = 35;
    exp_41_ram[2545] = 35;
    exp_41_ram[2546] = 35;
    exp_41_ram[2547] = 35;
    exp_41_ram[2548] = 35;
    exp_41_ram[2549] = 19;
    exp_41_ram[2550] = 35;
    exp_41_ram[2551] = 131;
    exp_41_ram[2552] = 3;
    exp_41_ram[2553] = 131;
    exp_41_ram[2554] = 3;
    exp_41_ram[2555] = 3;
    exp_41_ram[2556] = 131;
    exp_41_ram[2557] = 3;
    exp_41_ram[2558] = 131;
    exp_41_ram[2559] = 3;
    exp_41_ram[2560] = 131;
    exp_41_ram[2561] = 35;
    exp_41_ram[2562] = 35;
    exp_41_ram[2563] = 35;
    exp_41_ram[2564] = 35;
    exp_41_ram[2565] = 35;
    exp_41_ram[2566] = 35;
    exp_41_ram[2567] = 35;
    exp_41_ram[2568] = 35;
    exp_41_ram[2569] = 35;
    exp_41_ram[2570] = 3;
    exp_41_ram[2571] = 131;
    exp_41_ram[2572] = 3;
    exp_41_ram[2573] = 3;
    exp_41_ram[2574] = 131;
    exp_41_ram[2575] = 3;
    exp_41_ram[2576] = 131;
    exp_41_ram[2577] = 3;
    exp_41_ram[2578] = 131;
    exp_41_ram[2579] = 35;
    exp_41_ram[2580] = 35;
    exp_41_ram[2581] = 35;
    exp_41_ram[2582] = 35;
    exp_41_ram[2583] = 35;
    exp_41_ram[2584] = 35;
    exp_41_ram[2585] = 35;
    exp_41_ram[2586] = 35;
    exp_41_ram[2587] = 35;
    exp_41_ram[2588] = 147;
    exp_41_ram[2589] = 19;
    exp_41_ram[2590] = 239;
    exp_41_ram[2591] = 35;
    exp_41_ram[2592] = 35;
    exp_41_ram[2593] = 131;
    exp_41_ram[2594] = 99;
    exp_41_ram[2595] = 3;
    exp_41_ram[2596] = 131;
    exp_41_ram[2597] = 55;
    exp_41_ram[2598] = 19;
    exp_41_ram[2599] = 147;
    exp_41_ram[2600] = 51;
    exp_41_ram[2601] = 19;
    exp_41_ram[2602] = 51;
    exp_41_ram[2603] = 179;
    exp_41_ram[2604] = 179;
    exp_41_ram[2605] = 147;
    exp_41_ram[2606] = 35;
    exp_41_ram[2607] = 35;
    exp_41_ram[2608] = 111;
    exp_41_ram[2609] = 131;
    exp_41_ram[2610] = 99;
    exp_41_ram[2611] = 3;
    exp_41_ram[2612] = 131;
    exp_41_ram[2613] = 3;
    exp_41_ram[2614] = 3;
    exp_41_ram[2615] = 131;
    exp_41_ram[2616] = 3;
    exp_41_ram[2617] = 131;
    exp_41_ram[2618] = 3;
    exp_41_ram[2619] = 131;
    exp_41_ram[2620] = 35;
    exp_41_ram[2621] = 35;
    exp_41_ram[2622] = 35;
    exp_41_ram[2623] = 35;
    exp_41_ram[2624] = 35;
    exp_41_ram[2625] = 35;
    exp_41_ram[2626] = 35;
    exp_41_ram[2627] = 35;
    exp_41_ram[2628] = 35;
    exp_41_ram[2629] = 147;
    exp_41_ram[2630] = 19;
    exp_41_ram[2631] = 239;
    exp_41_ram[2632] = 147;
    exp_41_ram[2633] = 99;
    exp_41_ram[2634] = 55;
    exp_41_ram[2635] = 19;
    exp_41_ram[2636] = 147;
    exp_41_ram[2637] = 111;
    exp_41_ram[2638] = 19;
    exp_41_ram[2639] = 147;
    exp_41_ram[2640] = 3;
    exp_41_ram[2641] = 131;
    exp_41_ram[2642] = 51;
    exp_41_ram[2643] = 19;
    exp_41_ram[2644] = 51;
    exp_41_ram[2645] = 179;
    exp_41_ram[2646] = 179;
    exp_41_ram[2647] = 147;
    exp_41_ram[2648] = 35;
    exp_41_ram[2649] = 35;
    exp_41_ram[2650] = 111;
    exp_41_ram[2651] = 3;
    exp_41_ram[2652] = 131;
    exp_41_ram[2653] = 35;
    exp_41_ram[2654] = 35;
    exp_41_ram[2655] = 183;
    exp_41_ram[2656] = 131;
    exp_41_ram[2657] = 19;
    exp_41_ram[2658] = 147;
    exp_41_ram[2659] = 147;
    exp_41_ram[2660] = 3;
    exp_41_ram[2661] = 131;
    exp_41_ram[2662] = 51;
    exp_41_ram[2663] = 147;
    exp_41_ram[2664] = 179;
    exp_41_ram[2665] = 179;
    exp_41_ram[2666] = 179;
    exp_41_ram[2667] = 147;
    exp_41_ram[2668] = 35;
    exp_41_ram[2669] = 35;
    exp_41_ram[2670] = 131;
    exp_41_ram[2671] = 147;
    exp_41_ram[2672] = 131;
    exp_41_ram[2673] = 3;
    exp_41_ram[2674] = 19;
    exp_41_ram[2675] = 239;
    exp_41_ram[2676] = 3;
    exp_41_ram[2677] = 131;
    exp_41_ram[2678] = 3;
    exp_41_ram[2679] = 3;
    exp_41_ram[2680] = 131;
    exp_41_ram[2681] = 3;
    exp_41_ram[2682] = 131;
    exp_41_ram[2683] = 3;
    exp_41_ram[2684] = 131;
    exp_41_ram[2685] = 35;
    exp_41_ram[2686] = 35;
    exp_41_ram[2687] = 35;
    exp_41_ram[2688] = 35;
    exp_41_ram[2689] = 35;
    exp_41_ram[2690] = 35;
    exp_41_ram[2691] = 35;
    exp_41_ram[2692] = 35;
    exp_41_ram[2693] = 35;
    exp_41_ram[2694] = 131;
    exp_41_ram[2695] = 99;
    exp_41_ram[2696] = 131;
    exp_41_ram[2697] = 19;
    exp_41_ram[2698] = 35;
    exp_41_ram[2699] = 111;
    exp_41_ram[2700] = 131;
    exp_41_ram[2701] = 99;
    exp_41_ram[2702] = 3;
    exp_41_ram[2703] = 131;
    exp_41_ram[2704] = 3;
    exp_41_ram[2705] = 3;
    exp_41_ram[2706] = 131;
    exp_41_ram[2707] = 3;
    exp_41_ram[2708] = 131;
    exp_41_ram[2709] = 3;
    exp_41_ram[2710] = 131;
    exp_41_ram[2711] = 35;
    exp_41_ram[2712] = 35;
    exp_41_ram[2713] = 35;
    exp_41_ram[2714] = 35;
    exp_41_ram[2715] = 35;
    exp_41_ram[2716] = 35;
    exp_41_ram[2717] = 35;
    exp_41_ram[2718] = 35;
    exp_41_ram[2719] = 35;
    exp_41_ram[2720] = 147;
    exp_41_ram[2721] = 19;
    exp_41_ram[2722] = 239;
    exp_41_ram[2723] = 19;
    exp_41_ram[2724] = 131;
    exp_41_ram[2725] = 35;
    exp_41_ram[2726] = 111;
    exp_41_ram[2727] = 131;
    exp_41_ram[2728] = 35;
    exp_41_ram[2729] = 3;
    exp_41_ram[2730] = 131;
    exp_41_ram[2731] = 19;
    exp_41_ram[2732] = 147;
    exp_41_ram[2733] = 131;
    exp_41_ram[2734] = 3;
    exp_41_ram[2735] = 131;
    exp_41_ram[2736] = 3;
    exp_41_ram[2737] = 131;
    exp_41_ram[2738] = 19;
    exp_41_ram[2739] = 103;
    exp_41_ram[2740] = 19;
    exp_41_ram[2741] = 35;
    exp_41_ram[2742] = 35;
    exp_41_ram[2743] = 35;
    exp_41_ram[2744] = 35;
    exp_41_ram[2745] = 35;
    exp_41_ram[2746] = 35;
    exp_41_ram[2747] = 35;
    exp_41_ram[2748] = 35;
    exp_41_ram[2749] = 19;
    exp_41_ram[2750] = 35;
    exp_41_ram[2751] = 239;
    exp_41_ram[2752] = 19;
    exp_41_ram[2753] = 147;
    exp_41_ram[2754] = 183;
    exp_41_ram[2755] = 131;
    exp_41_ram[2756] = 19;
    exp_41_ram[2757] = 147;
    exp_41_ram[2758] = 19;
    exp_41_ram[2759] = 147;
    exp_41_ram[2760] = 19;
    exp_41_ram[2761] = 147;
    exp_41_ram[2762] = 239;
    exp_41_ram[2763] = 19;
    exp_41_ram[2764] = 147;
    exp_41_ram[2765] = 35;
    exp_41_ram[2766] = 183;
    exp_41_ram[2767] = 3;
    exp_41_ram[2768] = 131;
    exp_41_ram[2769] = 131;
    exp_41_ram[2770] = 179;
    exp_41_ram[2771] = 35;
    exp_41_ram[2772] = 131;
    exp_41_ram[2773] = 99;
    exp_41_ram[2774] = 131;
    exp_41_ram[2775] = 19;
    exp_41_ram[2776] = 147;
    exp_41_ram[2777] = 131;
    exp_41_ram[2778] = 35;
    exp_41_ram[2779] = 35;
    exp_41_ram[2780] = 131;
    exp_41_ram[2781] = 19;
    exp_41_ram[2782] = 147;
    exp_41_ram[2783] = 19;
    exp_41_ram[2784] = 147;
    exp_41_ram[2785] = 19;
    exp_41_ram[2786] = 147;
    exp_41_ram[2787] = 131;
    exp_41_ram[2788] = 3;
    exp_41_ram[2789] = 3;
    exp_41_ram[2790] = 131;
    exp_41_ram[2791] = 3;
    exp_41_ram[2792] = 131;
    exp_41_ram[2793] = 3;
    exp_41_ram[2794] = 131;
    exp_41_ram[2795] = 19;
    exp_41_ram[2796] = 103;
    exp_41_ram[2797] = 19;
    exp_41_ram[2798] = 35;
    exp_41_ram[2799] = 35;
    exp_41_ram[2800] = 35;
    exp_41_ram[2801] = 35;
    exp_41_ram[2802] = 19;
    exp_41_ram[2803] = 35;
    exp_41_ram[2804] = 35;
    exp_41_ram[2805] = 239;
    exp_41_ram[2806] = 19;
    exp_41_ram[2807] = 147;
    exp_41_ram[2808] = 183;
    exp_41_ram[2809] = 131;
    exp_41_ram[2810] = 19;
    exp_41_ram[2811] = 147;
    exp_41_ram[2812] = 19;
    exp_41_ram[2813] = 147;
    exp_41_ram[2814] = 19;
    exp_41_ram[2815] = 147;
    exp_41_ram[2816] = 239;
    exp_41_ram[2817] = 19;
    exp_41_ram[2818] = 147;
    exp_41_ram[2819] = 35;
    exp_41_ram[2820] = 35;
    exp_41_ram[2821] = 3;
    exp_41_ram[2822] = 131;
    exp_41_ram[2823] = 3;
    exp_41_ram[2824] = 131;
    exp_41_ram[2825] = 51;
    exp_41_ram[2826] = 19;
    exp_41_ram[2827] = 51;
    exp_41_ram[2828] = 179;
    exp_41_ram[2829] = 179;
    exp_41_ram[2830] = 147;
    exp_41_ram[2831] = 19;
    exp_41_ram[2832] = 147;
    exp_41_ram[2833] = 183;
    exp_41_ram[2834] = 35;
    exp_41_ram[2835] = 35;
    exp_41_ram[2836] = 19;
    exp_41_ram[2837] = 131;
    exp_41_ram[2838] = 3;
    exp_41_ram[2839] = 3;
    exp_41_ram[2840] = 131;
    exp_41_ram[2841] = 19;
    exp_41_ram[2842] = 103;
    exp_41_ram[2843] = 19;
    exp_41_ram[2844] = 35;
    exp_41_ram[2845] = 35;
    exp_41_ram[2846] = 19;
    exp_41_ram[2847] = 35;
    exp_41_ram[2848] = 183;
    exp_41_ram[2849] = 147;
    exp_41_ram[2850] = 3;
    exp_41_ram[2851] = 131;
    exp_41_ram[2852] = 3;
    exp_41_ram[2853] = 131;
    exp_41_ram[2854] = 3;
    exp_41_ram[2855] = 35;
    exp_41_ram[2856] = 35;
    exp_41_ram[2857] = 35;
    exp_41_ram[2858] = 35;
    exp_41_ram[2859] = 35;
    exp_41_ram[2860] = 131;
    exp_41_ram[2861] = 35;
    exp_41_ram[2862] = 183;
    exp_41_ram[2863] = 147;
    exp_41_ram[2864] = 3;
    exp_41_ram[2865] = 3;
    exp_41_ram[2866] = 131;
    exp_41_ram[2867] = 3;
    exp_41_ram[2868] = 3;
    exp_41_ram[2869] = 131;
    exp_41_ram[2870] = 3;
    exp_41_ram[2871] = 131;
    exp_41_ram[2872] = 3;
    exp_41_ram[2873] = 35;
    exp_41_ram[2874] = 35;
    exp_41_ram[2875] = 35;
    exp_41_ram[2876] = 35;
    exp_41_ram[2877] = 35;
    exp_41_ram[2878] = 35;
    exp_41_ram[2879] = 35;
    exp_41_ram[2880] = 35;
    exp_41_ram[2881] = 35;
    exp_41_ram[2882] = 131;
    exp_41_ram[2883] = 35;
    exp_41_ram[2884] = 35;
    exp_41_ram[2885] = 111;
    exp_41_ram[2886] = 131;
    exp_41_ram[2887] = 3;
    exp_41_ram[2888] = 147;
    exp_41_ram[2889] = 147;
    exp_41_ram[2890] = 51;
    exp_41_ram[2891] = 131;
    exp_41_ram[2892] = 179;
    exp_41_ram[2893] = 19;
    exp_41_ram[2894] = 179;
    exp_41_ram[2895] = 3;
    exp_41_ram[2896] = 183;
    exp_41_ram[2897] = 147;
    exp_41_ram[2898] = 131;
    exp_41_ram[2899] = 179;
    exp_41_ram[2900] = 35;
    exp_41_ram[2901] = 131;
    exp_41_ram[2902] = 147;
    exp_41_ram[2903] = 35;
    exp_41_ram[2904] = 3;
    exp_41_ram[2905] = 147;
    exp_41_ram[2906] = 227;
    exp_41_ram[2907] = 183;
    exp_41_ram[2908] = 147;
    exp_41_ram[2909] = 19;
    exp_41_ram[2910] = 163;
    exp_41_ram[2911] = 35;
    exp_41_ram[2912] = 111;
    exp_41_ram[2913] = 131;
    exp_41_ram[2914] = 3;
    exp_41_ram[2915] = 147;
    exp_41_ram[2916] = 147;
    exp_41_ram[2917] = 51;
    exp_41_ram[2918] = 131;
    exp_41_ram[2919] = 51;
    exp_41_ram[2920] = 131;
    exp_41_ram[2921] = 147;
    exp_41_ram[2922] = 147;
    exp_41_ram[2923] = 51;
    exp_41_ram[2924] = 3;
    exp_41_ram[2925] = 183;
    exp_41_ram[2926] = 147;
    exp_41_ram[2927] = 179;
    exp_41_ram[2928] = 35;
    exp_41_ram[2929] = 131;
    exp_41_ram[2930] = 147;
    exp_41_ram[2931] = 35;
    exp_41_ram[2932] = 3;
    exp_41_ram[2933] = 147;
    exp_41_ram[2934] = 227;
    exp_41_ram[2935] = 183;
    exp_41_ram[2936] = 147;
    exp_41_ram[2937] = 19;
    exp_41_ram[2938] = 163;
    exp_41_ram[2939] = 131;
    exp_41_ram[2940] = 131;
    exp_41_ram[2941] = 147;
    exp_41_ram[2942] = 19;
    exp_41_ram[2943] = 239;
    exp_41_ram[2944] = 19;
    exp_41_ram[2945] = 147;
    exp_41_ram[2946] = 35;
    exp_41_ram[2947] = 35;
    exp_41_ram[2948] = 131;
    exp_41_ram[2949] = 147;
    exp_41_ram[2950] = 147;
    exp_41_ram[2951] = 19;
    exp_41_ram[2952] = 183;
    exp_41_ram[2953] = 147;
    exp_41_ram[2954] = 35;
    exp_41_ram[2955] = 131;
    exp_41_ram[2956] = 147;
    exp_41_ram[2957] = 147;
    exp_41_ram[2958] = 19;
    exp_41_ram[2959] = 183;
    exp_41_ram[2960] = 147;
    exp_41_ram[2961] = 163;
    exp_41_ram[2962] = 183;
    exp_41_ram[2963] = 147;
    exp_41_ram[2964] = 19;
    exp_41_ram[2965] = 35;
    exp_41_ram[2966] = 131;
    exp_41_ram[2967] = 131;
    exp_41_ram[2968] = 147;
    exp_41_ram[2969] = 19;
    exp_41_ram[2970] = 239;
    exp_41_ram[2971] = 19;
    exp_41_ram[2972] = 147;
    exp_41_ram[2973] = 35;
    exp_41_ram[2974] = 35;
    exp_41_ram[2975] = 131;
    exp_41_ram[2976] = 147;
    exp_41_ram[2977] = 147;
    exp_41_ram[2978] = 19;
    exp_41_ram[2979] = 183;
    exp_41_ram[2980] = 147;
    exp_41_ram[2981] = 163;
    exp_41_ram[2982] = 131;
    exp_41_ram[2983] = 147;
    exp_41_ram[2984] = 147;
    exp_41_ram[2985] = 19;
    exp_41_ram[2986] = 183;
    exp_41_ram[2987] = 147;
    exp_41_ram[2988] = 35;
    exp_41_ram[2989] = 183;
    exp_41_ram[2990] = 147;
    exp_41_ram[2991] = 19;
    exp_41_ram[2992] = 163;
    exp_41_ram[2993] = 131;
    exp_41_ram[2994] = 131;
    exp_41_ram[2995] = 147;
    exp_41_ram[2996] = 19;
    exp_41_ram[2997] = 239;
    exp_41_ram[2998] = 19;
    exp_41_ram[2999] = 147;
    exp_41_ram[3000] = 35;
    exp_41_ram[3001] = 35;
    exp_41_ram[3002] = 131;
    exp_41_ram[3003] = 147;
    exp_41_ram[3004] = 147;
    exp_41_ram[3005] = 19;
    exp_41_ram[3006] = 183;
    exp_41_ram[3007] = 147;
    exp_41_ram[3008] = 35;
    exp_41_ram[3009] = 131;
    exp_41_ram[3010] = 147;
    exp_41_ram[3011] = 147;
    exp_41_ram[3012] = 19;
    exp_41_ram[3013] = 183;
    exp_41_ram[3014] = 147;
    exp_41_ram[3015] = 163;
    exp_41_ram[3016] = 183;
    exp_41_ram[3017] = 147;
    exp_41_ram[3018] = 19;
    exp_41_ram[3019] = 35;
    exp_41_ram[3020] = 131;
    exp_41_ram[3021] = 131;
    exp_41_ram[3022] = 147;
    exp_41_ram[3023] = 19;
    exp_41_ram[3024] = 239;
    exp_41_ram[3025] = 19;
    exp_41_ram[3026] = 147;
    exp_41_ram[3027] = 35;
    exp_41_ram[3028] = 35;
    exp_41_ram[3029] = 131;
    exp_41_ram[3030] = 147;
    exp_41_ram[3031] = 147;
    exp_41_ram[3032] = 19;
    exp_41_ram[3033] = 183;
    exp_41_ram[3034] = 147;
    exp_41_ram[3035] = 163;
    exp_41_ram[3036] = 131;
    exp_41_ram[3037] = 147;
    exp_41_ram[3038] = 147;
    exp_41_ram[3039] = 19;
    exp_41_ram[3040] = 183;
    exp_41_ram[3041] = 147;
    exp_41_ram[3042] = 35;
    exp_41_ram[3043] = 183;
    exp_41_ram[3044] = 147;
    exp_41_ram[3045] = 19;
    exp_41_ram[3046] = 163;
    exp_41_ram[3047] = 131;
    exp_41_ram[3048] = 131;
    exp_41_ram[3049] = 147;
    exp_41_ram[3050] = 147;
    exp_41_ram[3051] = 19;
    exp_41_ram[3052] = 239;
    exp_41_ram[3053] = 19;
    exp_41_ram[3054] = 147;
    exp_41_ram[3055] = 35;
    exp_41_ram[3056] = 35;
    exp_41_ram[3057] = 131;
    exp_41_ram[3058] = 147;
    exp_41_ram[3059] = 147;
    exp_41_ram[3060] = 19;
    exp_41_ram[3061] = 183;
    exp_41_ram[3062] = 147;
    exp_41_ram[3063] = 35;
    exp_41_ram[3064] = 131;
    exp_41_ram[3065] = 147;
    exp_41_ram[3066] = 19;
    exp_41_ram[3067] = 239;
    exp_41_ram[3068] = 19;
    exp_41_ram[3069] = 147;
    exp_41_ram[3070] = 35;
    exp_41_ram[3071] = 35;
    exp_41_ram[3072] = 131;
    exp_41_ram[3073] = 147;
    exp_41_ram[3074] = 147;
    exp_41_ram[3075] = 19;
    exp_41_ram[3076] = 183;
    exp_41_ram[3077] = 147;
    exp_41_ram[3078] = 163;
    exp_41_ram[3079] = 131;
    exp_41_ram[3080] = 147;
    exp_41_ram[3081] = 19;
    exp_41_ram[3082] = 239;
    exp_41_ram[3083] = 19;
    exp_41_ram[3084] = 147;
    exp_41_ram[3085] = 35;
    exp_41_ram[3086] = 35;
    exp_41_ram[3087] = 131;
    exp_41_ram[3088] = 147;
    exp_41_ram[3089] = 147;
    exp_41_ram[3090] = 19;
    exp_41_ram[3091] = 183;
    exp_41_ram[3092] = 147;
    exp_41_ram[3093] = 35;
    exp_41_ram[3094] = 131;
    exp_41_ram[3095] = 147;
    exp_41_ram[3096] = 147;
    exp_41_ram[3097] = 19;
    exp_41_ram[3098] = 183;
    exp_41_ram[3099] = 147;
    exp_41_ram[3100] = 163;
    exp_41_ram[3101] = 183;
    exp_41_ram[3102] = 147;
    exp_41_ram[3103] = 19;
    exp_41_ram[3104] = 35;
    exp_41_ram[3105] = 183;
    exp_41_ram[3106] = 147;
    exp_41_ram[3107] = 163;
    exp_41_ram[3108] = 183;
    exp_41_ram[3109] = 147;
    exp_41_ram[3110] = 19;
    exp_41_ram[3111] = 131;
    exp_41_ram[3112] = 3;
    exp_41_ram[3113] = 19;
    exp_41_ram[3114] = 103;
    exp_41_ram[3115] = 19;
    exp_41_ram[3116] = 35;
    exp_41_ram[3117] = 35;
    exp_41_ram[3118] = 19;
    exp_41_ram[3119] = 35;
    exp_41_ram[3120] = 3;
    exp_41_ram[3121] = 239;
    exp_41_ram[3122] = 147;
    exp_41_ram[3123] = 19;
    exp_41_ram[3124] = 239;
    exp_41_ram[3125] = 147;
    exp_41_ram[3126] = 19;
    exp_41_ram[3127] = 131;
    exp_41_ram[3128] = 3;
    exp_41_ram[3129] = 19;
    exp_41_ram[3130] = 103;
    exp_41_ram[3131] = 19;
    exp_41_ram[3132] = 35;
    exp_41_ram[3133] = 35;
    exp_41_ram[3134] = 35;
    exp_41_ram[3135] = 35;
    exp_41_ram[3136] = 35;
    exp_41_ram[3137] = 35;
    exp_41_ram[3138] = 35;
    exp_41_ram[3139] = 35;
    exp_41_ram[3140] = 35;
    exp_41_ram[3141] = 35;
    exp_41_ram[3142] = 19;
    exp_41_ram[3143] = 35;
    exp_41_ram[3144] = 35;
    exp_41_ram[3145] = 35;
    exp_41_ram[3146] = 147;
    exp_41_ram[3147] = 35;
    exp_41_ram[3148] = 147;
    exp_41_ram[3149] = 35;
    exp_41_ram[3150] = 131;
    exp_41_ram[3151] = 19;
    exp_41_ram[3152] = 239;
    exp_41_ram[3153] = 35;
    exp_41_ram[3154] = 3;
    exp_41_ram[3155] = 183;
    exp_41_ram[3156] = 147;
    exp_41_ram[3157] = 179;
    exp_41_ram[3158] = 35;
    exp_41_ram[3159] = 131;
    exp_41_ram[3160] = 19;
    exp_41_ram[3161] = 147;
    exp_41_ram[3162] = 131;
    exp_41_ram[3163] = 19;
    exp_41_ram[3164] = 99;
    exp_41_ram[3165] = 131;
    exp_41_ram[3166] = 19;
    exp_41_ram[3167] = 99;
    exp_41_ram[3168] = 131;
    exp_41_ram[3169] = 19;
    exp_41_ram[3170] = 99;
    exp_41_ram[3171] = 131;
    exp_41_ram[3172] = 147;
    exp_41_ram[3173] = 35;
    exp_41_ram[3174] = 131;
    exp_41_ram[3175] = 19;
    exp_41_ram[3176] = 131;
    exp_41_ram[3177] = 179;
    exp_41_ram[3178] = 35;
    exp_41_ram[3179] = 131;
    exp_41_ram[3180] = 19;
    exp_41_ram[3181] = 147;
    exp_41_ram[3182] = 3;
    exp_41_ram[3183] = 131;
    exp_41_ram[3184] = 51;
    exp_41_ram[3185] = 147;
    exp_41_ram[3186] = 179;
    exp_41_ram[3187] = 179;
    exp_41_ram[3188] = 179;
    exp_41_ram[3189] = 147;
    exp_41_ram[3190] = 35;
    exp_41_ram[3191] = 35;
    exp_41_ram[3192] = 111;
    exp_41_ram[3193] = 19;
    exp_41_ram[3194] = 35;
    exp_41_ram[3195] = 35;
    exp_41_ram[3196] = 131;
    exp_41_ram[3197] = 19;
    exp_41_ram[3198] = 131;
    exp_41_ram[3199] = 147;
    exp_41_ram[3200] = 19;
    exp_41_ram[3201] = 239;
    exp_41_ram[3202] = 35;
    exp_41_ram[3203] = 3;
    exp_41_ram[3204] = 183;
    exp_41_ram[3205] = 147;
    exp_41_ram[3206] = 179;
    exp_41_ram[3207] = 35;
    exp_41_ram[3208] = 131;
    exp_41_ram[3209] = 19;
    exp_41_ram[3210] = 147;
    exp_41_ram[3211] = 131;
    exp_41_ram[3212] = 19;
    exp_41_ram[3213] = 99;
    exp_41_ram[3214] = 131;
    exp_41_ram[3215] = 19;
    exp_41_ram[3216] = 99;
    exp_41_ram[3217] = 131;
    exp_41_ram[3218] = 19;
    exp_41_ram[3219] = 99;
    exp_41_ram[3220] = 131;
    exp_41_ram[3221] = 147;
    exp_41_ram[3222] = 35;
    exp_41_ram[3223] = 131;
    exp_41_ram[3224] = 19;
    exp_41_ram[3225] = 131;
    exp_41_ram[3226] = 179;
    exp_41_ram[3227] = 35;
    exp_41_ram[3228] = 131;
    exp_41_ram[3229] = 19;
    exp_41_ram[3230] = 131;
    exp_41_ram[3231] = 179;
    exp_41_ram[3232] = 35;
    exp_41_ram[3233] = 131;
    exp_41_ram[3234] = 19;
    exp_41_ram[3235] = 147;
    exp_41_ram[3236] = 3;
    exp_41_ram[3237] = 131;
    exp_41_ram[3238] = 51;
    exp_41_ram[3239] = 147;
    exp_41_ram[3240] = 179;
    exp_41_ram[3241] = 179;
    exp_41_ram[3242] = 179;
    exp_41_ram[3243] = 147;
    exp_41_ram[3244] = 35;
    exp_41_ram[3245] = 35;
    exp_41_ram[3246] = 111;
    exp_41_ram[3247] = 19;
    exp_41_ram[3248] = 131;
    exp_41_ram[3249] = 147;
    exp_41_ram[3250] = 35;
    exp_41_ram[3251] = 3;
    exp_41_ram[3252] = 183;
    exp_41_ram[3253] = 147;
    exp_41_ram[3254] = 19;
    exp_41_ram[3255] = 239;
    exp_41_ram[3256] = 19;
    exp_41_ram[3257] = 147;
    exp_41_ram[3258] = 35;
    exp_41_ram[3259] = 35;
    exp_41_ram[3260] = 131;
    exp_41_ram[3261] = 147;
    exp_41_ram[3262] = 35;
    exp_41_ram[3263] = 3;
    exp_41_ram[3264] = 131;
    exp_41_ram[3265] = 179;
    exp_41_ram[3266] = 35;
    exp_41_ram[3267] = 3;
    exp_41_ram[3268] = 147;
    exp_41_ram[3269] = 179;
    exp_41_ram[3270] = 35;
    exp_41_ram[3271] = 3;
    exp_41_ram[3272] = 131;
    exp_41_ram[3273] = 179;
    exp_41_ram[3274] = 35;
    exp_41_ram[3275] = 131;
    exp_41_ram[3276] = 35;
    exp_41_ram[3277] = 147;
    exp_41_ram[3278] = 35;
    exp_41_ram[3279] = 3;
    exp_41_ram[3280] = 183;
    exp_41_ram[3281] = 147;
    exp_41_ram[3282] = 19;
    exp_41_ram[3283] = 239;
    exp_41_ram[3284] = 19;
    exp_41_ram[3285] = 147;
    exp_41_ram[3286] = 35;
    exp_41_ram[3287] = 35;
    exp_41_ram[3288] = 131;
    exp_41_ram[3289] = 35;
    exp_41_ram[3290] = 131;
    exp_41_ram[3291] = 35;
    exp_41_ram[3292] = 147;
    exp_41_ram[3293] = 35;
    exp_41_ram[3294] = 131;
    exp_41_ram[3295] = 147;
    exp_41_ram[3296] = 19;
    exp_41_ram[3297] = 239;
    exp_41_ram[3298] = 19;
    exp_41_ram[3299] = 147;
    exp_41_ram[3300] = 35;
    exp_41_ram[3301] = 35;
    exp_41_ram[3302] = 131;
    exp_41_ram[3303] = 35;
    exp_41_ram[3304] = 131;
    exp_41_ram[3305] = 35;
    exp_41_ram[3306] = 147;
    exp_41_ram[3307] = 35;
    exp_41_ram[3308] = 131;
    exp_41_ram[3309] = 35;
    exp_41_ram[3310] = 131;
    exp_41_ram[3311] = 3;
    exp_41_ram[3312] = 3;
    exp_41_ram[3313] = 131;
    exp_41_ram[3314] = 3;
    exp_41_ram[3315] = 3;
    exp_41_ram[3316] = 131;
    exp_41_ram[3317] = 3;
    exp_41_ram[3318] = 131;
    exp_41_ram[3319] = 3;
    exp_41_ram[3320] = 35;
    exp_41_ram[3321] = 35;
    exp_41_ram[3322] = 35;
    exp_41_ram[3323] = 35;
    exp_41_ram[3324] = 35;
    exp_41_ram[3325] = 35;
    exp_41_ram[3326] = 35;
    exp_41_ram[3327] = 35;
    exp_41_ram[3328] = 35;
    exp_41_ram[3329] = 3;
    exp_41_ram[3330] = 131;
    exp_41_ram[3331] = 3;
    exp_41_ram[3332] = 3;
    exp_41_ram[3333] = 131;
    exp_41_ram[3334] = 3;
    exp_41_ram[3335] = 131;
    exp_41_ram[3336] = 3;
    exp_41_ram[3337] = 131;
    exp_41_ram[3338] = 3;
    exp_41_ram[3339] = 131;
    exp_41_ram[3340] = 19;
    exp_41_ram[3341] = 103;
    exp_41_ram[3342] = 19;
    exp_41_ram[3343] = 35;
    exp_41_ram[3344] = 35;
    exp_41_ram[3345] = 35;
    exp_41_ram[3346] = 35;
    exp_41_ram[3347] = 35;
    exp_41_ram[3348] = 19;
    exp_41_ram[3349] = 35;
    exp_41_ram[3350] = 147;
    exp_41_ram[3351] = 19;
    exp_41_ram[3352] = 35;
    exp_41_ram[3353] = 35;
    exp_41_ram[3354] = 131;
    exp_41_ram[3355] = 3;
    exp_41_ram[3356] = 131;
    exp_41_ram[3357] = 35;
    exp_41_ram[3358] = 35;
    exp_41_ram[3359] = 3;
    exp_41_ram[3360] = 131;
    exp_41_ram[3361] = 239;
    exp_41_ram[3362] = 147;
    exp_41_ram[3363] = 99;
    exp_41_ram[3364] = 55;
    exp_41_ram[3365] = 19;
    exp_41_ram[3366] = 147;
    exp_41_ram[3367] = 35;
    exp_41_ram[3368] = 35;
    exp_41_ram[3369] = 183;
    exp_41_ram[3370] = 131;
    exp_41_ram[3371] = 19;
    exp_41_ram[3372] = 147;
    exp_41_ram[3373] = 147;
    exp_41_ram[3374] = 3;
    exp_41_ram[3375] = 131;
    exp_41_ram[3376] = 51;
    exp_41_ram[3377] = 147;
    exp_41_ram[3378] = 179;
    exp_41_ram[3379] = 179;
    exp_41_ram[3380] = 179;
    exp_41_ram[3381] = 147;
    exp_41_ram[3382] = 19;
    exp_41_ram[3383] = 147;
    exp_41_ram[3384] = 3;
    exp_41_ram[3385] = 131;
    exp_41_ram[3386] = 51;
    exp_41_ram[3387] = 19;
    exp_41_ram[3388] = 51;
    exp_41_ram[3389] = 179;
    exp_41_ram[3390] = 179;
    exp_41_ram[3391] = 147;
    exp_41_ram[3392] = 35;
    exp_41_ram[3393] = 35;
    exp_41_ram[3394] = 183;
    exp_41_ram[3395] = 147;
    exp_41_ram[3396] = 147;
    exp_41_ram[3397] = 131;
    exp_41_ram[3398] = 3;
    exp_41_ram[3399] = 19;
    exp_41_ram[3400] = 239;
    exp_41_ram[3401] = 3;
    exp_41_ram[3402] = 131;
    exp_41_ram[3403] = 3;
    exp_41_ram[3404] = 3;
    exp_41_ram[3405] = 131;
    exp_41_ram[3406] = 3;
    exp_41_ram[3407] = 131;
    exp_41_ram[3408] = 3;
    exp_41_ram[3409] = 131;
    exp_41_ram[3410] = 35;
    exp_41_ram[3411] = 35;
    exp_41_ram[3412] = 35;
    exp_41_ram[3413] = 35;
    exp_41_ram[3414] = 35;
    exp_41_ram[3415] = 35;
    exp_41_ram[3416] = 35;
    exp_41_ram[3417] = 35;
    exp_41_ram[3418] = 35;
    exp_41_ram[3419] = 3;
    exp_41_ram[3420] = 131;
    exp_41_ram[3421] = 239;
    exp_41_ram[3422] = 19;
    exp_41_ram[3423] = 183;
    exp_41_ram[3424] = 147;
    exp_41_ram[3425] = 35;
    exp_41_ram[3426] = 183;
    exp_41_ram[3427] = 147;
    exp_41_ram[3428] = 19;
    exp_41_ram[3429] = 131;
    exp_41_ram[3430] = 3;
    exp_41_ram[3431] = 131;
    exp_41_ram[3432] = 3;
    exp_41_ram[3433] = 131;
    exp_41_ram[3434] = 19;
    exp_41_ram[3435] = 103;
    exp_41_ram[3436] = 19;
    exp_41_ram[3437] = 35;
    exp_41_ram[3438] = 35;
    exp_41_ram[3439] = 19;
    exp_41_ram[3440] = 35;
    exp_41_ram[3441] = 35;
    exp_41_ram[3442] = 3;
    exp_41_ram[3443] = 239;
    exp_41_ram[3444] = 147;
    exp_41_ram[3445] = 163;
    exp_41_ram[3446] = 131;
    exp_41_ram[3447] = 19;
    exp_41_ram[3448] = 147;
    exp_41_ram[3449] = 99;
    exp_41_ram[3450] = 3;
    exp_41_ram[3451] = 147;
    exp_41_ram[3452] = 147;
    exp_41_ram[3453] = 179;
    exp_41_ram[3454] = 147;
    exp_41_ram[3455] = 35;
    exp_41_ram[3456] = 3;
    exp_41_ram[3457] = 131;
    exp_41_ram[3458] = 179;
    exp_41_ram[3459] = 147;
    exp_41_ram[3460] = 35;
    exp_41_ram[3461] = 111;
    exp_41_ram[3462] = 19;
    exp_41_ram[3463] = 131;
    exp_41_ram[3464] = 19;
    exp_41_ram[3465] = 131;
    exp_41_ram[3466] = 3;
    exp_41_ram[3467] = 19;
    exp_41_ram[3468] = 103;
    exp_41_ram[3469] = 19;
    exp_41_ram[3470] = 35;
    exp_41_ram[3471] = 35;
    exp_41_ram[3472] = 19;
    exp_41_ram[3473] = 183;
    exp_41_ram[3474] = 131;
    exp_41_ram[3475] = 19;
    exp_41_ram[3476] = 239;
    exp_41_ram[3477] = 147;
    exp_41_ram[3478] = 19;
    exp_41_ram[3479] = 131;
    exp_41_ram[3480] = 3;
    exp_41_ram[3481] = 19;
    exp_41_ram[3482] = 103;
    exp_41_ram[3483] = 19;
    exp_41_ram[3484] = 35;
    exp_41_ram[3485] = 35;
    exp_41_ram[3486] = 35;
    exp_41_ram[3487] = 35;
    exp_41_ram[3488] = 19;
    exp_41_ram[3489] = 35;
    exp_41_ram[3490] = 239;
    exp_41_ram[3491] = 35;
    exp_41_ram[3492] = 35;
    exp_41_ram[3493] = 19;
    exp_41_ram[3494] = 239;
    exp_41_ram[3495] = 19;
    exp_41_ram[3496] = 147;
    exp_41_ram[3497] = 3;
    exp_41_ram[3498] = 131;
    exp_41_ram[3499] = 51;
    exp_41_ram[3500] = 19;
    exp_41_ram[3501] = 51;
    exp_41_ram[3502] = 179;
    exp_41_ram[3503] = 179;
    exp_41_ram[3504] = 147;
    exp_41_ram[3505] = 131;
    exp_41_ram[3506] = 19;
    exp_41_ram[3507] = 147;
    exp_41_ram[3508] = 19;
    exp_41_ram[3509] = 147;
    exp_41_ram[3510] = 227;
    exp_41_ram[3511] = 19;
    exp_41_ram[3512] = 147;
    exp_41_ram[3513] = 99;
    exp_41_ram[3514] = 147;
    exp_41_ram[3515] = 147;
    exp_41_ram[3516] = 227;
    exp_41_ram[3517] = 19;
    exp_41_ram[3518] = 19;
    exp_41_ram[3519] = 131;
    exp_41_ram[3520] = 3;
    exp_41_ram[3521] = 3;
    exp_41_ram[3522] = 131;
    exp_41_ram[3523] = 19;
    exp_41_ram[3524] = 103;
    exp_41_ram[3525] = 19;
    exp_41_ram[3526] = 35;
    exp_41_ram[3527] = 35;
    exp_41_ram[3528] = 19;
    exp_41_ram[3529] = 183;
    exp_41_ram[3530] = 19;
    exp_41_ram[3531] = 239;
    exp_41_ram[3532] = 19;
    exp_41_ram[3533] = 131;
    exp_41_ram[3534] = 3;
    exp_41_ram[3535] = 19;
    exp_41_ram[3536] = 103;
    exp_41_ram[3537] = 19;
    exp_41_ram[3538] = 35;
    exp_41_ram[3539] = 35;
    exp_41_ram[3540] = 19;
    exp_41_ram[3541] = 183;
    exp_41_ram[3542] = 19;
    exp_41_ram[3543] = 239;
    exp_41_ram[3544] = 147;
    exp_41_ram[3545] = 35;
    exp_41_ram[3546] = 35;
    exp_41_ram[3547] = 111;
    exp_41_ram[3548] = 131;
    exp_41_ram[3549] = 183;
    exp_41_ram[3550] = 19;
    exp_41_ram[3551] = 239;
    exp_41_ram[3552] = 111;
    exp_41_ram[3553] = 131;
    exp_41_ram[3554] = 147;
    exp_41_ram[3555] = 35;
    exp_41_ram[3556] = 183;
    exp_41_ram[3557] = 131;
    exp_41_ram[3558] = 147;
    exp_41_ram[3559] = 3;
    exp_41_ram[3560] = 239;
    exp_41_ram[3561] = 183;
    exp_41_ram[3562] = 3;
    exp_41_ram[3563] = 147;
    exp_41_ram[3564] = 179;
    exp_41_ram[3565] = 19;
    exp_41_ram[3566] = 239;
    exp_41_ram[3567] = 3;
    exp_41_ram[3568] = 147;
    exp_41_ram[3569] = 227;
    exp_41_ram[3570] = 111;
    exp_41_ram[3571] = 131;
    exp_41_ram[3572] = 147;
    exp_41_ram[3573] = 35;
    exp_41_ram[3574] = 183;
    exp_41_ram[3575] = 131;
    exp_41_ram[3576] = 147;
    exp_41_ram[3577] = 3;
    exp_41_ram[3578] = 239;
    exp_41_ram[3579] = 183;
    exp_41_ram[3580] = 3;
    exp_41_ram[3581] = 147;
    exp_41_ram[3582] = 179;
    exp_41_ram[3583] = 19;
    exp_41_ram[3584] = 239;
    exp_41_ram[3585] = 3;
    exp_41_ram[3586] = 147;
    exp_41_ram[3587] = 227;
    exp_41_ram[3588] = 131;
    exp_41_ram[3589] = 147;
    exp_41_ram[3590] = 35;
    exp_41_ram[3591] = 3;
    exp_41_ram[3592] = 147;
    exp_41_ram[3593] = 227;
    exp_41_ram[3594] = 183;
    exp_41_ram[3595] = 131;
    exp_41_ram[3596] = 147;
    exp_41_ram[3597] = 19;
    exp_41_ram[3598] = 239;
    exp_41_ram[3599] = 19;
    exp_41_ram[3600] = 131;
    exp_41_ram[3601] = 3;
    exp_41_ram[3602] = 19;
    exp_41_ram[3603] = 103;
    exp_41_ram[3604] = 19;
    exp_41_ram[3605] = 35;
    exp_41_ram[3606] = 35;
    exp_41_ram[3607] = 35;
    exp_41_ram[3608] = 35;
    exp_41_ram[3609] = 35;
    exp_41_ram[3610] = 35;
    exp_41_ram[3611] = 35;
    exp_41_ram[3612] = 35;
    exp_41_ram[3613] = 35;
    exp_41_ram[3614] = 35;
    exp_41_ram[3615] = 35;
    exp_41_ram[3616] = 35;
    exp_41_ram[3617] = 19;
    exp_41_ram[3618] = 147;
    exp_41_ram[3619] = 35;
    exp_41_ram[3620] = 19;
    exp_41_ram[3621] = 147;
    exp_41_ram[3622] = 35;
    exp_41_ram[3623] = 35;
    exp_41_ram[3624] = 239;
    exp_41_ram[3625] = 35;
    exp_41_ram[3626] = 35;
    exp_41_ram[3627] = 35;
    exp_41_ram[3628] = 111;
    exp_41_ram[3629] = 3;
    exp_41_ram[3630] = 183;
    exp_41_ram[3631] = 147;
    exp_41_ram[3632] = 179;
    exp_41_ram[3633] = 35;
    exp_41_ram[3634] = 3;
    exp_41_ram[3635] = 183;
    exp_41_ram[3636] = 147;
    exp_41_ram[3637] = 179;
    exp_41_ram[3638] = 35;
    exp_41_ram[3639] = 3;
    exp_41_ram[3640] = 183;
    exp_41_ram[3641] = 147;
    exp_41_ram[3642] = 179;
    exp_41_ram[3643] = 35;
    exp_41_ram[3644] = 3;
    exp_41_ram[3645] = 183;
    exp_41_ram[3646] = 147;
    exp_41_ram[3647] = 179;
    exp_41_ram[3648] = 35;
    exp_41_ram[3649] = 131;
    exp_41_ram[3650] = 147;
    exp_41_ram[3651] = 35;
    exp_41_ram[3652] = 239;
    exp_41_ram[3653] = 19;
    exp_41_ram[3654] = 147;
    exp_41_ram[3655] = 3;
    exp_41_ram[3656] = 131;
    exp_41_ram[3657] = 51;
    exp_41_ram[3658] = 19;
    exp_41_ram[3659] = 51;
    exp_41_ram[3660] = 179;
    exp_41_ram[3661] = 179;
    exp_41_ram[3662] = 147;
    exp_41_ram[3663] = 183;
    exp_41_ram[3664] = 131;
    exp_41_ram[3665] = 35;
    exp_41_ram[3666] = 35;
    exp_41_ram[3667] = 3;
    exp_41_ram[3668] = 131;
    exp_41_ram[3669] = 19;
    exp_41_ram[3670] = 147;
    exp_41_ram[3671] = 227;
    exp_41_ram[3672] = 19;
    exp_41_ram[3673] = 147;
    exp_41_ram[3674] = 99;
    exp_41_ram[3675] = 147;
    exp_41_ram[3676] = 147;
    exp_41_ram[3677] = 227;
    exp_41_ram[3678] = 131;
    exp_41_ram[3679] = 183;
    exp_41_ram[3680] = 19;
    exp_41_ram[3681] = 239;
    exp_41_ram[3682] = 239;
    exp_41_ram[3683] = 35;
    exp_41_ram[3684] = 35;
    exp_41_ram[3685] = 35;
    exp_41_ram[3686] = 111;
    exp_41_ram[3687] = 3;
    exp_41_ram[3688] = 131;
    exp_41_ram[3689] = 183;
    exp_41_ram[3690] = 147;
    exp_41_ram[3691] = 51;
    exp_41_ram[3692] = 147;
    exp_41_ram[3693] = 179;
    exp_41_ram[3694] = 51;
    exp_41_ram[3695] = 183;
    exp_41_ram[3696] = 147;
    exp_41_ram[3697] = 179;
    exp_41_ram[3698] = 179;
    exp_41_ram[3699] = 19;
    exp_41_ram[3700] = 179;
    exp_41_ram[3701] = 147;
    exp_41_ram[3702] = 35;
    exp_41_ram[3703] = 35;
    exp_41_ram[3704] = 3;
    exp_41_ram[3705] = 131;
    exp_41_ram[3706] = 183;
    exp_41_ram[3707] = 147;
    exp_41_ram[3708] = 51;
    exp_41_ram[3709] = 147;
    exp_41_ram[3710] = 179;
    exp_41_ram[3711] = 51;
    exp_41_ram[3712] = 183;
    exp_41_ram[3713] = 147;
    exp_41_ram[3714] = 179;
    exp_41_ram[3715] = 179;
    exp_41_ram[3716] = 19;
    exp_41_ram[3717] = 179;
    exp_41_ram[3718] = 147;
    exp_41_ram[3719] = 35;
    exp_41_ram[3720] = 35;
    exp_41_ram[3721] = 3;
    exp_41_ram[3722] = 131;
    exp_41_ram[3723] = 183;
    exp_41_ram[3724] = 147;
    exp_41_ram[3725] = 51;
    exp_41_ram[3726] = 147;
    exp_41_ram[3727] = 179;
    exp_41_ram[3728] = 51;
    exp_41_ram[3729] = 183;
    exp_41_ram[3730] = 147;
    exp_41_ram[3731] = 179;
    exp_41_ram[3732] = 179;
    exp_41_ram[3733] = 19;
    exp_41_ram[3734] = 179;
    exp_41_ram[3735] = 147;
    exp_41_ram[3736] = 35;
    exp_41_ram[3737] = 35;
    exp_41_ram[3738] = 3;
    exp_41_ram[3739] = 131;
    exp_41_ram[3740] = 183;
    exp_41_ram[3741] = 147;
    exp_41_ram[3742] = 51;
    exp_41_ram[3743] = 147;
    exp_41_ram[3744] = 179;
    exp_41_ram[3745] = 51;
    exp_41_ram[3746] = 183;
    exp_41_ram[3747] = 147;
    exp_41_ram[3748] = 179;
    exp_41_ram[3749] = 179;
    exp_41_ram[3750] = 19;
    exp_41_ram[3751] = 179;
    exp_41_ram[3752] = 147;
    exp_41_ram[3753] = 35;
    exp_41_ram[3754] = 35;
    exp_41_ram[3755] = 131;
    exp_41_ram[3756] = 147;
    exp_41_ram[3757] = 35;
    exp_41_ram[3758] = 239;
    exp_41_ram[3759] = 19;
    exp_41_ram[3760] = 147;
    exp_41_ram[3761] = 3;
    exp_41_ram[3762] = 131;
    exp_41_ram[3763] = 51;
    exp_41_ram[3764] = 19;
    exp_41_ram[3765] = 51;
    exp_41_ram[3766] = 179;
    exp_41_ram[3767] = 179;
    exp_41_ram[3768] = 147;
    exp_41_ram[3769] = 183;
    exp_41_ram[3770] = 131;
    exp_41_ram[3771] = 35;
    exp_41_ram[3772] = 35;
    exp_41_ram[3773] = 3;
    exp_41_ram[3774] = 131;
    exp_41_ram[3775] = 19;
    exp_41_ram[3776] = 147;
    exp_41_ram[3777] = 227;
    exp_41_ram[3778] = 19;
    exp_41_ram[3779] = 147;
    exp_41_ram[3780] = 99;
    exp_41_ram[3781] = 147;
    exp_41_ram[3782] = 147;
    exp_41_ram[3783] = 227;
    exp_41_ram[3784] = 131;
    exp_41_ram[3785] = 183;
    exp_41_ram[3786] = 19;
    exp_41_ram[3787] = 239;
    exp_41_ram[3788] = 239;
    exp_41_ram[3789] = 35;
    exp_41_ram[3790] = 35;
    exp_41_ram[3791] = 35;
    exp_41_ram[3792] = 111;
    exp_41_ram[3793] = 3;
    exp_41_ram[3794] = 183;
    exp_41_ram[3795] = 147;
    exp_41_ram[3796] = 179;
    exp_41_ram[3797] = 35;
    exp_41_ram[3798] = 3;
    exp_41_ram[3799] = 183;
    exp_41_ram[3800] = 147;
    exp_41_ram[3801] = 179;
    exp_41_ram[3802] = 35;
    exp_41_ram[3803] = 3;
    exp_41_ram[3804] = 183;
    exp_41_ram[3805] = 147;
    exp_41_ram[3806] = 179;
    exp_41_ram[3807] = 35;
    exp_41_ram[3808] = 3;
    exp_41_ram[3809] = 183;
    exp_41_ram[3810] = 147;
    exp_41_ram[3811] = 179;
    exp_41_ram[3812] = 35;
    exp_41_ram[3813] = 131;
    exp_41_ram[3814] = 147;
    exp_41_ram[3815] = 35;
    exp_41_ram[3816] = 239;
    exp_41_ram[3817] = 19;
    exp_41_ram[3818] = 147;
    exp_41_ram[3819] = 3;
    exp_41_ram[3820] = 131;
    exp_41_ram[3821] = 51;
    exp_41_ram[3822] = 19;
    exp_41_ram[3823] = 51;
    exp_41_ram[3824] = 179;
    exp_41_ram[3825] = 179;
    exp_41_ram[3826] = 147;
    exp_41_ram[3827] = 183;
    exp_41_ram[3828] = 131;
    exp_41_ram[3829] = 35;
    exp_41_ram[3830] = 35;
    exp_41_ram[3831] = 3;
    exp_41_ram[3832] = 131;
    exp_41_ram[3833] = 19;
    exp_41_ram[3834] = 147;
    exp_41_ram[3835] = 227;
    exp_41_ram[3836] = 19;
    exp_41_ram[3837] = 147;
    exp_41_ram[3838] = 99;
    exp_41_ram[3839] = 147;
    exp_41_ram[3840] = 147;
    exp_41_ram[3841] = 227;
    exp_41_ram[3842] = 131;
    exp_41_ram[3843] = 183;
    exp_41_ram[3844] = 19;
    exp_41_ram[3845] = 239;
    exp_41_ram[3846] = 239;
    exp_41_ram[3847] = 35;
    exp_41_ram[3848] = 35;
    exp_41_ram[3849] = 35;
    exp_41_ram[3850] = 111;
    exp_41_ram[3851] = 3;
    exp_41_ram[3852] = 131;
    exp_41_ram[3853] = 55;
    exp_41_ram[3854] = 19;
    exp_41_ram[3855] = 147;
    exp_41_ram[3856] = 19;
    exp_41_ram[3857] = 147;
    exp_41_ram[3858] = 239;
    exp_41_ram[3859] = 19;
    exp_41_ram[3860] = 147;
    exp_41_ram[3861] = 35;
    exp_41_ram[3862] = 35;
    exp_41_ram[3863] = 3;
    exp_41_ram[3864] = 131;
    exp_41_ram[3865] = 55;
    exp_41_ram[3866] = 19;
    exp_41_ram[3867] = 147;
    exp_41_ram[3868] = 19;
    exp_41_ram[3869] = 147;
    exp_41_ram[3870] = 239;
    exp_41_ram[3871] = 19;
    exp_41_ram[3872] = 147;
    exp_41_ram[3873] = 35;
    exp_41_ram[3874] = 35;
    exp_41_ram[3875] = 3;
    exp_41_ram[3876] = 131;
    exp_41_ram[3877] = 55;
    exp_41_ram[3878] = 19;
    exp_41_ram[3879] = 147;
    exp_41_ram[3880] = 19;
    exp_41_ram[3881] = 147;
    exp_41_ram[3882] = 239;
    exp_41_ram[3883] = 19;
    exp_41_ram[3884] = 147;
    exp_41_ram[3885] = 35;
    exp_41_ram[3886] = 35;
    exp_41_ram[3887] = 3;
    exp_41_ram[3888] = 131;
    exp_41_ram[3889] = 55;
    exp_41_ram[3890] = 19;
    exp_41_ram[3891] = 147;
    exp_41_ram[3892] = 19;
    exp_41_ram[3893] = 147;
    exp_41_ram[3894] = 239;
    exp_41_ram[3895] = 19;
    exp_41_ram[3896] = 147;
    exp_41_ram[3897] = 35;
    exp_41_ram[3898] = 35;
    exp_41_ram[3899] = 131;
    exp_41_ram[3900] = 147;
    exp_41_ram[3901] = 35;
    exp_41_ram[3902] = 239;
    exp_41_ram[3903] = 19;
    exp_41_ram[3904] = 147;
    exp_41_ram[3905] = 3;
    exp_41_ram[3906] = 131;
    exp_41_ram[3907] = 51;
    exp_41_ram[3908] = 19;
    exp_41_ram[3909] = 51;
    exp_41_ram[3910] = 179;
    exp_41_ram[3911] = 179;
    exp_41_ram[3912] = 147;
    exp_41_ram[3913] = 183;
    exp_41_ram[3914] = 131;
    exp_41_ram[3915] = 19;
    exp_41_ram[3916] = 147;
    exp_41_ram[3917] = 19;
    exp_41_ram[3918] = 147;
    exp_41_ram[3919] = 227;
    exp_41_ram[3920] = 19;
    exp_41_ram[3921] = 147;
    exp_41_ram[3922] = 99;
    exp_41_ram[3923] = 147;
    exp_41_ram[3924] = 147;
    exp_41_ram[3925] = 227;
    exp_41_ram[3926] = 131;
    exp_41_ram[3927] = 183;
    exp_41_ram[3928] = 19;
    exp_41_ram[3929] = 239;
    exp_41_ram[3930] = 19;
    exp_41_ram[3931] = 131;
    exp_41_ram[3932] = 3;
    exp_41_ram[3933] = 3;
    exp_41_ram[3934] = 131;
    exp_41_ram[3935] = 3;
    exp_41_ram[3936] = 131;
    exp_41_ram[3937] = 3;
    exp_41_ram[3938] = 131;
    exp_41_ram[3939] = 3;
    exp_41_ram[3940] = 131;
    exp_41_ram[3941] = 3;
    exp_41_ram[3942] = 131;
    exp_41_ram[3943] = 19;
    exp_41_ram[3944] = 103;
    exp_41_ram[3945] = 19;
    exp_41_ram[3946] = 35;
    exp_41_ram[3947] = 35;
    exp_41_ram[3948] = 35;
    exp_41_ram[3949] = 35;
    exp_41_ram[3950] = 35;
    exp_41_ram[3951] = 35;
    exp_41_ram[3952] = 19;
    exp_41_ram[3953] = 183;
    exp_41_ram[3954] = 19;
    exp_41_ram[3955] = 239;
    exp_41_ram[3956] = 239;
    exp_41_ram[3957] = 147;
    exp_41_ram[3958] = 147;
    exp_41_ram[3959] = 35;
    exp_41_ram[3960] = 183;
    exp_41_ram[3961] = 19;
    exp_41_ram[3962] = 239;
    exp_41_ram[3963] = 239;
    exp_41_ram[3964] = 147;
    exp_41_ram[3965] = 147;
    exp_41_ram[3966] = 35;
    exp_41_ram[3967] = 183;
    exp_41_ram[3968] = 19;
    exp_41_ram[3969] = 239;
    exp_41_ram[3970] = 239;
    exp_41_ram[3971] = 147;
    exp_41_ram[3972] = 35;
    exp_41_ram[3973] = 183;
    exp_41_ram[3974] = 19;
    exp_41_ram[3975] = 239;
    exp_41_ram[3976] = 239;
    exp_41_ram[3977] = 147;
    exp_41_ram[3978] = 35;
    exp_41_ram[3979] = 183;
    exp_41_ram[3980] = 19;
    exp_41_ram[3981] = 239;
    exp_41_ram[3982] = 239;
    exp_41_ram[3983] = 147;
    exp_41_ram[3984] = 35;
    exp_41_ram[3985] = 147;
    exp_41_ram[3986] = 35;
    exp_41_ram[3987] = 147;
    exp_41_ram[3988] = 35;
    exp_41_ram[3989] = 147;
    exp_41_ram[3990] = 19;
    exp_41_ram[3991] = 239;
    exp_41_ram[3992] = 19;
    exp_41_ram[3993] = 147;
    exp_41_ram[3994] = 35;
    exp_41_ram[3995] = 35;
    exp_41_ram[3996] = 3;
    exp_41_ram[3997] = 131;
    exp_41_ram[3998] = 19;
    exp_41_ram[3999] = 147;
    exp_41_ram[4000] = 239;
    exp_41_ram[4001] = 239;
    exp_41_ram[4002] = 35;
    exp_41_ram[4003] = 35;
    exp_41_ram[4004] = 35;
    exp_41_ram[4005] = 111;
    exp_41_ram[4006] = 19;
    exp_41_ram[4007] = 239;
    exp_41_ram[4008] = 19;
    exp_41_ram[4009] = 147;
    exp_41_ram[4010] = 3;
    exp_41_ram[4011] = 131;
    exp_41_ram[4012] = 19;
    exp_41_ram[4013] = 147;
    exp_41_ram[4014] = 239;
    exp_41_ram[4015] = 19;
    exp_41_ram[4016] = 147;
    exp_41_ram[4017] = 183;
    exp_41_ram[4018] = 131;
    exp_41_ram[4019] = 19;
    exp_41_ram[4020] = 239;
    exp_41_ram[4021] = 19;
    exp_41_ram[4022] = 147;
    exp_41_ram[4023] = 19;
    exp_41_ram[4024] = 147;
    exp_41_ram[4025] = 19;
    exp_41_ram[4026] = 147;
    exp_41_ram[4027] = 239;
    exp_41_ram[4028] = 147;
    exp_41_ram[4029] = 227;
    exp_41_ram[4030] = 183;
    exp_41_ram[4031] = 131;
    exp_41_ram[4032] = 19;
    exp_41_ram[4033] = 147;
    exp_41_ram[4034] = 3;
    exp_41_ram[4035] = 131;
    exp_41_ram[4036] = 51;
    exp_41_ram[4037] = 147;
    exp_41_ram[4038] = 179;
    exp_41_ram[4039] = 179;
    exp_41_ram[4040] = 179;
    exp_41_ram[4041] = 147;
    exp_41_ram[4042] = 35;
    exp_41_ram[4043] = 35;
    exp_41_ram[4044] = 19;
    exp_41_ram[4045] = 239;
    exp_41_ram[4046] = 19;
    exp_41_ram[4047] = 147;
    exp_41_ram[4048] = 35;
    exp_41_ram[4049] = 35;
    exp_41_ram[4050] = 147;
    exp_41_ram[4051] = 19;
    exp_41_ram[4052] = 239;
    exp_41_ram[4053] = 147;
    exp_41_ram[4054] = 19;
    exp_41_ram[4055] = 239;
    exp_41_ram[4056] = 131;
    exp_41_ram[4057] = 147;
    exp_41_ram[4058] = 35;
    exp_41_ram[4059] = 3;
    exp_41_ram[4060] = 147;
    exp_41_ram[4061] = 227;
    exp_41_ram[4062] = 19;
    exp_41_ram[4063] = 19;
    exp_41_ram[4064] = 131;
    exp_41_ram[4065] = 3;
    exp_41_ram[4066] = 3;
    exp_41_ram[4067] = 131;
    exp_41_ram[4068] = 3;
    exp_41_ram[4069] = 131;
    exp_41_ram[4070] = 19;
    exp_41_ram[4071] = 103;
    exp_41_ram[4072] = 19;
    exp_41_ram[4073] = 35;
    exp_41_ram[4074] = 35;
    exp_41_ram[4075] = 19;
    exp_41_ram[4076] = 183;
    exp_41_ram[4077] = 19;
    exp_41_ram[4078] = 239;
    exp_41_ram[4079] = 183;
    exp_41_ram[4080] = 19;
    exp_41_ram[4081] = 239;
    exp_41_ram[4082] = 183;
    exp_41_ram[4083] = 19;
    exp_41_ram[4084] = 239;
    exp_41_ram[4085] = 183;
    exp_41_ram[4086] = 19;
    exp_41_ram[4087] = 239;
    exp_41_ram[4088] = 183;
    exp_41_ram[4089] = 19;
    exp_41_ram[4090] = 239;
    exp_41_ram[4091] = 239;
    exp_41_ram[4092] = 147;
    exp_41_ram[4093] = 163;
    exp_41_ram[4094] = 131;
    exp_41_ram[4095] = 19;
    exp_41_ram[4096] = 99;
    exp_41_ram[4097] = 19;
    exp_41_ram[4098] = 227;
    exp_41_ram[4099] = 19;
    exp_41_ram[4100] = 99;
    exp_41_ram[4101] = 19;
    exp_41_ram[4102] = 227;
    exp_41_ram[4103] = 19;
    exp_41_ram[4104] = 99;
    exp_41_ram[4105] = 19;
    exp_41_ram[4106] = 99;
    exp_41_ram[4107] = 111;
    exp_41_ram[4108] = 239;
    exp_41_ram[4109] = 111;
    exp_41_ram[4110] = 239;
    exp_41_ram[4111] = 111;
    exp_41_ram[4112] = 239;
    exp_41_ram[4113] = 111;
    exp_41_ram[4114] = 239;
    exp_41_ram[4115] = 19;
    exp_41_ram[4116] = 111;
    exp_41_ram[4117] = 19;
    exp_41_ram[4118] = 147;
    exp_41_ram[4119] = 51;
    exp_41_ram[4120] = 19;
    exp_41_ram[4121] = 179;
    exp_41_ram[4122] = 99;
    exp_41_ram[4123] = 99;
    exp_41_ram[4124] = 19;
    exp_41_ram[4125] = 179;
    exp_41_ram[4126] = 19;
    exp_41_ram[4127] = 103;
    exp_41_ram[4128] = 227;
    exp_41_ram[4129] = 19;
    exp_41_ram[4130] = 179;
    exp_41_ram[4131] = 111;
    exp_41_ram[4132] = 128;
    exp_41_ram[4133] = 8;
    exp_41_ram[4134] = 12;
    exp_41_ram[4135] = 16;
    exp_41_ram[4136] = 40;
    exp_41_ram[4137] = 112;
    exp_41_ram[4138] = 112;
    exp_41_ram[4139] = 76;
    exp_41_ram[4140] = 112;
    exp_41_ram[4141] = 112;
    exp_41_ram[4142] = 112;
    exp_41_ram[4143] = 112;
    exp_41_ram[4144] = 112;
    exp_41_ram[4145] = 112;
    exp_41_ram[4146] = 112;
    exp_41_ram[4147] = 4;
    exp_41_ram[4148] = 112;
    exp_41_ram[4149] = 224;
    exp_41_ram[4150] = 112;
    exp_41_ram[4151] = 112;
    exp_41_ram[4152] = 188;
    exp_41_ram[4153] = 20;
    exp_41_ram[4154] = 172;
    exp_41_ram[4155] = 116;
    exp_41_ram[4156] = 172;
    exp_41_ram[4157] = 208;
    exp_41_ram[4158] = 172;
    exp_41_ram[4159] = 172;
    exp_41_ram[4160] = 172;
    exp_41_ram[4161] = 172;
    exp_41_ram[4162] = 172;
    exp_41_ram[4163] = 172;
    exp_41_ram[4164] = 172;
    exp_41_ram[4165] = 88;
    exp_41_ram[4166] = 172;
    exp_41_ram[4167] = 172;
    exp_41_ram[4168] = 172;
    exp_41_ram[4169] = 172;
    exp_41_ram[4170] = 172;
    exp_41_ram[4171] = 144;
    exp_41_ram[4172] = 212;
    exp_41_ram[4173] = 8;
    exp_41_ram[4174] = 8;
    exp_41_ram[4175] = 8;
    exp_41_ram[4176] = 8;
    exp_41_ram[4177] = 8;
    exp_41_ram[4178] = 8;
    exp_41_ram[4179] = 8;
    exp_41_ram[4180] = 8;
    exp_41_ram[4181] = 8;
    exp_41_ram[4182] = 8;
    exp_41_ram[4183] = 8;
    exp_41_ram[4184] = 8;
    exp_41_ram[4185] = 8;
    exp_41_ram[4186] = 8;
    exp_41_ram[4187] = 8;
    exp_41_ram[4188] = 8;
    exp_41_ram[4189] = 8;
    exp_41_ram[4190] = 8;
    exp_41_ram[4191] = 8;
    exp_41_ram[4192] = 8;
    exp_41_ram[4193] = 8;
    exp_41_ram[4194] = 8;
    exp_41_ram[4195] = 8;
    exp_41_ram[4196] = 8;
    exp_41_ram[4197] = 8;
    exp_41_ram[4198] = 8;
    exp_41_ram[4199] = 8;
    exp_41_ram[4200] = 8;
    exp_41_ram[4201] = 8;
    exp_41_ram[4202] = 8;
    exp_41_ram[4203] = 8;
    exp_41_ram[4204] = 8;
    exp_41_ram[4205] = 8;
    exp_41_ram[4206] = 8;
    exp_41_ram[4207] = 8;
    exp_41_ram[4208] = 8;
    exp_41_ram[4209] = 8;
    exp_41_ram[4210] = 8;
    exp_41_ram[4211] = 8;
    exp_41_ram[4212] = 8;
    exp_41_ram[4213] = 8;
    exp_41_ram[4214] = 8;
    exp_41_ram[4215] = 8;
    exp_41_ram[4216] = 8;
    exp_41_ram[4217] = 8;
    exp_41_ram[4218] = 8;
    exp_41_ram[4219] = 8;
    exp_41_ram[4220] = 8;
    exp_41_ram[4221] = 8;
    exp_41_ram[4222] = 8;
    exp_41_ram[4223] = 236;
    exp_41_ram[4224] = 8;
    exp_41_ram[4225] = 8;
    exp_41_ram[4226] = 8;
    exp_41_ram[4227] = 8;
    exp_41_ram[4228] = 8;
    exp_41_ram[4229] = 8;
    exp_41_ram[4230] = 8;
    exp_41_ram[4231] = 8;
    exp_41_ram[4232] = 8;
    exp_41_ram[4233] = 236;
    exp_41_ram[4234] = 56;
    exp_41_ram[4235] = 236;
    exp_41_ram[4236] = 8;
    exp_41_ram[4237] = 8;
    exp_41_ram[4238] = 8;
    exp_41_ram[4239] = 8;
    exp_41_ram[4240] = 236;
    exp_41_ram[4241] = 8;
    exp_41_ram[4242] = 8;
    exp_41_ram[4243] = 8;
    exp_41_ram[4244] = 8;
    exp_41_ram[4245] = 8;
    exp_41_ram[4246] = 236;
    exp_41_ram[4247] = 104;
    exp_41_ram[4248] = 8;
    exp_41_ram[4249] = 8;
    exp_41_ram[4250] = 20;
    exp_41_ram[4251] = 8;
    exp_41_ram[4252] = 236;
    exp_41_ram[4253] = 8;
    exp_41_ram[4254] = 8;
    exp_41_ram[4255] = 236;
    exp_41_ram[4256] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_39) begin
      exp_41_ram[exp_35] <= exp_37;
    end
  end
  assign exp_41 = exp_41_ram[exp_36];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_67) begin
        exp_41_ram[exp_63] <= exp_65;
    end
  end
  assign exp_69 = exp_41_ram[exp_64];
  assign exp_68 = exp_100;
  assign exp_100 = 1;
  assign exp_64 = exp_99;
  assign exp_99 = exp_16[31:2];
  assign exp_67 = exp_92;
  assign exp_63 = exp_91;
  assign exp_65 = exp_91;
  assign exp_40 = exp_135;
  assign exp_135 = 1;
  assign exp_36 = exp_134;
  assign exp_134 = exp_18[31:2];
  assign exp_39 = exp_109;
  assign exp_109 = exp_107 & exp_108;
  assign exp_107 = exp_22 & exp_23;
  assign exp_108 = exp_24[0:0];
  assign exp_35 = exp_105;
  assign exp_105 = exp_18[31:2];
  assign exp_37 = exp_106;
  assign exp_106 = exp_19[7:0];
  assign exp_126 = 1;
  assign exp_149 = exp_187;

  reg [31:0] exp_187_reg;
  always@(*) begin
    case (exp_185)
      0:exp_187_reg <= exp_165;
      1:exp_187_reg <= exp_175;
      default:exp_187_reg <= exp_186;
    endcase
  end
  assign exp_187 = exp_187_reg;
  assign exp_185 = exp_147[2:2];
  assign exp_147 = exp_9;
  assign exp_186 = 0;

      reg [31:0] exp_165_reg = 0;
      always@(posedge clk) begin
        if (exp_164) begin
          exp_165_reg <= exp_172;
        end
      end
      assign exp_165 = exp_165_reg;
    
  reg [31:0] exp_172_reg;
  always@(*) begin
    case (exp_167)
      0:exp_172_reg <= exp_169;
      1:exp_172_reg <= exp_170;
      default:exp_172_reg <= exp_171;
    endcase
  end
  assign exp_172 = exp_172_reg;
  assign exp_167 = exp_165 == exp_166;
  assign exp_166 = 4294967295;
  assign exp_171 = 0;
  assign exp_169 = exp_165 + exp_168;
  assign exp_168 = 1;
  assign exp_170 = 0;
  assign exp_164 = 1;

      reg [31:0] exp_175_reg = 0;
      always@(posedge clk) begin
        if (exp_174) begin
          exp_175_reg <= exp_182;
        end
      end
      assign exp_175 = exp_175_reg;
    
  reg [31:0] exp_182_reg;
  always@(*) begin
    case (exp_177)
      0:exp_182_reg <= exp_179;
      1:exp_182_reg <= exp_180;
      default:exp_182_reg <= exp_181;
    endcase
  end
  assign exp_182 = exp_182_reg;
  assign exp_177 = exp_175 == exp_176;
  assign exp_176 = 4294967295;
  assign exp_181 = 0;
  assign exp_179 = exp_175 + exp_178;
  assign exp_178 = 1;
  assign exp_180 = 0;
  assign exp_174 = exp_167 & exp_173;
  assign exp_173 = 1;
  assign exp_190 = exp_274;
  assign exp_274 = exp_271;

      reg [7:0] exp_271_reg = 0;
      always@(posedge clk) begin
        if (exp_270) begin
          exp_271_reg <= exp_273;
        end
      end
      assign exp_271 = exp_271_reg;
      assign exp_273 = {exp_212, exp_272};  assign exp_272 = exp_271[7:1];
  assign exp_270 = exp_235 & exp_269;
  assign exp_269 = exp_236 == exp_268;
  assign exp_268 = 0;
  assign exp_277 = exp_376;
  assign exp_376 = 0;
  assign exp_379 = exp_396;
  assign exp_396 = 0;
  assign exp_613 = exp_400[15:8];
  assign exp_614 = exp_400[23:16];
  assign exp_615 = exp_400[31:24];
  assign exp_627 = $signed(exp_626);
  assign exp_626 = exp_625 + exp_621;
  assign exp_625 = 0;

  reg [15:0] exp_621_reg;
  always@(*) begin
    case (exp_611)
      0:exp_621_reg <= exp_618;
      1:exp_621_reg <= exp_619;
      default:exp_621_reg <= exp_620;
    endcase
  end
  assign exp_621 = exp_621_reg;
  assign exp_620 = 0;
  assign exp_618 = exp_400[15:0];
  assign exp_619 = exp_400[31:16];
  assign exp_628 = 0;
  assign exp_629 = exp_617;
  assign exp_630 = exp_621;
  assign exp_631 = 0;
  assign exp_632 = 0;

  reg [31:0] exp_991_reg;
  always@(*) begin
    case (exp_781)
      0:exp_991_reg <= exp_987;
      1:exp_991_reg <= exp_989;
      default:exp_991_reg <= exp_990;
    endcase
  end
  assign exp_991 = exp_991_reg;
  assign exp_990 = 0;

  reg [31:0] exp_987_reg;
  always@(*) begin
    case (exp_758)
      0:exp_987_reg <= exp_982;
      1:exp_987_reg <= exp_983;
      default:exp_987_reg <= exp_986;
    endcase
  end
  assign exp_987 = exp_987_reg;
  assign exp_758 = exp_757 & exp_755;
  assign exp_757 = exp_750 == exp_756;
  assign exp_756 = 0;
  assign exp_986 = 0;
  assign exp_982 = exp_981[63:32];

  reg [63:0] exp_981_reg;
  always@(*) begin
    case (exp_978)
      0:exp_981_reg <= exp_977;
      1:exp_981_reg <= exp_979;
      default:exp_981_reg <= exp_980;
    endcase
  end
  assign exp_981 = exp_981_reg;

      reg [0:0] exp_978_reg = 0;
      always@(posedge clk) begin
        if (exp_963) begin
          exp_978_reg <= exp_961;
        end
      end
      assign exp_978 = exp_978_reg;
    
      reg [0:0] exp_961_reg = 0;
      always@(posedge clk) begin
        if (exp_940) begin
          exp_961_reg <= exp_938;
        end
      end
      assign exp_961 = exp_961_reg;
    
      reg [0:0] exp_938_reg = 0;
      always@(posedge clk) begin
        if (exp_920) begin
          exp_938_reg <= exp_935;
        end
      end
      assign exp_938 = exp_938_reg;
      assign exp_935 = exp_933 ^ exp_934;
  assign exp_933 = exp_915 & exp_898;
  assign exp_915 = exp_914 + exp_913;
  assign exp_914 = 0;
  assign exp_913 = exp_911[31:31];

      reg [31:0] exp_911_reg = 0;
      always@(posedge clk) begin
        if (exp_910) begin
          exp_911_reg <= exp_528;
        end
      end
      assign exp_911 = exp_911_reg;
      assign exp_910 = exp_900 == exp_909;
  assign exp_909 = 0;
  assign exp_898 = exp_897 | exp_764;
  assign exp_897 = exp_758 | exp_761;
  assign exp_761 = exp_760 & exp_755;
  assign exp_760 = exp_750 == exp_759;
  assign exp_759 = 1;
  assign exp_764 = exp_763 & exp_755;
  assign exp_763 = exp_750 == exp_762;
  assign exp_762 = 2;
  assign exp_934 = exp_918 & exp_899;
  assign exp_918 = exp_917 + exp_916;
  assign exp_917 = 0;
  assign exp_916 = exp_912[31:31];

      reg [31:0] exp_912_reg = 0;
      always@(posedge clk) begin
        if (exp_910) begin
          exp_912_reg <= exp_529;
        end
      end
      assign exp_912 = exp_912_reg;
      assign exp_899 = exp_758 | exp_761;
  assign exp_920 = exp_900 == exp_919;
  assign exp_919 = 1;
  assign exp_940 = exp_900 == exp_939;
  assign exp_939 = 2;
  assign exp_963 = exp_900 == exp_962;
  assign exp_962 = 3;
  assign exp_980 = 0;

      reg [63:0] exp_977_reg = 0;
      always@(posedge clk) begin
        if (exp_963) begin
          exp_977_reg <= exp_976;
        end
      end
      assign exp_977 = exp_977_reg;
      assign exp_976 = exp_972 + exp_975;
  assign exp_972 = exp_968 + exp_971;
  assign exp_968 = exp_964 + exp_967;
  assign exp_964 = exp_957;

      reg [31:0] exp_957_reg = 0;
      always@(posedge clk) begin
        if (exp_940) begin
          exp_957_reg <= exp_944;
        end
      end
      assign exp_957 = exp_957_reg;
      assign exp_944 = exp_942 * exp_943;
  assign exp_942 = exp_941;
  assign exp_941 = exp_936[15:0];

      reg [31:0] exp_936_reg = 0;
      always@(posedge clk) begin
        if (exp_920) begin
          exp_936_reg <= exp_926;
        end
      end
      assign exp_936 = exp_936_reg;
      assign exp_926 = exp_925 + exp_924;
  assign exp_925 = 0;

  reg [31:0] exp_924_reg;
  always@(*) begin
    case (exp_921)
      0:exp_924_reg <= exp_911;
      1:exp_924_reg <= exp_922;
      default:exp_924_reg <= exp_923;
    endcase
  end
  assign exp_924 = exp_924_reg;
  assign exp_921 = exp_915 & exp_898;
  assign exp_923 = 0;
  assign exp_922 = -exp_911;
  assign exp_943 = exp_937[15:0];

      reg [31:0] exp_937_reg = 0;
      always@(posedge clk) begin
        if (exp_920) begin
          exp_937_reg <= exp_932;
        end
      end
      assign exp_937 = exp_937_reg;
      assign exp_932 = exp_931 + exp_930;
  assign exp_931 = 0;

  reg [31:0] exp_930_reg;
  always@(*) begin
    case (exp_927)
      0:exp_930_reg <= exp_912;
      1:exp_930_reg <= exp_928;
      default:exp_930_reg <= exp_929;
    endcase
  end
  assign exp_930 = exp_930_reg;
  assign exp_927 = exp_918 & exp_899;
  assign exp_929 = 0;
  assign exp_928 = -exp_912;
  assign exp_967 = exp_965 << exp_966;
  assign exp_965 = exp_958;

      reg [31:0] exp_958_reg = 0;
      always@(posedge clk) begin
        if (exp_940) begin
          exp_958_reg <= exp_948;
        end
      end
      assign exp_958 = exp_958_reg;
      assign exp_948 = exp_946 * exp_947;
  assign exp_946 = exp_945;
  assign exp_945 = exp_936[15:0];
  assign exp_947 = exp_937[31:16];
  assign exp_966 = 16;
  assign exp_971 = exp_969 << exp_970;
  assign exp_969 = exp_959;

      reg [31:0] exp_959_reg = 0;
      always@(posedge clk) begin
        if (exp_940) begin
          exp_959_reg <= exp_952;
        end
      end
      assign exp_959 = exp_959_reg;
      assign exp_952 = exp_950 * exp_951;
  assign exp_950 = exp_949;
  assign exp_949 = exp_936[31:16];
  assign exp_951 = exp_937[15:0];
  assign exp_970 = 16;
  assign exp_975 = exp_973 << exp_974;
  assign exp_973 = exp_960;

      reg [31:0] exp_960_reg = 0;
      always@(posedge clk) begin
        if (exp_940) begin
          exp_960_reg <= exp_956;
        end
      end
      assign exp_960 = exp_960_reg;
      assign exp_956 = exp_954 * exp_955;
  assign exp_954 = exp_953;
  assign exp_953 = exp_936[31:16];
  assign exp_955 = exp_937[31:16];
  assign exp_974 = 32;
  assign exp_979 = -exp_977;
  assign exp_983 = exp_981[31:0];

  reg [31:0] exp_989_reg;
  always@(*) begin
    case (exp_782)
      0:exp_989_reg <= exp_892;
      1:exp_989_reg <= exp_893;
      default:exp_989_reg <= exp_988;
    endcase
  end
  assign exp_989 = exp_989_reg;
  assign exp_782 = exp_750[1:1];
  assign exp_988 = 0;

      reg [31:0] exp_892_reg = 0;
      always@(posedge clk) begin
        if (exp_801) begin
          exp_892_reg <= exp_886;
        end
      end
      assign exp_892 = exp_892_reg;
    
  reg [31:0] exp_886_reg;
  always@(*) begin
    case (exp_882)
      0:exp_886_reg <= exp_873;
      1:exp_886_reg <= exp_884;
      default:exp_886_reg <= exp_885;
    endcase
  end
  assign exp_886 = exp_886_reg;
  assign exp_882 = exp_881 & exp_784;
  assign exp_881 = exp_830 == exp_880;

      reg [31:0] exp_830_reg = 0;
      always@(posedge clk) begin
        if (exp_815) begin
          exp_830_reg <= exp_827;
        end
      end
      assign exp_830 = exp_830_reg;
      assign exp_827 = exp_826 + exp_825;
  assign exp_826 = 0;

  reg [31:0] exp_825_reg;
  always@(*) begin
    case (exp_822)
      0:exp_825_reg <= exp_807;
      1:exp_825_reg <= exp_823;
      default:exp_825_reg <= exp_824;
    endcase
  end
  assign exp_825 = exp_825_reg;
  assign exp_822 = exp_813 & exp_784;
  assign exp_813 = exp_812 + exp_811;
  assign exp_812 = 0;
  assign exp_811 = exp_807[31:31];

      reg [31:0] exp_807_reg = 0;
      always@(posedge clk) begin
        if (exp_805) begin
          exp_807_reg <= exp_529;
        end
      end
      assign exp_807 = exp_807_reg;
      assign exp_805 = exp_787 == exp_804;
  assign exp_804 = 0;
  assign exp_784 = ~exp_783;
  assign exp_783 = exp_750[0:0];
  assign exp_824 = 0;
  assign exp_823 = -exp_807;
  assign exp_815 = exp_787 == exp_814;
  assign exp_814 = 1;
  assign exp_880 = 0;
  assign exp_885 = 0;
  assign exp_873 = exp_872 + exp_871;
  assign exp_872 = 0;

  reg [31:0] exp_871_reg;
  always@(*) begin
    case (exp_868)
      0:exp_871_reg <= exp_866;
      1:exp_871_reg <= exp_869;
      default:exp_871_reg <= exp_870;
    endcase
  end
  assign exp_871 = exp_871_reg;
  assign exp_868 = exp_832 & exp_784;

      reg [0:0] exp_832_reg = 0;
      always@(posedge clk) begin
        if (exp_815) begin
          exp_832_reg <= exp_828;
        end
      end
      assign exp_832 = exp_832_reg;
      assign exp_828 = exp_810 ^ exp_813;
  assign exp_810 = exp_809 + exp_808;
  assign exp_809 = 0;
  assign exp_808 = exp_806[31:31];

      reg [31:0] exp_806_reg = 0;
      always@(posedge clk) begin
        if (exp_805) begin
          exp_806_reg <= exp_528;
        end
      end
      assign exp_806 = exp_806_reg;
      assign exp_870 = 0;

      reg [31:0] exp_866_reg = 0;
      always@(posedge clk) begin
        if (exp_799) begin
          exp_866_reg <= exp_836;
        end
      end
      assign exp_866 = exp_866_reg;
    
      reg [31:0] exp_836_reg = 0;
      always@(posedge clk) begin
        if (exp_835) begin
          exp_836_reg <= exp_863;
        end
      end
      assign exp_836 = exp_836_reg;
    
  reg [31:0] exp_863_reg;
  always@(*) begin
    case (exp_797)
      0:exp_863_reg <= exp_855;
      1:exp_863_reg <= exp_861;
      default:exp_863_reg <= exp_862;
    endcase
  end
  assign exp_863 = exp_863_reg;
  assign exp_797 = exp_787 == exp_796;
  assign exp_796 = 2;
  assign exp_862 = 0;

  reg [31:0] exp_855_reg;
  always@(*) begin
    case (exp_845)
      0:exp_855_reg <= exp_849;
      1:exp_855_reg <= exp_853;
      default:exp_855_reg <= exp_854;
    endcase
  end
  assign exp_855 = exp_855_reg;
  assign exp_845 = ~exp_844;
  assign exp_844 = exp_843[32:32];
  assign exp_843 = exp_842 - exp_830;
  assign exp_842 = exp_841;
  assign exp_841 = {exp_839, exp_840};  assign exp_839 = exp_834[31:0];

      reg [31:0] exp_834_reg = 0;
      always@(posedge clk) begin
        if (exp_833) begin
          exp_834_reg <= exp_860;
        end
      end
      assign exp_834 = exp_834_reg;
    
  reg [32:0] exp_860_reg;
  always@(*) begin
    case (exp_797)
      0:exp_860_reg <= exp_847;
      1:exp_860_reg <= exp_858;
      default:exp_860_reg <= exp_859;
    endcase
  end
  assign exp_860 = exp_860_reg;
  assign exp_859 = 0;

  reg [32:0] exp_847_reg;
  always@(*) begin
    case (exp_845)
      0:exp_847_reg <= exp_841;
      1:exp_847_reg <= exp_843;
      default:exp_847_reg <= exp_846;
    endcase
  end
  assign exp_847 = exp_847_reg;
  assign exp_846 = 0;
  assign exp_858 = 0;
  assign exp_833 = 1;
  assign exp_840 = exp_838[31:31];

      reg [31:0] exp_838_reg = 0;
      always@(posedge clk) begin
        if (exp_837) begin
          exp_838_reg <= exp_865;
        end
      end
      assign exp_838 = exp_838_reg;
    
  reg [31:0] exp_865_reg;
  always@(*) begin
    case (exp_797)
      0:exp_865_reg <= exp_857;
      1:exp_865_reg <= exp_829;
      default:exp_865_reg <= exp_864;
    endcase
  end
  assign exp_865 = exp_865_reg;
  assign exp_864 = 0;
  assign exp_857 = exp_838 << exp_856;
  assign exp_856 = 1;

      reg [31:0] exp_829_reg = 0;
      always@(posedge clk) begin
        if (exp_815) begin
          exp_829_reg <= exp_821;
        end
      end
      assign exp_829 = exp_829_reg;
      assign exp_821 = exp_820 + exp_819;
  assign exp_820 = 0;

  reg [31:0] exp_819_reg;
  always@(*) begin
    case (exp_816)
      0:exp_819_reg <= exp_806;
      1:exp_819_reg <= exp_817;
      default:exp_819_reg <= exp_818;
    endcase
  end
  assign exp_819 = exp_819_reg;
  assign exp_816 = exp_810 & exp_784;
  assign exp_818 = 0;
  assign exp_817 = -exp_806;
  assign exp_837 = 1;
  assign exp_854 = 0;
  assign exp_849 = exp_836 << exp_848;
  assign exp_848 = 1;
  assign exp_853 = exp_851 | exp_852;
  assign exp_851 = exp_836 << exp_850;
  assign exp_850 = 1;
  assign exp_852 = 1;
  assign exp_861 = 0;
  assign exp_835 = 1;
  assign exp_799 = exp_787 == exp_798;
  assign exp_798 = 35;
  assign exp_869 = -exp_866;
  assign exp_884 = $signed(exp_883);
  assign exp_883 = -1;
  assign exp_801 = exp_787 == exp_800;
  assign exp_800 = 36;

      reg [31:0] exp_893_reg = 0;
      always@(posedge clk) begin
        if (exp_801) begin
          exp_893_reg <= exp_891;
        end
      end
      assign exp_893 = exp_893_reg;
    
  reg [31:0] exp_891_reg;
  always@(*) begin
    case (exp_889)
      0:exp_891_reg <= exp_879;
      1:exp_891_reg <= exp_806;
      default:exp_891_reg <= exp_890;
    endcase
  end
  assign exp_891 = exp_891_reg;
  assign exp_889 = exp_888 & exp_784;
  assign exp_888 = exp_830 == exp_887;
  assign exp_887 = 0;
  assign exp_890 = 0;
  assign exp_879 = exp_878 + exp_877;
  assign exp_878 = 0;

  reg [31:0] exp_877_reg;
  always@(*) begin
    case (exp_874)
      0:exp_877_reg <= exp_867;
      1:exp_877_reg <= exp_875;
      default:exp_877_reg <= exp_876;
    endcase
  end
  assign exp_877 = exp_877_reg;
  assign exp_874 = exp_831 & exp_784;

      reg [0:0] exp_831_reg = 0;
      always@(posedge clk) begin
        if (exp_815) begin
          exp_831_reg <= exp_810;
        end
      end
      assign exp_831 = exp_831_reg;
      assign exp_876 = 0;

      reg [31:0] exp_867_reg = 0;
      always@(posedge clk) begin
        if (exp_799) begin
          exp_867_reg <= exp_834;
        end
      end
      assign exp_867 = exp_867_reg;
      assign exp_875 = -exp_867;
  assign exp_462 = $signed(exp_461);
  assign exp_461 = 0;
  assign exp_691 = exp_526 != exp_527;
  assign exp_704 = 0;
  assign exp_705 = 0;
  assign exp_692 = $signed(exp_526) < $signed(exp_527);
  assign exp_693 = $signed(exp_526) >= $signed(exp_527);
  assign exp_698 = exp_695 < exp_697;
  assign exp_695 = exp_694 + exp_526;
  assign exp_694 = 0;
  assign exp_697 = exp_696 + exp_527;
  assign exp_696 = 0;
  assign exp_703 = exp_700 >= exp_702;
  assign exp_700 = exp_699 + exp_526;
  assign exp_699 = 0;
  assign exp_702 = exp_701 + exp_527;
  assign exp_701 = 0;
  assign exp_1018 = 0;
  assign exp_1017 = exp_416 + exp_1016;
  assign exp_1016 = 4;

  reg [32:0] exp_748_reg;
  always@(*) begin
    case (exp_549)
      0:exp_748_reg <= exp_738;
      1:exp_748_reg <= exp_746;
      default:exp_748_reg <= exp_747;
    endcase
  end
  assign exp_748 = exp_748_reg;
  assign exp_747 = 0;
  assign exp_738 = exp_737 + exp_535;

  reg [31:0] exp_737_reg;
  always@(*) begin
    case (exp_547)
      0:exp_737_reg <= exp_723;
      1:exp_737_reg <= exp_735;
      default:exp_737_reg <= exp_736;
    endcase
  end
  assign exp_737 = exp_737_reg;
  assign exp_736 = 0;
  assign exp_723 = $signed(exp_722);
  assign exp_722 = exp_721 + exp_720;
  assign exp_721 = 0;
  assign exp_720 = {exp_719, exp_716};  assign exp_719 = {exp_718, exp_715};  assign exp_718 = {exp_717, exp_714};  assign exp_717 = {exp_712, exp_713};  assign exp_712 = exp_534[31:31];
  assign exp_713 = exp_534[7:7];
  assign exp_714 = exp_534[30:25];
  assign exp_715 = exp_534[11:8];
  assign exp_716 = 0;
  assign exp_735 = $signed(exp_734);
  assign exp_734 = exp_733 + exp_732;
  assign exp_733 = 0;
  assign exp_732 = {exp_731, exp_728};  assign exp_731 = {exp_730, exp_727};  assign exp_730 = {exp_729, exp_726};  assign exp_729 = {exp_724, exp_725};  assign exp_724 = exp_534[31:31];
  assign exp_725 = exp_534[19:12];
  assign exp_726 = exp_534[20:20];
  assign exp_727 = exp_534[30:21];
  assign exp_728 = 0;

      reg [31:0] exp_535_reg = 0;
      always@(posedge clk) begin
        if (exp_525) begin
          exp_535_reg <= exp_418;
        end
      end
      assign exp_535 = exp_535_reg;
      assign exp_746 = exp_745 & exp_744;
  assign exp_745 = $signed(exp_743);
  assign exp_743 = exp_526 + exp_742;
  assign exp_742 = $signed(exp_741);
  assign exp_741 = exp_740 + exp_739;
  assign exp_740 = 0;
  assign exp_739 = exp_534[31:20];
  assign exp_744 = 4294967294;
  assign exp_415 = exp_408 & exp_406;
  assign exp_88 = exp_92;
  assign exp_84 = exp_91;
  assign exp_86 = exp_91;
  assign exp_17 = exp_417;
  assign exp_550 = 3;
  assign exp_280 = exp_12;
  assign exp_313 = exp_301 & exp_312;
  assign exp_312 = ~exp_310;
  assign exp_310 = exp_304 & exp_301;
  assign exp_304 = exp_302 == exp_303;

      reg [8:0] exp_302_reg = 0;
      always@(posedge clk) begin
        if (exp_301) begin
          exp_302_reg <= exp_309;
        end
      end
      assign exp_302 = exp_302_reg;
    
  reg [8:0] exp_309_reg;
  always@(*) begin
    case (exp_304)
      0:exp_309_reg <= exp_306;
      1:exp_309_reg <= exp_307;
      default:exp_309_reg <= exp_308;
    endcase
  end
  assign exp_309 = exp_309_reg;
  assign exp_308 = 0;
  assign exp_306 = exp_302 + exp_305;
  assign exp_305 = 1;
  assign exp_307 = 0;
  assign exp_303 = 433;
  assign exp_300 = 1;
  assign exp_339 = exp_316 & exp_338;
  assign exp_338 = ~exp_337;
  assign exp_337 = exp_325 & exp_335;
  assign exp_325 = exp_319 & exp_316;
  assign exp_319 = exp_317 == exp_318;

      reg [8:0] exp_317_reg = 0;
      always@(posedge clk) begin
        if (exp_316) begin
          exp_317_reg <= exp_324;
        end
      end
      assign exp_317 = exp_317_reg;
    
  reg [8:0] exp_324_reg;
  always@(*) begin
    case (exp_319)
      0:exp_324_reg <= exp_321;
      1:exp_324_reg <= exp_322;
      default:exp_324_reg <= exp_323;
    endcase
  end
  assign exp_324 = exp_324_reg;
  assign exp_323 = 0;
  assign exp_321 = exp_317 + exp_320;
  assign exp_320 = 1;
  assign exp_322 = 0;
  assign exp_318 = 433;
  assign exp_335 = exp_329 & exp_326;
  assign exp_329 = exp_327 == exp_328;

      reg [2:0] exp_327_reg = 0;
      always@(posedge clk) begin
        if (exp_326) begin
          exp_327_reg <= exp_334;
        end
      end
      assign exp_327 = exp_327_reg;
    
  reg [2:0] exp_334_reg;
  always@(*) begin
    case (exp_329)
      0:exp_334_reg <= exp_331;
      1:exp_334_reg <= exp_332;
      default:exp_334_reg <= exp_333;
    endcase
  end
  assign exp_334 = exp_334_reg;
  assign exp_333 = 0;
  assign exp_331 = exp_327 + exp_330;
  assign exp_330 = 1;
  assign exp_332 = 0;
  assign exp_326 = exp_316 & exp_325;
  assign exp_328 = 7;
  assign exp_315 = 1;
  assign exp_355 = exp_342 & exp_354;
  assign exp_354 = ~exp_351;
  assign exp_351 = exp_345 & exp_342;
  assign exp_345 = exp_343 == exp_344;

      reg [8:0] exp_343_reg = 0;
      always@(posedge clk) begin
        if (exp_342) begin
          exp_343_reg <= exp_350;
        end
      end
      assign exp_343 = exp_343_reg;
    
  reg [8:0] exp_350_reg;
  always@(*) begin
    case (exp_345)
      0:exp_350_reg <= exp_347;
      1:exp_350_reg <= exp_348;
      default:exp_350_reg <= exp_349;
    endcase
  end
  assign exp_350 = exp_350_reg;
  assign exp_349 = 0;
  assign exp_347 = exp_343 + exp_346;
  assign exp_346 = 1;
  assign exp_348 = 0;
  assign exp_344 = 433;
  assign exp_341 = 1;
  assign exp_298 = exp_296 & exp_297;
  assign exp_297 = ~exp_293;
  assign exp_295 = 1;
  assign exp_374 = 0;

  reg [0:0] exp_371_reg;
  always@(*) begin
    case (exp_301)
      0:exp_371_reg <= exp_368;
      1:exp_371_reg <= exp_369;
      default:exp_371_reg <= exp_370;
    endcase
  end
  assign exp_371 = exp_371_reg;
  assign exp_370 = 0;
  assign exp_368 = exp_359[0:0];

      reg [7:0] exp_359_reg = 0;
      always@(posedge clk) begin
        if (exp_358) begin
          exp_359_reg <= exp_367;
        end
      end
      assign exp_359 = exp_359_reg;
    
  reg [7:0] exp_367_reg;
  always@(*) begin
    case (exp_365)
      0:exp_367_reg <= exp_364;
      1:exp_367_reg <= exp_292;
      default:exp_367_reg <= exp_366;
    endcase
  end
  assign exp_367 = exp_367_reg;
  assign exp_365 = exp_296 & exp_293;
  assign exp_366 = 0;

  reg [7:0] exp_364_reg;
  always@(*) begin
    case (exp_360)
      0:exp_364_reg <= exp_359;
      1:exp_364_reg <= exp_362;
      default:exp_364_reg <= exp_363;
    endcase
  end
  assign exp_364 = exp_364_reg;
  assign exp_360 = exp_316 & exp_325;
  assign exp_363 = 0;
  assign exp_362 = exp_359 >> exp_361;
  assign exp_361 = 1;
  assign exp_292 = exp_276[7:0];
  assign exp_276 = exp_10;
  assign exp_358 = 1;
  assign exp_369 = 0;
  assign exp_373 = 1;

      reg [31:0] exp_395_reg = 0;
      always@(posedge clk) begin
        if (exp_394) begin
          exp_395_reg <= exp_378;
        end
      end
      assign exp_395 = exp_395_reg;
      assign exp_378 = exp_10;
  assign exp_394 = exp_381 & exp_382;
  assign exp_381 = exp_389;
  assign exp_389 = exp_11 & exp_388;
  assign exp_382 = exp_12;
  assign stdout_tx = exp_375;
  assign leds_out = exp_395;

endmodule