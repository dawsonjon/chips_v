
module soc(clk, stdin_valid_in, stdin_in, stdout_ready_in, stdin_ready_out, stdout_valid_out, stdout_out, leds_out);
  input [0:0] stdin_valid_in;
  input [31:0] stdin_in;
  input [0:0] stdout_ready_in;
  input [0:0] clk;
  output [0:0] stdin_ready_out;
  output [0:0] stdout_valid_out;
  output [31:0] stdout_out;
  output [31:0] leds_out;
  wire [0:0] exp_245;
  wire [0:0] exp_228;
  wire [0:0] exp_236;
  wire [0:0] exp_5;
  wire [0:0] exp_250;
  wire [0:0] exp_597;
  wire [0:0] exp_534;
  wire [0:0] exp_399;
  wire [6:0] exp_384;
  wire [31:0] exp_382;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [11:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_264;
  wire [32:0] exp_867;
  wire [0:0] exp_863;
  wire [0:0] exp_559;
  wire [0:0] exp_537;
  wire [0:0] exp_395;
  wire [6:0] exp_394;
  wire [0:0] exp_397;
  wire [6:0] exp_396;
  wire [0:0] exp_558;
  wire [0:0] exp_403;
  wire [6:0] exp_402;
  wire [0:0] exp_557;
  wire [0:0] exp_556;
  wire [0:0] exp_555;
  wire [2:0] exp_385;
  wire [0:0] exp_554;
  wire [0:0] exp_538;
  wire [31:0] exp_374;
  wire [31:0] exp_312;
  wire [0:0] exp_308;
  wire [4:0] exp_288;
  wire [0:0] exp_307;
  wire [0:0] exp_311;
  wire [31:0] exp_304;
  wire [0:0] exp_285;
  wire [0:0] exp_858;
  wire [0:0] exp_857;
  wire [0:0] exp_856;
  wire [0:0] exp_855;
  wire [4:0] exp_267;
  wire [4:0] exp_850;
  wire [0:0] exp_849;
  wire [0:0] exp_441;
  wire [0:0] exp_440;
  wire [0:0] exp_439;
  wire [0:0] exp_438;
  wire [0:0] exp_437;
  wire [0:0] exp_436;
  wire [0:0] exp_387;
  wire [4:0] exp_386;
  wire [0:0] exp_389;
  wire [5:0] exp_388;
  wire [0:0] exp_391;
  wire [5:0] exp_390;
  wire [0:0] exp_393;
  wire [4:0] exp_392;
  wire [0:0] exp_844;
  wire [0:0] exp_843;
  wire [0:0] exp_629;
  wire [0:0] exp_603;
  wire [0:0] exp_601;
  wire [6:0] exp_599;
  wire [5:0] exp_600;
  wire [0:0] exp_602;
  wire [0:0] exp_628;
  wire [2:0] exp_598;
  wire [0:0] exp_842;
  wire [0:0] exp_840;
  wire [0:0] exp_833;
  wire [2:0] exp_748;
  wire [2:0] exp_755;
  wire [0:0] exp_750;
  wire [2:0] exp_749;
  wire [0:0] exp_754;
  wire [2:0] exp_752;
  wire [0:0] exp_751;
  wire [0:0] exp_753;
  wire [0:0] exp_744;
  wire [0:0] exp_743;
  wire [0:0] exp_742;
  wire [2:0] exp_832;
  wire [0:0] exp_841;
  wire [0:0] exp_651;
  wire [5:0] exp_635;
  wire [5:0] exp_642;
  wire [0:0] exp_637;
  wire [5:0] exp_636;
  wire [0:0] exp_641;
  wire [5:0] exp_639;
  wire [0:0] exp_638;
  wire [0:0] exp_640;
  wire [5:0] exp_650;
  wire [0:0] exp_262;
  wire [0:0] exp_261;
  wire [0:0] exp_259;
  wire [0:0] exp_258;
  wire [0:0] exp_256;
  wire [0:0] exp_257;
  wire [0:0] exp_255;
  wire [0:0] exp_868;
  wire [0:0] exp_254;
  wire [0:0] exp_253;
  wire [0:0] exp_872;
  wire [0:0] exp_871;
  wire [0:0] exp_870;
  wire [0:0] exp_869;
  wire [0:0] exp_249;
  wire [0:0] exp_240;
  wire [0:0] exp_235;
  wire [0:0] exp_232;
  wire [31:0] exp_1;
  wire [31:0] exp_246;
  wire [31:0] exp_453;
  wire [31:0] exp_452;
  wire [31:0] exp_451;
  wire [31:0] exp_450;
  wire [11:0] exp_449;
  wire [11:0] exp_448;
  wire [11:0] exp_447;
  wire [0:0] exp_401;
  wire [5:0] exp_400;
  wire [0:0] exp_446;
  wire [11:0] exp_442;
  wire [11:0] exp_445;
  wire [6:0] exp_443;
  wire [4:0] exp_444;
  wire [31:0] exp_231;
  wire [0:0] exp_234;
  wire [31:0] exp_233;
  wire [0:0] exp_239;
  wire [0:0] exp_218;
  wire [0:0] exp_213;
  wire [0:0] exp_210;
  wire [31:0] exp_209;
  wire [0:0] exp_212;
  wire [31:0] exp_211;
  wire [0:0] exp_217;
  wire [0:0] exp_196;
  wire [0:0] exp_191;
  wire [0:0] exp_188;
  wire [31:0] exp_187;
  wire [0:0] exp_190;
  wire [31:0] exp_189;
  wire [0:0] exp_195;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [31:0] exp_146;
  wire [0:0] exp_149;
  wire [31:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [13:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_251;
  wire [0:0] exp_536;
  wire [0:0] exp_535;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_176;
  wire [0:0] exp_183;
  wire [0:0] exp_198;
  wire [0:0] exp_205;
  wire [0:0] exp_223;
  wire [0:0] exp_227;
  wire [0:0] exp_243;
  wire [0:0] exp_846;
  wire [0:0] exp_845;
  wire [0:0] exp_260;
  wire [0:0] exp_303;
  wire [31:0] exp_275;
  wire [0:0] exp_274;
  wire [1:0] exp_283;
  wire [4:0] exp_270;
  wire [0:0] exp_273;
  wire [0:0] exp_852;
  wire [0:0] exp_851;
  wire [4:0] exp_269;
  wire [31:0] exp_271;
  wire [31:0] exp_848;
  wire [0:0] exp_847;
  wire [31:0] exp_484;
  wire [0:0] exp_483;
  wire [31:0] exp_435;
  wire [2:0] exp_378;
  wire [2:0] exp_369;
  wire [0:0] exp_366;
  wire [0:0] exp_300;
  wire [6:0] exp_290;
  wire [6:0] exp_299;
  wire [0:0] exp_302;
  wire [6:0] exp_301;
  wire [0:0] exp_368;
  wire [2:0] exp_356;
  wire [0:0] exp_298;
  wire [4:0] exp_297;
  wire [0:0] exp_355;
  wire [2:0] exp_343;
  wire [0:0] exp_296;
  wire [5:0] exp_295;
  wire [0:0] exp_342;
  wire [2:0] exp_292;
  wire [0:0] exp_341;
  wire [0:0] exp_354;
  wire [0:0] exp_367;
  wire [0:0] exp_373;
  wire [0:0] exp_434;
  wire [31:0] exp_414;
  wire [0:0] exp_380;
  wire [0:0] exp_372;
  wire [0:0] exp_358;
  wire [0:0] exp_345;
  wire [0:0] exp_331;
  wire [0:0] exp_329;
  wire [0:0] exp_330;
  wire [0:0] exp_294;
  wire [4:0] exp_293;
  wire [0:0] exp_344;
  wire [0:0] exp_357;
  wire [0:0] exp_371;
  wire [0:0] exp_370;
  wire [0:0] exp_413;
  wire [31:0] exp_411;
  wire [31:0] exp_376;
  wire [31:0] exp_362;
  wire [0:0] exp_359;
  wire [0:0] exp_361;
  wire [31:0] exp_351;
  wire [0:0] exp_350;
  wire [31:0] exp_337;
  wire [0:0] exp_336;
  wire [31:0] exp_335;
  wire [31:0] exp_333;
  wire [19:0] exp_332;
  wire [3:0] exp_334;
  wire [31:0] exp_349;
  wire [31:0] exp_347;
  wire [19:0] exp_346;
  wire [3:0] exp_348;
  wire [31:0] exp_360;
  wire [31:0] exp_377;
  wire [31:0] exp_365;
  wire [0:0] exp_363;
  wire [0:0] exp_364;
  wire [31:0] exp_353;
  wire [0:0] exp_352;
  wire [31:0] exp_340;
  wire [0:0] exp_339;
  wire [31:0] exp_324;
  wire [0:0] exp_323;
  wire [31:0] exp_318;
  wire [0:0] exp_314;
  wire [4:0] exp_289;
  wire [0:0] exp_313;
  wire [0:0] exp_317;
  wire [31:0] exp_306;
  wire [0:0] exp_286;
  wire [0:0] exp_862;
  wire [0:0] exp_861;
  wire [0:0] exp_860;
  wire [0:0] exp_859;
  wire [4:0] exp_268;
  wire [0:0] exp_305;
  wire [31:0] exp_282;
  wire [0:0] exp_281;
  wire [1:0] exp_284;
  wire [4:0] exp_277;
  wire [0:0] exp_280;
  wire [0:0] exp_854;
  wire [0:0] exp_853;
  wire [4:0] exp_276;
  wire [31:0] exp_278;
  wire [31:0] exp_287;
  wire [31:0] exp_316;
  wire [0:0] exp_315;
  wire [31:0] exp_322;
  wire [31:0] exp_319;
  wire [31:0] exp_321;
  wire [11:0] exp_320;
  wire [31:0] exp_338;
  wire [31:0] exp_266;
  wire [0:0] exp_265;
  wire [31:0] exp_412;
  wire [31:0] exp_416;
  wire [31:0] exp_415;
  wire [5:0] exp_410;
  wire [5:0] exp_409;
  wire [5:0] exp_408;
  wire [4:0] exp_379;
  wire [4:0] exp_328;
  wire [0:0] exp_327;
  wire [4:0] exp_326;
  wire [4:0] exp_291;
  wire [31:0] exp_432;
  wire [1:0] exp_418;
  wire [0:0] exp_417;
  wire [31:0] exp_433;
  wire [1:0] exp_424;
  wire [0:0] exp_423;
  wire [31:0] exp_420;
  wire [31:0] exp_419;
  wire [31:0] exp_422;
  wire [31:0] exp_421;
  wire [31:0] exp_425;
  wire [31:0] exp_429;
  wire [32:0] exp_428;
  wire [32:0] exp_426;
  wire [0:0] exp_407;
  wire [0:0] exp_381;
  wire [0:0] exp_325;
  wire [0:0] exp_406;
  wire [0:0] exp_405;
  wire [0:0] exp_404;
  wire [32:0] exp_427;
  wire [31:0] exp_430;
  wire [31:0] exp_431;
  wire [31:0] exp_482;
  wire [0:0] exp_481;
  wire [31:0] exp_472;
  wire [7:0] exp_471;
  wire [7:0] exp_470;
  wire [7:0] exp_465;
  wire [1:0] exp_456;
  wire [1:0] exp_455;
  wire [1:0] exp_454;
  wire [0:0] exp_464;
  wire [7:0] exp_460;
  wire [31:0] exp_248;
  wire [31:0] exp_238;
  wire [0:0] exp_237;
  wire [31:0] exp_216;
  wire [0:0] exp_215;
  wire [31:0] exp_194;
  wire [0:0] exp_193;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [11:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_252;
  wire [3:0] exp_533;
  wire [0:0] exp_532;
  wire [3:0] exp_520;
  wire [3:0] exp_516;
  wire [1:0] exp_519;
  wire [1:0] exp_518;
  wire [1:0] exp_517;
  wire [3:0] exp_525;
  wire [3:0] exp_521;
  wire [0:0] exp_524;
  wire [0:0] exp_523;
  wire [0:0] exp_522;
  wire [3:0] exp_526;
  wire [3:0] exp_527;
  wire [3:0] exp_528;
  wire [3:0] exp_529;
  wire [3:0] exp_530;
  wire [3:0] exp_531;
  wire [11:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_247;
  wire [31:0] exp_515;
  wire [0:0] exp_514;
  wire [31:0] exp_502;
  wire [0:0] exp_501;
  wire [31:0] exp_488;
  wire [7:0] exp_487;
  wire [7:0] exp_486;
  wire [7:0] exp_485;
  wire [31:0] exp_375;
  wire [31:0] exp_496;
  wire [3:0] exp_495;
  wire [31:0] exp_498;
  wire [4:0] exp_497;
  wire [31:0] exp_500;
  wire [4:0] exp_499;
  wire [31:0] exp_506;
  wire [0:0] exp_459;
  wire [0:0] exp_458;
  wire [0:0] exp_457;
  wire [0:0] exp_505;
  wire [31:0] exp_492;
  wire [15:0] exp_491;
  wire [15:0] exp_490;
  wire [15:0] exp_489;
  wire [31:0] exp_504;
  wire [4:0] exp_503;
  wire [31:0] exp_508;
  wire [31:0] exp_507;
  wire [31:0] exp_494;
  wire [31:0] exp_493;
  wire [31:0] exp_509;
  wire [31:0] exp_510;
  wire [31:0] exp_511;
  wire [31:0] exp_512;
  wire [31:0] exp_513;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [11:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [11:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [11:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [11:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [11:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [11:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [11:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [11:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [11:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [11:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [11:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [11:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_179;
  wire [0:0] exp_177;
  wire [31:0] exp_139;
  wire [0:0] exp_178;
  wire [31:0] exp_157;
  wire [31:0] exp_164;
  wire [0:0] exp_159;
  wire [31:0] exp_158;
  wire [0:0] exp_163;
  wire [31:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [31:0] exp_167;
  wire [31:0] exp_174;
  wire [0:0] exp_169;
  wire [31:0] exp_168;
  wire [0:0] exp_173;
  wire [31:0] exp_171;
  wire [0:0] exp_170;
  wire [0:0] exp_172;
  wire [0:0] exp_166;
  wire [0:0] exp_165;
  wire [31:0] exp_182;
  wire [31:0] exp_201;
  wire [31:0] exp_204;
  wire [31:0] exp_222;
  wire [31:0] exp_226;
  wire [31:0] exp_241;
  wire [7:0] exp_461;
  wire [7:0] exp_462;
  wire [7:0] exp_463;
  wire [31:0] exp_475;
  wire [15:0] exp_474;
  wire [15:0] exp_473;
  wire [15:0] exp_469;
  wire [0:0] exp_468;
  wire [15:0] exp_466;
  wire [15:0] exp_467;
  wire [31:0] exp_476;
  wire [31:0] exp_477;
  wire [31:0] exp_478;
  wire [31:0] exp_479;
  wire [31:0] exp_480;
  wire [31:0] exp_839;
  wire [0:0] exp_838;
  wire [31:0] exp_835;
  wire [0:0] exp_606;
  wire [0:0] exp_605;
  wire [0:0] exp_604;
  wire [0:0] exp_834;
  wire [31:0] exp_830;
  wire [63:0] exp_829;
  wire [0:0] exp_826;
  wire [0:0] exp_809;
  wire [0:0] exp_786;
  wire [0:0] exp_783;
  wire [0:0] exp_781;
  wire [0:0] exp_763;
  wire [0:0] exp_762;
  wire [0:0] exp_761;
  wire [31:0] exp_759;
  wire [0:0] exp_758;
  wire [0:0] exp_757;
  wire [0:0] exp_746;
  wire [0:0] exp_745;
  wire [0:0] exp_609;
  wire [0:0] exp_608;
  wire [0:0] exp_607;
  wire [0:0] exp_612;
  wire [0:0] exp_611;
  wire [1:0] exp_610;
  wire [0:0] exp_782;
  wire [0:0] exp_766;
  wire [0:0] exp_765;
  wire [0:0] exp_764;
  wire [31:0] exp_760;
  wire [0:0] exp_747;
  wire [0:0] exp_768;
  wire [0:0] exp_767;
  wire [0:0] exp_788;
  wire [1:0] exp_787;
  wire [0:0] exp_811;
  wire [1:0] exp_810;
  wire [0:0] exp_828;
  wire [63:0] exp_825;
  wire [63:0] exp_824;
  wire [63:0] exp_820;
  wire [63:0] exp_816;
  wire [63:0] exp_812;
  wire [31:0] exp_805;
  wire [31:0] exp_792;
  wire [31:0] exp_790;
  wire [15:0] exp_789;
  wire [31:0] exp_784;
  wire [31:0] exp_774;
  wire [31:0] exp_773;
  wire [31:0] exp_772;
  wire [0:0] exp_769;
  wire [0:0] exp_771;
  wire [31:0] exp_770;
  wire [15:0] exp_791;
  wire [31:0] exp_785;
  wire [31:0] exp_780;
  wire [31:0] exp_779;
  wire [31:0] exp_778;
  wire [0:0] exp_775;
  wire [0:0] exp_777;
  wire [31:0] exp_776;
  wire [63:0] exp_815;
  wire [63:0] exp_813;
  wire [31:0] exp_806;
  wire [31:0] exp_796;
  wire [31:0] exp_794;
  wire [15:0] exp_793;
  wire [15:0] exp_795;
  wire [4:0] exp_814;
  wire [63:0] exp_819;
  wire [63:0] exp_817;
  wire [31:0] exp_807;
  wire [31:0] exp_800;
  wire [31:0] exp_798;
  wire [15:0] exp_797;
  wire [15:0] exp_799;
  wire [4:0] exp_818;
  wire [63:0] exp_823;
  wire [63:0] exp_821;
  wire [31:0] exp_808;
  wire [31:0] exp_804;
  wire [31:0] exp_802;
  wire [15:0] exp_801;
  wire [15:0] exp_803;
  wire [5:0] exp_822;
  wire [63:0] exp_827;
  wire [31:0] exp_831;
  wire [31:0] exp_837;
  wire [0:0] exp_630;
  wire [0:0] exp_836;
  wire [31:0] exp_740;
  wire [31:0] exp_734;
  wire [0:0] exp_730;
  wire [0:0] exp_729;
  wire [31:0] exp_678;
  wire [31:0] exp_675;
  wire [31:0] exp_674;
  wire [31:0] exp_673;
  wire [0:0] exp_670;
  wire [0:0] exp_661;
  wire [0:0] exp_660;
  wire [0:0] exp_659;
  wire [31:0] exp_655;
  wire [0:0] exp_653;
  wire [0:0] exp_652;
  wire [0:0] exp_632;
  wire [0:0] exp_631;
  wire [0:0] exp_672;
  wire [31:0] exp_671;
  wire [0:0] exp_663;
  wire [0:0] exp_662;
  wire [0:0] exp_728;
  wire [0:0] exp_733;
  wire [31:0] exp_721;
  wire [31:0] exp_720;
  wire [31:0] exp_719;
  wire [0:0] exp_716;
  wire [0:0] exp_680;
  wire [0:0] exp_676;
  wire [0:0] exp_658;
  wire [0:0] exp_657;
  wire [0:0] exp_656;
  wire [31:0] exp_654;
  wire [0:0] exp_718;
  wire [31:0] exp_714;
  wire [31:0] exp_684;
  wire [31:0] exp_711;
  wire [0:0] exp_645;
  wire [1:0] exp_644;
  wire [0:0] exp_710;
  wire [31:0] exp_703;
  wire [0:0] exp_693;
  wire [0:0] exp_692;
  wire [32:0] exp_691;
  wire [32:0] exp_690;
  wire [32:0] exp_689;
  wire [31:0] exp_687;
  wire [31:0] exp_682;
  wire [32:0] exp_708;
  wire [0:0] exp_707;
  wire [32:0] exp_695;
  wire [0:0] exp_694;
  wire [0:0] exp_706;
  wire [0:0] exp_681;
  wire [0:0] exp_688;
  wire [31:0] exp_686;
  wire [31:0] exp_713;
  wire [0:0] exp_712;
  wire [31:0] exp_705;
  wire [0:0] exp_704;
  wire [31:0] exp_677;
  wire [31:0] exp_669;
  wire [31:0] exp_668;
  wire [31:0] exp_667;
  wire [0:0] exp_664;
  wire [0:0] exp_666;
  wire [31:0] exp_665;
  wire [0:0] exp_685;
  wire [0:0] exp_702;
  wire [31:0] exp_697;
  wire [0:0] exp_696;
  wire [31:0] exp_701;
  wire [31:0] exp_699;
  wire [0:0] exp_698;
  wire [0:0] exp_700;
  wire [0:0] exp_709;
  wire [0:0] exp_683;
  wire [0:0] exp_647;
  wire [5:0] exp_646;
  wire [31:0] exp_717;
  wire [31:0] exp_732;
  wire [0:0] exp_731;
  wire [0:0] exp_649;
  wire [5:0] exp_648;
  wire [31:0] exp_741;
  wire [31:0] exp_739;
  wire [0:0] exp_737;
  wire [0:0] exp_736;
  wire [0:0] exp_735;
  wire [0:0] exp_738;
  wire [31:0] exp_727;
  wire [31:0] exp_726;
  wire [31:0] exp_725;
  wire [0:0] exp_722;
  wire [0:0] exp_679;
  wire [0:0] exp_724;
  wire [31:0] exp_715;
  wire [31:0] exp_723;
  wire [31:0] exp_310;
  wire [0:0] exp_309;
  wire [0:0] exp_539;
  wire [0:0] exp_552;
  wire [0:0] exp_553;
  wire [0:0] exp_540;
  wire [0:0] exp_541;
  wire [0:0] exp_546;
  wire [31:0] exp_543;
  wire [31:0] exp_542;
  wire [31:0] exp_545;
  wire [31:0] exp_544;
  wire [0:0] exp_551;
  wire [31:0] exp_548;
  wire [31:0] exp_547;
  wire [31:0] exp_550;
  wire [31:0] exp_549;
  wire [0:0] exp_866;
  wire [31:0] exp_865;
  wire [2:0] exp_864;
  wire [32:0] exp_596;
  wire [0:0] exp_595;
  wire [31:0] exp_586;
  wire [31:0] exp_585;
  wire [0:0] exp_584;
  wire [31:0] exp_571;
  wire [12:0] exp_570;
  wire [12:0] exp_569;
  wire [12:0] exp_568;
  wire [11:0] exp_567;
  wire [7:0] exp_566;
  wire [1:0] exp_565;
  wire [0:0] exp_560;
  wire [0:0] exp_561;
  wire [5:0] exp_562;
  wire [3:0] exp_563;
  wire [0:0] exp_564;
  wire [31:0] exp_583;
  wire [20:0] exp_582;
  wire [20:0] exp_581;
  wire [20:0] exp_580;
  wire [19:0] exp_579;
  wire [9:0] exp_578;
  wire [8:0] exp_577;
  wire [0:0] exp_572;
  wire [7:0] exp_573;
  wire [0:0] exp_574;
  wire [9:0] exp_575;
  wire [0:0] exp_576;
  wire [31:0] exp_383;
  wire [32:0] exp_594;
  wire [32:0] exp_593;
  wire [31:0] exp_591;
  wire [31:0] exp_590;
  wire [11:0] exp_589;
  wire [11:0] exp_588;
  wire [11:0] exp_587;
  wire [32:0] exp_592;
  wire [0:0] exp_263;
  wire [0:0] exp_80;
  wire [11:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_398;
  wire [0:0] exp_244;
  wire [0:0] exp_229;
  wire [0:0] exp_200;
  wire [0:0] exp_184;
  wire [0:0] exp_192;
  wire [0:0] exp_185;
  wire [31:0] exp_181;
  wire [31:0] exp_221;
  wire [31:0] exp_203;
  wire [0:0] exp_220;
  wire [0:0] exp_206;
  wire [0:0] exp_214;
  wire [0:0] exp_207;

  assign exp_245 = exp_228 & exp_244;
  assign exp_228 = exp_236;
  assign exp_236 = exp_5 & exp_235;
  assign exp_5 = exp_250;
  assign exp_250 = exp_597;
  assign exp_597 = exp_534 & exp_262;
  assign exp_534 = exp_399 | exp_401;
  assign exp_399 = exp_384 == exp_398;
  assign exp_384 = exp_382[6:0];

      reg [31:0] exp_382_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_382_reg <= exp_96;
        end
      end
      assign exp_382 = exp_382_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_264;

      reg [31:0] exp_264_reg = 0;
      always@(posedge clk) begin
        if (exp_263) begin
          exp_264_reg <= exp_867;
        end
      end
      assign exp_264 = exp_264_reg;
    
  reg [32:0] exp_867_reg;
  always@(*) begin
    case (exp_863)
      0:exp_867_reg <= exp_865;
      1:exp_867_reg <= exp_596;
      default:exp_867_reg <= exp_866;
    endcase
  end
  assign exp_867 = exp_867_reg;
  assign exp_863 = exp_559 & exp_262;
  assign exp_559 = exp_537 | exp_558;
  assign exp_537 = exp_395 | exp_397;
  assign exp_395 = exp_384 == exp_394;
  assign exp_394 = 111;
  assign exp_397 = exp_384 == exp_396;
  assign exp_396 = 103;

  reg [0:0] exp_558_reg;
  always@(*) begin
    case (exp_403)
      0:exp_558_reg <= exp_556;
      1:exp_558_reg <= exp_555;
      default:exp_558_reg <= exp_557;
    endcase
  end
  assign exp_558 = exp_558_reg;
  assign exp_403 = exp_384 == exp_402;
  assign exp_402 = 99;
  assign exp_557 = 0;
  assign exp_556 = 0;

  reg [0:0] exp_555_reg;
  always@(*) begin
    case (exp_385)
      0:exp_555_reg <= exp_538;
      1:exp_555_reg <= exp_539;
      2:exp_555_reg <= exp_552;
      3:exp_555_reg <= exp_553;
      4:exp_555_reg <= exp_540;
      5:exp_555_reg <= exp_541;
      6:exp_555_reg <= exp_546;
      7:exp_555_reg <= exp_551;
      default:exp_555_reg <= exp_554;
    endcase
  end
  assign exp_555 = exp_555_reg;
  assign exp_385 = exp_382[14:12];
  assign exp_554 = 0;
  assign exp_538 = exp_374 == exp_375;

      reg [31:0] exp_374_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_374_reg <= exp_312;
        end
      end
      assign exp_374 = exp_374_reg;
    
  reg [31:0] exp_312_reg;
  always@(*) begin
    case (exp_308)
      0:exp_312_reg <= exp_304;
      1:exp_312_reg <= exp_310;
      default:exp_312_reg <= exp_311;
    endcase
  end
  assign exp_312 = exp_312_reg;
  assign exp_308 = exp_288 == exp_307;
  assign exp_288 = exp_96[19:15];
  assign exp_307 = 0;
  assign exp_311 = 0;

  reg [31:0] exp_304_reg;
  always@(*) begin
    case (exp_285)
      0:exp_304_reg <= exp_275;
      1:exp_304_reg <= exp_287;
      default:exp_304_reg <= exp_303;
    endcase
  end
  assign exp_304 = exp_304_reg;
  assign exp_285 = exp_858;
  assign exp_858 = exp_857 & exp_254;
  assign exp_857 = exp_856 & exp_262;
  assign exp_856 = exp_855 & exp_849;
  assign exp_855 = exp_267 == exp_850;
  assign exp_267 = exp_96[19:15];
  assign exp_850 = exp_382[11:7];
  assign exp_849 = exp_441 | exp_844;
  assign exp_441 = exp_440 | exp_399;
  assign exp_440 = exp_439 | exp_393;
  assign exp_439 = exp_438 | exp_391;
  assign exp_438 = exp_437 | exp_397;
  assign exp_437 = exp_436 | exp_395;
  assign exp_436 = exp_387 | exp_389;
  assign exp_387 = exp_384 == exp_386;
  assign exp_386 = 19;
  assign exp_389 = exp_384 == exp_388;
  assign exp_388 = 51;
  assign exp_391 = exp_384 == exp_390;
  assign exp_390 = 55;
  assign exp_393 = exp_384 == exp_392;
  assign exp_392 = 23;
  assign exp_844 = exp_843 & exp_603;

  reg [0:0] exp_843_reg;
  always@(*) begin
    case (exp_629)
      0:exp_843_reg <= exp_840;
      1:exp_843_reg <= exp_841;
      default:exp_843_reg <= exp_842;
    endcase
  end
  assign exp_843 = exp_843_reg;
  assign exp_629 = exp_603 & exp_628;
  assign exp_603 = exp_601 & exp_602;
  assign exp_601 = exp_599 == exp_600;
  assign exp_599 = exp_382[6:0];
  assign exp_600 = 51;
  assign exp_602 = exp_382[25:25];
  assign exp_628 = exp_598[2:2];
  assign exp_598 = exp_382[14:12];
  assign exp_842 = 0;
  assign exp_840 = exp_833 & exp_603;
  assign exp_833 = exp_748 == exp_832;

      reg [2:0] exp_748_reg = 0;
      always@(posedge clk) begin
        if (exp_744) begin
          exp_748_reg <= exp_755;
        end
      end
      assign exp_748 = exp_748_reg;
    
  reg [2:0] exp_755_reg;
  always@(*) begin
    case (exp_750)
      0:exp_755_reg <= exp_752;
      1:exp_755_reg <= exp_753;
      default:exp_755_reg <= exp_754;
    endcase
  end
  assign exp_755 = exp_755_reg;
  assign exp_750 = exp_748 == exp_749;
  assign exp_749 = 4;
  assign exp_754 = 0;
  assign exp_752 = exp_748 + exp_751;
  assign exp_751 = 1;
  assign exp_753 = 0;
  assign exp_744 = exp_603 & exp_743;
  assign exp_743 = ~exp_742;
  assign exp_742 = exp_598[2:2];
  assign exp_832 = 4;
  assign exp_841 = exp_651 & exp_603;
  assign exp_651 = exp_635 == exp_650;

      reg [5:0] exp_635_reg = 0;
      always@(posedge clk) begin
        if (exp_629) begin
          exp_635_reg <= exp_642;
        end
      end
      assign exp_635 = exp_635_reg;
    
  reg [5:0] exp_642_reg;
  always@(*) begin
    case (exp_637)
      0:exp_642_reg <= exp_639;
      1:exp_642_reg <= exp_640;
      default:exp_642_reg <= exp_641;
    endcase
  end
  assign exp_642 = exp_642_reg;
  assign exp_637 = exp_635 == exp_636;
  assign exp_636 = 37;
  assign exp_641 = 0;
  assign exp_639 = exp_635 + exp_638;
  assign exp_638 = 1;
  assign exp_640 = 0;
  assign exp_650 = 37;

      reg [0:0] exp_262_reg = 0;
      always@(posedge clk) begin
        if (exp_254) begin
          exp_262_reg <= exp_261;
        end
      end
      assign exp_262 = exp_262_reg;
      assign exp_261 = exp_259 & exp_260;

      reg [0:0] exp_259_reg = 0;
      always@(posedge clk) begin
        if (exp_254) begin
          exp_259_reg <= exp_258;
        end
      end
      assign exp_259 = exp_259_reg;
      assign exp_258 = exp_256 & exp_257;
  assign exp_256 = 1;
  assign exp_257 = ~exp_255;
  assign exp_255 = exp_868;
  assign exp_868 = exp_262 & exp_559;
  assign exp_254 = ~exp_253;
  assign exp_253 = exp_872;
  assign exp_872 = exp_262 & exp_871;
  assign exp_871 = exp_870 | exp_846;
  assign exp_870 = exp_250 & exp_869;
  assign exp_869 = ~exp_249;
  assign exp_249 = exp_240;

  reg [0:0] exp_240_reg;
  always@(*) begin
    case (exp_235)
      0:exp_240_reg <= exp_218;
      1:exp_240_reg <= exp_227;
      default:exp_240_reg <= exp_239;
    endcase
  end
  assign exp_240 = exp_240_reg;
  assign exp_235 = exp_232 & exp_234;
  assign exp_232 = exp_1 >= exp_231;
  assign exp_1 = exp_246;
  assign exp_246 = exp_453;
  assign exp_453 = exp_452 + exp_451;
  assign exp_452 = 0;
  assign exp_451 = exp_374 + exp_450;
  assign exp_450 = $signed(exp_449);
  assign exp_449 = exp_448 + exp_447;
  assign exp_448 = 0;

  reg [11:0] exp_447_reg;
  always@(*) begin
    case (exp_401)
      0:exp_447_reg <= exp_442;
      1:exp_447_reg <= exp_445;
      default:exp_447_reg <= exp_446;
    endcase
  end
  assign exp_447 = exp_447_reg;
  assign exp_401 = exp_384 == exp_400;
  assign exp_400 = 35;
  assign exp_446 = 0;
  assign exp_442 = exp_382[31:20];
  assign exp_445 = {exp_443, exp_444};  assign exp_443 = exp_382[31:25];
  assign exp_444 = exp_382[11:7];
  assign exp_231 = 2147483664;
  assign exp_234 = exp_1 <= exp_233;
  assign exp_233 = 2147483664;
  assign exp_239 = 0;

  reg [0:0] exp_218_reg;
  always@(*) begin
    case (exp_213)
      0:exp_218_reg <= exp_196;
      1:exp_218_reg <= exp_205;
      default:exp_218_reg <= exp_217;
    endcase
  end
  assign exp_218 = exp_218_reg;
  assign exp_213 = exp_210 & exp_212;
  assign exp_210 = exp_1 >= exp_209;
  assign exp_209 = 2147483660;
  assign exp_212 = exp_1 <= exp_211;
  assign exp_211 = 2147483660;
  assign exp_217 = 0;

  reg [0:0] exp_196_reg;
  always@(*) begin
    case (exp_191)
      0:exp_196_reg <= exp_155;
      1:exp_196_reg <= exp_183;
      default:exp_196_reg <= exp_195;
    endcase
  end
  assign exp_196 = exp_196_reg;
  assign exp_191 = exp_188 & exp_190;
  assign exp_188 = exp_1 >= exp_187;
  assign exp_187 = 2147483656;
  assign exp_190 = exp_1 <= exp_189;
  assign exp_189 = 2147483656;
  assign exp_195 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 2147483648;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 2147483652;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 16380;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_251;
  assign exp_251 = exp_536;
  assign exp_536 = exp_535 + exp_401;
  assign exp_535 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_176;
  assign exp_176 = 1;
  assign exp_183 = exp_198;
  assign exp_198 = stdout_ready_in;
  assign exp_205 = exp_223;
  assign exp_223 = 1;
  assign exp_227 = exp_243;
  assign exp_243 = stdin_valid_in;
  assign exp_846 = exp_603 & exp_845;
  assign exp_845 = ~exp_843;
  assign exp_260 = ~exp_255;
  assign exp_303 = 0;

  //Create RAM
  reg [31:0] exp_275_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_273) begin
      exp_275_ram[exp_269] <= exp_271;
    end
  end
  assign exp_275 = exp_275_ram[exp_270];
  assign exp_274 = exp_283;
  assign exp_283 = 1;
  assign exp_270 = exp_267;
  assign exp_273 = exp_852;
  assign exp_852 = exp_851 & exp_254;
  assign exp_851 = exp_849 & exp_262;
  assign exp_269 = exp_850;
  assign exp_271 = exp_848;

  reg [31:0] exp_848_reg;
  always@(*) begin
    case (exp_844)
      0:exp_848_reg <= exp_484;
      1:exp_848_reg <= exp_839;
      default:exp_848_reg <= exp_847;
    endcase
  end
  assign exp_848 = exp_848_reg;
  assign exp_847 = 0;

  reg [31:0] exp_484_reg;
  always@(*) begin
    case (exp_399)
      0:exp_484_reg <= exp_435;
      1:exp_484_reg <= exp_482;
      default:exp_484_reg <= exp_483;
    endcase
  end
  assign exp_484 = exp_484_reg;
  assign exp_483 = 0;

  reg [31:0] exp_435_reg;
  always@(*) begin
    case (exp_378)
      0:exp_435_reg <= exp_414;
      1:exp_435_reg <= exp_416;
      2:exp_435_reg <= exp_432;
      3:exp_435_reg <= exp_433;
      4:exp_435_reg <= exp_425;
      5:exp_435_reg <= exp_429;
      6:exp_435_reg <= exp_430;
      7:exp_435_reg <= exp_431;
      default:exp_435_reg <= exp_434;
    endcase
  end
  assign exp_435 = exp_435_reg;

      reg [2:0] exp_378_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_378_reg <= exp_369;
        end
      end
      assign exp_378 = exp_378_reg;
    
  reg [2:0] exp_369_reg;
  always@(*) begin
    case (exp_366)
      0:exp_369_reg <= exp_356;
      1:exp_369_reg <= exp_367;
      default:exp_369_reg <= exp_368;
    endcase
  end
  assign exp_369 = exp_369_reg;
  assign exp_366 = exp_300 | exp_302;
  assign exp_300 = exp_290 == exp_299;
  assign exp_290 = exp_96[6:0];
  assign exp_299 = 111;
  assign exp_302 = exp_290 == exp_301;
  assign exp_301 = 103;
  assign exp_368 = 0;

  reg [2:0] exp_356_reg;
  always@(*) begin
    case (exp_298)
      0:exp_356_reg <= exp_343;
      1:exp_356_reg <= exp_354;
      default:exp_356_reg <= exp_355;
    endcase
  end
  assign exp_356 = exp_356_reg;
  assign exp_298 = exp_290 == exp_297;
  assign exp_297 = 23;
  assign exp_355 = 0;

  reg [2:0] exp_343_reg;
  always@(*) begin
    case (exp_296)
      0:exp_343_reg <= exp_292;
      1:exp_343_reg <= exp_341;
      default:exp_343_reg <= exp_342;
    endcase
  end
  assign exp_343 = exp_343_reg;
  assign exp_296 = exp_290 == exp_295;
  assign exp_295 = 55;
  assign exp_342 = 0;
  assign exp_292 = exp_96[14:12];
  assign exp_341 = 0;
  assign exp_354 = 0;
  assign exp_367 = 0;
  assign exp_373 = exp_254 & exp_259;
  assign exp_434 = 0;

  reg [31:0] exp_414_reg;
  always@(*) begin
    case (exp_380)
      0:exp_414_reg <= exp_411;
      1:exp_414_reg <= exp_412;
      default:exp_414_reg <= exp_413;
    endcase
  end
  assign exp_414 = exp_414_reg;

      reg [0:0] exp_380_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_380_reg <= exp_372;
        end
      end
      assign exp_380 = exp_380_reg;
      assign exp_372 = exp_358 & exp_371;
  assign exp_358 = exp_345 & exp_357;
  assign exp_345 = exp_331 & exp_344;
  assign exp_331 = exp_329 & exp_330;
  assign exp_329 = exp_96[30:30];
  assign exp_330 = ~exp_294;
  assign exp_294 = exp_290 == exp_293;
  assign exp_293 = 19;
  assign exp_344 = ~exp_296;
  assign exp_357 = ~exp_298;
  assign exp_371 = ~exp_370;
  assign exp_370 = exp_300 | exp_302;
  assign exp_413 = 0;
  assign exp_411 = exp_376 + exp_377;

      reg [31:0] exp_376_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_376_reg <= exp_362;
        end
      end
      assign exp_376 = exp_376_reg;
    
  reg [31:0] exp_362_reg;
  always@(*) begin
    case (exp_359)
      0:exp_362_reg <= exp_351;
      1:exp_362_reg <= exp_360;
      default:exp_362_reg <= exp_361;
    endcase
  end
  assign exp_362 = exp_362_reg;
  assign exp_359 = exp_300 | exp_302;
  assign exp_361 = 0;

  reg [31:0] exp_351_reg;
  always@(*) begin
    case (exp_298)
      0:exp_351_reg <= exp_337;
      1:exp_351_reg <= exp_349;
      default:exp_351_reg <= exp_350;
    endcase
  end
  assign exp_351 = exp_351_reg;
  assign exp_350 = 0;

  reg [31:0] exp_337_reg;
  always@(*) begin
    case (exp_296)
      0:exp_337_reg <= exp_312;
      1:exp_337_reg <= exp_335;
      default:exp_337_reg <= exp_336;
    endcase
  end
  assign exp_337 = exp_337_reg;
  assign exp_336 = 0;
  assign exp_335 = exp_333 << exp_334;
  assign exp_333 = exp_332;
  assign exp_332 = exp_96[31:12];
  assign exp_334 = 12;
  assign exp_349 = exp_347 << exp_348;
  assign exp_347 = exp_346;
  assign exp_346 = exp_96[31:12];
  assign exp_348 = 12;
  assign exp_360 = 4;

      reg [31:0] exp_377_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_377_reg <= exp_365;
        end
      end
      assign exp_377 = exp_377_reg;
    
  reg [31:0] exp_365_reg;
  always@(*) begin
    case (exp_363)
      0:exp_365_reg <= exp_353;
      1:exp_365_reg <= exp_266;
      default:exp_365_reg <= exp_364;
    endcase
  end
  assign exp_365 = exp_365_reg;
  assign exp_363 = exp_300 | exp_302;
  assign exp_364 = 0;

  reg [31:0] exp_353_reg;
  always@(*) begin
    case (exp_298)
      0:exp_353_reg <= exp_340;
      1:exp_353_reg <= exp_266;
      default:exp_353_reg <= exp_352;
    endcase
  end
  assign exp_353 = exp_353_reg;
  assign exp_352 = 0;

  reg [31:0] exp_340_reg;
  always@(*) begin
    case (exp_296)
      0:exp_340_reg <= exp_324;
      1:exp_340_reg <= exp_338;
      default:exp_340_reg <= exp_339;
    endcase
  end
  assign exp_340 = exp_340_reg;
  assign exp_339 = 0;

  reg [31:0] exp_324_reg;
  always@(*) begin
    case (exp_294)
      0:exp_324_reg <= exp_318;
      1:exp_324_reg <= exp_322;
      default:exp_324_reg <= exp_323;
    endcase
  end
  assign exp_324 = exp_324_reg;
  assign exp_323 = 0;

  reg [31:0] exp_318_reg;
  always@(*) begin
    case (exp_314)
      0:exp_318_reg <= exp_306;
      1:exp_318_reg <= exp_316;
      default:exp_318_reg <= exp_317;
    endcase
  end
  assign exp_318 = exp_318_reg;
  assign exp_314 = exp_289 == exp_313;
  assign exp_289 = exp_96[24:20];
  assign exp_313 = 0;
  assign exp_317 = 0;

  reg [31:0] exp_306_reg;
  always@(*) begin
    case (exp_286)
      0:exp_306_reg <= exp_282;
      1:exp_306_reg <= exp_287;
      default:exp_306_reg <= exp_305;
    endcase
  end
  assign exp_306 = exp_306_reg;
  assign exp_286 = exp_862;
  assign exp_862 = exp_861 & exp_254;
  assign exp_861 = exp_860 & exp_262;
  assign exp_860 = exp_859 & exp_849;
  assign exp_859 = exp_268 == exp_850;
  assign exp_268 = exp_96[24:20];
  assign exp_305 = 0;

  //Create RAM
  reg [31:0] exp_282_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_280) begin
      exp_282_ram[exp_276] <= exp_278;
    end
  end
  assign exp_282 = exp_282_ram[exp_277];
  assign exp_281 = exp_284;
  assign exp_284 = 1;
  assign exp_277 = exp_268;
  assign exp_280 = exp_854;
  assign exp_854 = exp_853 & exp_254;
  assign exp_853 = exp_849 & exp_262;
  assign exp_276 = exp_850;
  assign exp_278 = exp_848;
  assign exp_287 = exp_848;
  assign exp_316 = $signed(exp_315);
  assign exp_315 = 0;
  assign exp_322 = exp_319 + exp_321;
  assign exp_319 = 0;
  assign exp_321 = $signed(exp_320);
  assign exp_320 = exp_96[31:20];
  assign exp_338 = 0;

      reg [31:0] exp_266_reg = 0;
      always@(posedge clk) begin
        if (exp_265) begin
          exp_266_reg <= exp_264;
        end
      end
      assign exp_266 = exp_266_reg;
      assign exp_265 = exp_256 & exp_254;
  assign exp_412 = exp_376 - exp_377;
  assign exp_416 = exp_376 << exp_415;
  assign exp_415 = $signed(exp_410);
  assign exp_410 = exp_409 + exp_408;
  assign exp_409 = 0;
  assign exp_408 = exp_379;

      reg [4:0] exp_379_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_379_reg <= exp_328;
        end
      end
      assign exp_379 = exp_379_reg;
    
  reg [4:0] exp_328_reg;
  always@(*) begin
    case (exp_294)
      0:exp_328_reg <= exp_326;
      1:exp_328_reg <= exp_291;
      default:exp_328_reg <= exp_327;
    endcase
  end
  assign exp_328 = exp_328_reg;
  assign exp_327 = 0;
  assign exp_326 = exp_324[4:0];
  assign exp_291 = exp_96[24:20];
  assign exp_432 = $signed(exp_418);
  assign exp_418 = exp_417;
  assign exp_417 = $signed(exp_376) < $signed(exp_377);
  assign exp_433 = $signed(exp_424);
  assign exp_424 = exp_423;
  assign exp_423 = exp_420 < exp_422;
  assign exp_420 = exp_419 + exp_376;
  assign exp_419 = 0;
  assign exp_422 = exp_421 + exp_377;
  assign exp_421 = 0;
  assign exp_425 = exp_376 ^ exp_377;
  assign exp_429 = exp_428[31:0];
  assign exp_428 = $signed(exp_426) >>> $signed(exp_427);
  assign exp_426 = {exp_407, exp_376};
  reg [0:0] exp_407_reg;
  always@(*) begin
    case (exp_381)
      0:exp_407_reg <= exp_405;
      1:exp_407_reg <= exp_404;
      default:exp_407_reg <= exp_406;
    endcase
  end
  assign exp_407 = exp_407_reg;

      reg [0:0] exp_381_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_381_reg <= exp_325;
        end
      end
      assign exp_381 = exp_381_reg;
      assign exp_325 = exp_96[30:30];
  assign exp_406 = 0;
  assign exp_405 = 0;
  assign exp_404 = exp_376[31:31];
  assign exp_427 = $signed(exp_410);
  assign exp_430 = exp_376 | exp_377;
  assign exp_431 = exp_376 & exp_377;

  reg [31:0] exp_482_reg;
  always@(*) begin
    case (exp_385)
      0:exp_482_reg <= exp_472;
      1:exp_482_reg <= exp_475;
      2:exp_482_reg <= exp_248;
      3:exp_482_reg <= exp_476;
      4:exp_482_reg <= exp_477;
      5:exp_482_reg <= exp_478;
      6:exp_482_reg <= exp_479;
      7:exp_482_reg <= exp_480;
      default:exp_482_reg <= exp_481;
    endcase
  end
  assign exp_482 = exp_482_reg;
  assign exp_481 = 0;
  assign exp_472 = $signed(exp_471);
  assign exp_471 = exp_470 + exp_465;
  assign exp_470 = 0;

  reg [7:0] exp_465_reg;
  always@(*) begin
    case (exp_456)
      0:exp_465_reg <= exp_460;
      1:exp_465_reg <= exp_461;
      2:exp_465_reg <= exp_462;
      3:exp_465_reg <= exp_463;
      default:exp_465_reg <= exp_464;
    endcase
  end
  assign exp_465 = exp_465_reg;
  assign exp_456 = exp_455 + exp_454;
  assign exp_455 = 0;
  assign exp_454 = exp_453[1:0];
  assign exp_464 = 0;
  assign exp_460 = exp_248[7:0];
  assign exp_248 = exp_238;

  reg [31:0] exp_238_reg;
  always@(*) begin
    case (exp_235)
      0:exp_238_reg <= exp_216;
      1:exp_238_reg <= exp_226;
      default:exp_238_reg <= exp_237;
    endcase
  end
  assign exp_238 = exp_238_reg;
  assign exp_237 = 0;

  reg [31:0] exp_216_reg;
  always@(*) begin
    case (exp_213)
      0:exp_216_reg <= exp_194;
      1:exp_216_reg <= exp_204;
      default:exp_216_reg <= exp_215;
    endcase
  end
  assign exp_216 = exp_216_reg;
  assign exp_215 = 0;

  reg [31:0] exp_194_reg;
  always@(*) begin
    case (exp_191)
      0:exp_194_reg <= exp_153;
      1:exp_194_reg <= exp_182;
      default:exp_194_reg <= exp_193;
    endcase
  end
  assign exp_194 = exp_194_reg;
  assign exp_193 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 0;
    exp_54_ram[32] = 255;
    exp_54_ram[33] = 39;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 0;
    exp_54_ram[36] = 0;
    exp_54_ram[37] = 0;
    exp_54_ram[38] = 0;
    exp_54_ram[39] = 0;
    exp_54_ram[40] = 40;
    exp_54_ram[41] = 113;
    exp_54_ram[42] = 14;
    exp_54_ram[43] = 0;
    exp_54_ram[44] = 12;
    exp_54_ram[45] = 15;
    exp_54_ram[46] = 0;
    exp_54_ram[47] = 0;
    exp_54_ram[48] = 0;
    exp_54_ram[49] = 0;
    exp_54_ram[50] = 0;
    exp_54_ram[51] = 2;
    exp_54_ram[52] = 0;
    exp_54_ram[53] = 64;
    exp_54_ram[54] = 0;
    exp_54_ram[55] = 0;
    exp_54_ram[56] = 0;
    exp_54_ram[57] = 0;
    exp_54_ram[58] = 0;
    exp_54_ram[59] = 0;
    exp_54_ram[60] = 1;
    exp_54_ram[61] = 3;
    exp_54_ram[62] = 1;
    exp_54_ram[63] = 1;
    exp_54_ram[64] = 1;
    exp_54_ram[65] = 3;
    exp_54_ram[66] = 0;
    exp_54_ram[67] = 2;
    exp_54_ram[68] = 1;
    exp_54_ram[69] = 0;
    exp_54_ram[70] = 0;
    exp_54_ram[71] = 1;
    exp_54_ram[72] = 255;
    exp_54_ram[73] = 1;
    exp_54_ram[74] = 0;
    exp_54_ram[75] = 255;
    exp_54_ram[76] = 1;
    exp_54_ram[77] = 64;
    exp_54_ram[78] = 3;
    exp_54_ram[79] = 1;
    exp_54_ram[80] = 1;
    exp_54_ram[81] = 3;
    exp_54_ram[82] = 1;
    exp_54_ram[83] = 0;
    exp_54_ram[84] = 2;
    exp_54_ram[85] = 0;
    exp_54_ram[86] = 0;
    exp_54_ram[87] = 0;
    exp_54_ram[88] = 255;
    exp_54_ram[89] = 1;
    exp_54_ram[90] = 0;
    exp_54_ram[91] = 255;
    exp_54_ram[92] = 1;
    exp_54_ram[93] = 0;
    exp_54_ram[94] = 0;
    exp_54_ram[95] = 14;
    exp_54_ram[96] = 1;
    exp_54_ram[97] = 1;
    exp_54_ram[98] = 242;
    exp_54_ram[99] = 1;
    exp_54_ram[100] = 243;
    exp_54_ram[101] = 0;
    exp_54_ram[102] = 0;
    exp_54_ram[103] = 2;
    exp_54_ram[104] = 0;
    exp_54_ram[105] = 12;
    exp_54_ram[106] = 15;
    exp_54_ram[107] = 1;
    exp_54_ram[108] = 0;
    exp_54_ram[109] = 0;
    exp_54_ram[110] = 0;
    exp_54_ram[111] = 0;
    exp_54_ram[112] = 2;
    exp_54_ram[113] = 0;
    exp_54_ram[114] = 64;
    exp_54_ram[115] = 10;
    exp_54_ram[116] = 65;
    exp_54_ram[117] = 0;
    exp_54_ram[118] = 1;
    exp_54_ram[119] = 1;
    exp_54_ram[120] = 1;
    exp_54_ram[121] = 1;
    exp_54_ram[122] = 3;
    exp_54_ram[123] = 3;
    exp_54_ram[124] = 1;
    exp_54_ram[125] = 0;
    exp_54_ram[126] = 2;
    exp_54_ram[127] = 0;
    exp_54_ram[128] = 1;
    exp_54_ram[129] = 1;
    exp_54_ram[130] = 255;
    exp_54_ram[131] = 1;
    exp_54_ram[132] = 1;
    exp_54_ram[133] = 255;
    exp_54_ram[134] = 1;
    exp_54_ram[135] = 65;
    exp_54_ram[136] = 3;
    exp_54_ram[137] = 1;
    exp_54_ram[138] = 1;
    exp_54_ram[139] = 3;
    exp_54_ram[140] = 1;
    exp_54_ram[141] = 0;
    exp_54_ram[142] = 2;
    exp_54_ram[143] = 0;
    exp_54_ram[144] = 0;
    exp_54_ram[145] = 0;
    exp_54_ram[146] = 255;
    exp_54_ram[147] = 1;
    exp_54_ram[148] = 0;
    exp_54_ram[149] = 255;
    exp_54_ram[150] = 1;
    exp_54_ram[151] = 0;
    exp_54_ram[152] = 0;
    exp_54_ram[153] = 1;
    exp_54_ram[154] = 1;
    exp_54_ram[155] = 244;
    exp_54_ram[156] = 1;
    exp_54_ram[157] = 244;
    exp_54_ram[158] = 0;
    exp_54_ram[159] = 0;
    exp_54_ram[160] = 0;
    exp_54_ram[161] = 0;
    exp_54_ram[162] = 0;
    exp_54_ram[163] = 1;
    exp_54_ram[164] = 0;
    exp_54_ram[165] = 3;
    exp_54_ram[166] = 1;
    exp_54_ram[167] = 1;
    exp_54_ram[168] = 1;
    exp_54_ram[169] = 3;
    exp_54_ram[170] = 1;
    exp_54_ram[171] = 0;
    exp_54_ram[172] = 2;
    exp_54_ram[173] = 0;
    exp_54_ram[174] = 0;
    exp_54_ram[175] = 1;
    exp_54_ram[176] = 255;
    exp_54_ram[177] = 1;
    exp_54_ram[178] = 0;
    exp_54_ram[179] = 255;
    exp_54_ram[180] = 1;
    exp_54_ram[181] = 64;
    exp_54_ram[182] = 3;
    exp_54_ram[183] = 1;
    exp_54_ram[184] = 1;
    exp_54_ram[185] = 3;
    exp_54_ram[186] = 1;
    exp_54_ram[187] = 2;
    exp_54_ram[188] = 0;
    exp_54_ram[189] = 0;
    exp_54_ram[190] = 0;
    exp_54_ram[191] = 1;
    exp_54_ram[192] = 255;
    exp_54_ram[193] = 1;
    exp_54_ram[194] = 0;
    exp_54_ram[195] = 255;
    exp_54_ram[196] = 1;
    exp_54_ram[197] = 1;
    exp_54_ram[198] = 64;
    exp_54_ram[199] = 0;
    exp_54_ram[200] = 235;
    exp_54_ram[201] = 24;
    exp_54_ram[202] = 0;
    exp_54_ram[203] = 4;
    exp_54_ram[204] = 15;
    exp_54_ram[205] = 0;
    exp_54_ram[206] = 0;
    exp_54_ram[207] = 0;
    exp_54_ram[208] = 113;
    exp_54_ram[209] = 0;
    exp_54_ram[210] = 0;
    exp_54_ram[211] = 2;
    exp_54_ram[212] = 0;
    exp_54_ram[213] = 64;
    exp_54_ram[214] = 2;
    exp_54_ram[215] = 0;
    exp_54_ram[216] = 240;
    exp_54_ram[217] = 0;
    exp_54_ram[218] = 0;
    exp_54_ram[219] = 239;
    exp_54_ram[220] = 1;
    exp_54_ram[221] = 1;
    exp_54_ram[222] = 252;
    exp_54_ram[223] = 1;
    exp_54_ram[224] = 251;
    exp_54_ram[225] = 0;
    exp_54_ram[226] = 0;
    exp_54_ram[227] = 0;
    exp_54_ram[228] = 0;
    exp_54_ram[229] = 1;
    exp_54_ram[230] = 3;
    exp_54_ram[231] = 0;
    exp_54_ram[232] = 0;
    exp_54_ram[233] = 0;
    exp_54_ram[234] = 0;
    exp_54_ram[235] = 1;
    exp_54_ram[236] = 1;
    exp_54_ram[237] = 1;
    exp_54_ram[238] = 3;
    exp_54_ram[239] = 1;
    exp_54_ram[240] = 0;
    exp_54_ram[241] = 3;
    exp_54_ram[242] = 0;
    exp_54_ram[243] = 1;
    exp_54_ram[244] = 1;
    exp_54_ram[245] = 255;
    exp_54_ram[246] = 1;
    exp_54_ram[247] = 1;
    exp_54_ram[248] = 255;
    exp_54_ram[249] = 1;
    exp_54_ram[250] = 65;
    exp_54_ram[251] = 3;
    exp_54_ram[252] = 3;
    exp_54_ram[253] = 1;
    exp_54_ram[254] = 2;
    exp_54_ram[255] = 1;
    exp_54_ram[256] = 1;
    exp_54_ram[257] = 0;
    exp_54_ram[258] = 0;
    exp_54_ram[259] = 1;
    exp_54_ram[260] = 1;
    exp_54_ram[261] = 255;
    exp_54_ram[262] = 1;
    exp_54_ram[263] = 1;
    exp_54_ram[264] = 255;
    exp_54_ram[265] = 1;
    exp_54_ram[266] = 1;
    exp_54_ram[267] = 0;
    exp_54_ram[268] = 0;
    exp_54_ram[269] = 255;
    exp_54_ram[270] = 0;
    exp_54_ram[271] = 1;
    exp_54_ram[272] = 0;
    exp_54_ram[273] = 1;
    exp_54_ram[274] = 65;
    exp_54_ram[275] = 2;
    exp_54_ram[276] = 2;
    exp_54_ram[277] = 1;
    exp_54_ram[278] = 2;
    exp_54_ram[279] = 0;
    exp_54_ram[280] = 1;
    exp_54_ram[281] = 2;
    exp_54_ram[282] = 0;
    exp_54_ram[283] = 1;
    exp_54_ram[284] = 1;
    exp_54_ram[285] = 0;
    exp_54_ram[286] = 2;
    exp_54_ram[287] = 206;
    exp_54_ram[288] = 0;
    exp_54_ram[289] = 255;
    exp_54_ram[290] = 0;
    exp_54_ram[291] = 1;
    exp_54_ram[292] = 0;
    exp_54_ram[293] = 0;
    exp_54_ram[294] = 1;
    exp_54_ram[295] = 0;
    exp_54_ram[296] = 220;
    exp_54_ram[297] = 255;
    exp_54_ram[298] = 205;
    exp_54_ram[299] = 0;
    exp_54_ram[300] = 0;
    exp_54_ram[301] = 218;
    exp_54_ram[302] = 0;
    exp_54_ram[303] = 0;
    exp_54_ram[304] = 0;
    exp_54_ram[305] = 0;
    exp_54_ram[306] = 0;
    exp_54_ram[307] = 0;
    exp_54_ram[308] = 0;
    exp_54_ram[309] = 254;
    exp_54_ram[310] = 0;
    exp_54_ram[311] = 6;
    exp_54_ram[312] = 6;
    exp_54_ram[313] = 0;
    exp_54_ram[314] = 0;
    exp_54_ram[315] = 255;
    exp_54_ram[316] = 2;
    exp_54_ram[317] = 0;
    exp_54_ram[318] = 0;
    exp_54_ram[319] = 0;
    exp_54_ram[320] = 0;
    exp_54_ram[321] = 0;
    exp_54_ram[322] = 254;
    exp_54_ram[323] = 0;
    exp_54_ram[324] = 0;
    exp_54_ram[325] = 64;
    exp_54_ram[326] = 0;
    exp_54_ram[327] = 0;
    exp_54_ram[328] = 0;
    exp_54_ram[329] = 254;
    exp_54_ram[330] = 0;
    exp_54_ram[331] = 0;
    exp_54_ram[332] = 251;
    exp_54_ram[333] = 0;
    exp_54_ram[334] = 0;
    exp_54_ram[335] = 64;
    exp_54_ram[336] = 0;
    exp_54_ram[337] = 64;
    exp_54_ram[338] = 249;
    exp_54_ram[339] = 64;
    exp_54_ram[340] = 0;
    exp_54_ram[341] = 249;
    exp_54_ram[342] = 64;
    exp_54_ram[343] = 0;
    exp_54_ram[344] = 0;
    exp_54_ram[345] = 0;
    exp_54_ram[346] = 0;
    exp_54_ram[347] = 247;
    exp_54_ram[348] = 0;
    exp_54_ram[349] = 0;
    exp_54_ram[350] = 64;
    exp_54_ram[351] = 254;
    exp_54_ram[352] = 64;
    exp_54_ram[353] = 246;
    exp_54_ram[354] = 64;
    exp_54_ram[355] = 0;
    exp_54_ram[356] = 108;
    exp_54_ram[357] = 111;
    exp_54_ram[358] = 33;
    exp_54_ram[359] = 0;
    exp_54_ram[360] = 110;
    exp_54_ram[361] = 32;
    exp_54_ram[362] = 103;
    exp_54_ram[363] = 114;
    exp_54_ram[364] = 114;
    exp_54_ram[365] = 109;
    exp_54_ram[366] = 46;
    exp_54_ram[367] = 0;
    exp_54_ram[368] = 0;
    exp_54_ram[369] = 51;
    exp_54_ram[370] = 105;
    exp_54_ram[371] = 110;
    exp_54_ram[372] = 101;
    exp_54_ram[373] = 117;
    exp_54_ram[374] = 112;
    exp_54_ram[375] = 115;
    exp_54_ram[376] = 32;
    exp_54_ram[377] = 101;
    exp_54_ram[378] = 100;
    exp_54_ram[379] = 0;
    exp_54_ram[380] = 54;
    exp_54_ram[381] = 105;
    exp_54_ram[382] = 110;
    exp_54_ram[383] = 101;
    exp_54_ram[384] = 117;
    exp_54_ram[385] = 112;
    exp_54_ram[386] = 115;
    exp_54_ram[387] = 32;
    exp_54_ram[388] = 101;
    exp_54_ram[389] = 100;
    exp_54_ram[390] = 0;
    exp_54_ram[391] = 51;
    exp_54_ram[392] = 105;
    exp_54_ram[393] = 110;
    exp_54_ram[394] = 101;
    exp_54_ram[395] = 105;
    exp_54_ram[396] = 101;
    exp_54_ram[397] = 110;
    exp_54_ram[398] = 115;
    exp_54_ram[399] = 110;
    exp_54_ram[400] = 0;
    exp_54_ram[401] = 54;
    exp_54_ram[402] = 105;
    exp_54_ram[403] = 110;
    exp_54_ram[404] = 101;
    exp_54_ram[405] = 105;
    exp_54_ram[406] = 101;
    exp_54_ram[407] = 110;
    exp_54_ram[408] = 115;
    exp_54_ram[409] = 110;
    exp_54_ram[410] = 0;
    exp_54_ram[411] = 103;
    exp_54_ram[412] = 110;
    exp_54_ram[413] = 117;
    exp_54_ram[414] = 0;
    exp_54_ram[415] = 108;
    exp_54_ram[416] = 0;
    exp_54_ram[417] = 115;
    exp_54_ram[418] = 0;
    exp_54_ram[419] = 111;
    exp_54_ram[420] = 101;
    exp_54_ram[421] = 48;
    exp_54_ram[422] = 37;
    exp_54_ram[423] = 32;
    exp_54_ram[424] = 120;
    exp_54_ram[425] = 0;
    exp_54_ram[426] = 105;
    exp_54_ram[427] = 86;
    exp_54_ram[428] = 109;
    exp_54_ram[429] = 0;
    exp_54_ram[430] = 32;
    exp_54_ram[431] = 108;
    exp_54_ram[432] = 111;
    exp_54_ram[433] = 0;
    exp_54_ram[434] = 75;
    exp_54_ram[435] = 104;
    exp_54_ram[436] = 105;
    exp_54_ram[437] = 0;
    exp_54_ram[438] = 83;
    exp_54_ram[439] = 32;
    exp_54_ram[440] = 99;
    exp_54_ram[441] = 0;
    exp_54_ram[442] = 84;
    exp_54_ram[443] = 32;
    exp_54_ram[444] = 116;
    exp_54_ram[445] = 105;
    exp_54_ram[446] = 105;
    exp_54_ram[447] = 0;
    exp_54_ram[448] = 84;
    exp_54_ram[449] = 32;
    exp_54_ram[450] = 111;
    exp_54_ram[451] = 0;
    exp_54_ram[452] = 2;
    exp_54_ram[453] = 3;
    exp_54_ram[454] = 4;
    exp_54_ram[455] = 4;
    exp_54_ram[456] = 5;
    exp_54_ram[457] = 5;
    exp_54_ram[458] = 5;
    exp_54_ram[459] = 5;
    exp_54_ram[460] = 6;
    exp_54_ram[461] = 6;
    exp_54_ram[462] = 6;
    exp_54_ram[463] = 6;
    exp_54_ram[464] = 6;
    exp_54_ram[465] = 6;
    exp_54_ram[466] = 6;
    exp_54_ram[467] = 6;
    exp_54_ram[468] = 7;
    exp_54_ram[469] = 7;
    exp_54_ram[470] = 7;
    exp_54_ram[471] = 7;
    exp_54_ram[472] = 7;
    exp_54_ram[473] = 7;
    exp_54_ram[474] = 7;
    exp_54_ram[475] = 7;
    exp_54_ram[476] = 7;
    exp_54_ram[477] = 7;
    exp_54_ram[478] = 7;
    exp_54_ram[479] = 7;
    exp_54_ram[480] = 7;
    exp_54_ram[481] = 7;
    exp_54_ram[482] = 7;
    exp_54_ram[483] = 7;
    exp_54_ram[484] = 8;
    exp_54_ram[485] = 8;
    exp_54_ram[486] = 8;
    exp_54_ram[487] = 8;
    exp_54_ram[488] = 8;
    exp_54_ram[489] = 8;
    exp_54_ram[490] = 8;
    exp_54_ram[491] = 8;
    exp_54_ram[492] = 8;
    exp_54_ram[493] = 8;
    exp_54_ram[494] = 8;
    exp_54_ram[495] = 8;
    exp_54_ram[496] = 8;
    exp_54_ram[497] = 8;
    exp_54_ram[498] = 8;
    exp_54_ram[499] = 8;
    exp_54_ram[500] = 8;
    exp_54_ram[501] = 8;
    exp_54_ram[502] = 8;
    exp_54_ram[503] = 8;
    exp_54_ram[504] = 8;
    exp_54_ram[505] = 8;
    exp_54_ram[506] = 8;
    exp_54_ram[507] = 8;
    exp_54_ram[508] = 8;
    exp_54_ram[509] = 8;
    exp_54_ram[510] = 8;
    exp_54_ram[511] = 8;
    exp_54_ram[512] = 8;
    exp_54_ram[513] = 8;
    exp_54_ram[514] = 8;
    exp_54_ram[515] = 8;
    exp_54_ram[516] = 0;
    exp_54_ram[517] = 0;
    exp_54_ram[518] = 0;
    exp_54_ram[519] = 62;
    exp_54_ram[520] = 0;
    exp_54_ram[521] = 0;
    exp_54_ram[522] = 0;
    exp_54_ram[523] = 0;
    exp_54_ram[524] = 0;
    exp_54_ram[525] = 0;
    exp_54_ram[526] = 0;
    exp_54_ram[527] = 0;
    exp_54_ram[528] = 0;
    exp_54_ram[529] = 0;
    exp_54_ram[530] = 254;
    exp_54_ram[531] = 255;
    exp_54_ram[532] = 0;
    exp_54_ram[533] = 0;
    exp_54_ram[534] = 61;
    exp_54_ram[535] = 0;
    exp_54_ram[536] = 0;
    exp_54_ram[537] = 252;
    exp_54_ram[538] = 0;
    exp_54_ram[539] = 0;
    exp_54_ram[540] = 0;
    exp_54_ram[541] = 0;
    exp_54_ram[542] = 0;
    exp_54_ram[543] = 1;
    exp_54_ram[544] = 0;
    exp_54_ram[545] = 255;
    exp_54_ram[546] = 0;
    exp_54_ram[547] = 0;
    exp_54_ram[548] = 0;
    exp_54_ram[549] = 0;
    exp_54_ram[550] = 247;
    exp_54_ram[551] = 0;
    exp_54_ram[552] = 0;
    exp_54_ram[553] = 0;
    exp_54_ram[554] = 1;
    exp_54_ram[555] = 0;
    exp_54_ram[556] = 0;
    exp_54_ram[557] = 0;
    exp_54_ram[558] = 0;
    exp_54_ram[559] = 0;
    exp_54_ram[560] = 253;
    exp_54_ram[561] = 252;
    exp_54_ram[562] = 2;
    exp_54_ram[563] = 2;
    exp_54_ram[564] = 3;
    exp_54_ram[565] = 3;
    exp_54_ram[566] = 3;
    exp_54_ram[567] = 1;
    exp_54_ram[568] = 1;
    exp_54_ram[569] = 0;
    exp_54_ram[570] = 2;
    exp_54_ram[571] = 3;
    exp_54_ram[572] = 3;
    exp_54_ram[573] = 1;
    exp_54_ram[574] = 1;
    exp_54_ram[575] = 1;
    exp_54_ram[576] = 0;
    exp_54_ram[577] = 0;
    exp_54_ram[578] = 0;
    exp_54_ram[579] = 0;
    exp_54_ram[580] = 0;
    exp_54_ram[581] = 0;
    exp_54_ram[582] = 0;
    exp_54_ram[583] = 0;
    exp_54_ram[584] = 14;
    exp_54_ram[585] = 1;
    exp_54_ram[586] = 14;
    exp_54_ram[587] = 0;
    exp_54_ram[588] = 16;
    exp_54_ram[589] = 0;
    exp_54_ram[590] = 0;
    exp_54_ram[591] = 0;
    exp_54_ram[592] = 0;
    exp_54_ram[593] = 0;
    exp_54_ram[594] = 3;
    exp_54_ram[595] = 15;
    exp_54_ram[596] = 0;
    exp_54_ram[597] = 0;
    exp_54_ram[598] = 9;
    exp_54_ram[599] = 15;
    exp_54_ram[600] = 6;
    exp_54_ram[601] = 3;
    exp_54_ram[602] = 15;
    exp_54_ram[603] = 0;
    exp_54_ram[604] = 0;
    exp_54_ram[605] = 0;
    exp_54_ram[606] = 0;
    exp_54_ram[607] = 240;
    exp_54_ram[608] = 0;
    exp_54_ram[609] = 3;
    exp_54_ram[610] = 255;
    exp_54_ram[611] = 3;
    exp_54_ram[612] = 251;
    exp_54_ram[613] = 3;
    exp_54_ram[614] = 3;
    exp_54_ram[615] = 3;
    exp_54_ram[616] = 3;
    exp_54_ram[617] = 2;
    exp_54_ram[618] = 2;
    exp_54_ram[619] = 2;
    exp_54_ram[620] = 2;
    exp_54_ram[621] = 1;
    exp_54_ram[622] = 1;
    exp_54_ram[623] = 1;
    exp_54_ram[624] = 1;
    exp_54_ram[625] = 0;
    exp_54_ram[626] = 4;
    exp_54_ram[627] = 0;
    exp_54_ram[628] = 0;
    exp_54_ram[629] = 3;
    exp_54_ram[630] = 249;
    exp_54_ram[631] = 5;
    exp_54_ram[632] = 248;
    exp_54_ram[633] = 251;
    exp_54_ram[634] = 0;
    exp_54_ram[635] = 0;
    exp_54_ram[636] = 0;
    exp_54_ram[637] = 0;
    exp_54_ram[638] = 232;
    exp_54_ram[639] = 248;
    exp_54_ram[640] = 0;
    exp_54_ram[641] = 8;
    exp_54_ram[642] = 242;
    exp_54_ram[643] = 59;
    exp_54_ram[644] = 0;
    exp_54_ram[645] = 160;
    exp_54_ram[646] = 0;
    exp_54_ram[647] = 241;
    exp_54_ram[648] = 0;
    exp_54_ram[649] = 40;
    exp_54_ram[650] = 251;
    exp_54_ram[651] = 4;
    exp_54_ram[652] = 4;
    exp_54_ram[653] = 3;
    exp_54_ram[654] = 3;
    exp_54_ram[655] = 3;
    exp_54_ram[656] = 3;
    exp_54_ram[657] = 3;
    exp_54_ram[658] = 3;
    exp_54_ram[659] = 1;
    exp_54_ram[660] = 0;
    exp_54_ram[661] = 4;
    exp_54_ram[662] = 5;
    exp_54_ram[663] = 3;
    exp_54_ram[664] = 3;
    exp_54_ram[665] = 0;
    exp_54_ram[666] = 0;
    exp_54_ram[667] = 0;
    exp_54_ram[668] = 0;
    exp_54_ram[669] = 0;
    exp_54_ram[670] = 2;
    exp_54_ram[671] = 0;
    exp_54_ram[672] = 0;
    exp_54_ram[673] = 6;
    exp_54_ram[674] = 7;
    exp_54_ram[675] = 0;
    exp_54_ram[676] = 0;
    exp_54_ram[677] = 0;
    exp_54_ram[678] = 1;
    exp_54_ram[679] = 7;
    exp_54_ram[680] = 0;
    exp_54_ram[681] = 0;
    exp_54_ram[682] = 3;
    exp_54_ram[683] = 6;
    exp_54_ram[684] = 0;
    exp_54_ram[685] = 1;
    exp_54_ram[686] = 0;
    exp_54_ram[687] = 6;
    exp_54_ram[688] = 4;
    exp_54_ram[689] = 4;
    exp_54_ram[690] = 4;
    exp_54_ram[691] = 4;
    exp_54_ram[692] = 3;
    exp_54_ram[693] = 3;
    exp_54_ram[694] = 3;
    exp_54_ram[695] = 3;
    exp_54_ram[696] = 2;
    exp_54_ram[697] = 2;
    exp_54_ram[698] = 2;
    exp_54_ram[699] = 2;
    exp_54_ram[700] = 1;
    exp_54_ram[701] = 0;
    exp_54_ram[702] = 5;
    exp_54_ram[703] = 0;
    exp_54_ram[704] = 0;
    exp_54_ram[705] = 0;
    exp_54_ram[706] = 0;
    exp_54_ram[707] = 215;
    exp_54_ram[708] = 0;
    exp_54_ram[709] = 0;
    exp_54_ram[710] = 250;
    exp_54_ram[711] = 0;
    exp_54_ram[712] = 246;
    exp_54_ram[713] = 2;
    exp_54_ram[714] = 0;
    exp_54_ram[715] = 1;
    exp_54_ram[716] = 0;
    exp_54_ram[717] = 0;
    exp_54_ram[718] = 1;
    exp_54_ram[719] = 253;
    exp_54_ram[720] = 2;
    exp_54_ram[721] = 5;
    exp_54_ram[722] = 8;
    exp_54_ram[723] = 6;
    exp_54_ram[724] = 14;
    exp_54_ram[725] = 2;
    exp_54_ram[726] = 13;
    exp_54_ram[727] = 5;
    exp_54_ram[728] = 250;
    exp_54_ram[729] = 0;
    exp_54_ram[730] = 0;
    exp_54_ram[731] = 11;
    exp_54_ram[732] = 3;
    exp_54_ram[733] = 0;
    exp_54_ram[734] = 0;
    exp_54_ram[735] = 250;
    exp_54_ram[736] = 244;
    exp_54_ram[737] = 6;
    exp_54_ram[738] = 248;
    exp_54_ram[739] = 0;
    exp_54_ram[740] = 0;
    exp_54_ram[741] = 14;
    exp_54_ram[742] = 0;
    exp_54_ram[743] = 0;
    exp_54_ram[744] = 0;
    exp_54_ram[745] = 2;
    exp_54_ram[746] = 0;
    exp_54_ram[747] = 0;
    exp_54_ram[748] = 205;
    exp_54_ram[749] = 0;
    exp_54_ram[750] = 0;
    exp_54_ram[751] = 0;
    exp_54_ram[752] = 0;
    exp_54_ram[753] = 0;
    exp_54_ram[754] = 255;
    exp_54_ram[755] = 65;
    exp_54_ram[756] = 0;
    exp_54_ram[757] = 0;
    exp_54_ram[758] = 206;
    exp_54_ram[759] = 7;
    exp_54_ram[760] = 11;
    exp_54_ram[761] = 2;
    exp_54_ram[762] = 6;
    exp_54_ram[763] = 10;
    exp_54_ram[764] = 7;
    exp_54_ram[765] = 242;
    exp_54_ram[766] = 0;
    exp_54_ram[767] = 0;
    exp_54_ram[768] = 0;
    exp_54_ram[769] = 4;
    exp_54_ram[770] = 0;
    exp_54_ram[771] = 240;
    exp_54_ram[772] = 7;
    exp_54_ram[773] = 240;
    exp_54_ram[774] = 0;
    exp_54_ram[775] = 0;
    exp_54_ram[776] = 1;
    exp_54_ram[777] = 7;
    exp_54_ram[778] = 0;
    exp_54_ram[779] = 0;
    exp_54_ram[780] = 0;
    exp_54_ram[781] = 2;
    exp_54_ram[782] = 237;
    exp_54_ram[783] = 0;
    exp_54_ram[784] = 0;
    exp_54_ram[785] = 0;
    exp_54_ram[786] = 0;
    exp_54_ram[787] = 0;
    exp_54_ram[788] = 195;
    exp_54_ram[789] = 0;
    exp_54_ram[790] = 0;
    exp_54_ram[791] = 235;
    exp_54_ram[792] = 0;
    exp_54_ram[793] = 0;
    exp_54_ram[794] = 0;
    exp_54_ram[795] = 0;
    exp_54_ram[796] = 193;
    exp_54_ram[797] = 0;
    exp_54_ram[798] = 0;
    exp_54_ram[799] = 0;
    exp_54_ram[800] = 248;
    exp_54_ram[801] = 0;
    exp_54_ram[802] = 0;
    exp_54_ram[803] = 0;
    exp_54_ram[804] = 244;
    exp_54_ram[805] = 0;
    exp_54_ram[806] = 0;
    exp_54_ram[807] = 0;
    exp_54_ram[808] = 0;
    exp_54_ram[809] = 242;
    exp_54_ram[810] = 0;
    exp_54_ram[811] = 0;
    exp_54_ram[812] = 0;
    exp_54_ram[813] = 254;
    exp_54_ram[814] = 0;
    exp_54_ram[815] = 0;
    exp_54_ram[816] = 0;
    exp_54_ram[817] = 252;
    exp_54_ram[818] = 2;
    exp_54_ram[819] = 0;
    exp_54_ram[820] = 2;
    exp_54_ram[821] = 0;
    exp_54_ram[822] = 61;
    exp_54_ram[823] = 2;
    exp_54_ram[824] = 2;
    exp_54_ram[825] = 0;
    exp_54_ram[826] = 2;
    exp_54_ram[827] = 0;
    exp_54_ram[828] = 2;
    exp_54_ram[829] = 3;
    exp_54_ram[830] = 3;
    exp_54_ram[831] = 0;
    exp_54_ram[832] = 210;
    exp_54_ram[833] = 1;
    exp_54_ram[834] = 4;
    exp_54_ram[835] = 0;
    exp_54_ram[836] = 0;
    exp_54_ram[837] = 0;
    exp_54_ram[838] = 0;
    exp_54_ram[839] = 67;
    exp_54_ram[840] = 0;
    exp_54_ram[841] = 0;
    exp_54_ram[842] = 0;
    exp_54_ram[843] = 0;
    exp_54_ram[844] = 0;
    exp_54_ram[845] = 0;
    exp_54_ram[846] = 61;
    exp_54_ram[847] = 0;
    exp_54_ram[848] = 0;
    exp_54_ram[849] = 255;
    exp_54_ram[850] = 0;
    exp_54_ram[851] = 0;
    exp_54_ram[852] = 0;
    exp_54_ram[853] = 255;
    exp_54_ram[854] = 0;
    exp_54_ram[855] = 252;
    exp_54_ram[856] = 0;
    exp_54_ram[857] = 0;
    exp_54_ram[858] = 0;
    exp_54_ram[859] = 1;
    exp_54_ram[860] = 0;
    exp_54_ram[861] = 0;
    exp_54_ram[862] = 0;
    exp_54_ram[863] = 0;
    exp_54_ram[864] = 0;
    exp_54_ram[865] = 253;
    exp_54_ram[866] = 0;
    exp_54_ram[867] = 0;
    exp_54_ram[868] = 2;
    exp_54_ram[869] = 0;
    exp_54_ram[870] = 0;
    exp_54_ram[871] = 0;
    exp_54_ram[872] = 255;
    exp_54_ram[873] = 0;
    exp_54_ram[874] = 0;
    exp_54_ram[875] = 0;
    exp_54_ram[876] = 0;
    exp_54_ram[877] = 247;
    exp_54_ram[878] = 0;
    exp_54_ram[879] = 67;
    exp_54_ram[880] = 64;
    exp_54_ram[881] = 255;
    exp_54_ram[882] = 255;
    exp_54_ram[883] = 0;
    exp_54_ram[884] = 0;
    exp_54_ram[885] = 0;
    exp_54_ram[886] = 255;
    exp_54_ram[887] = 0;
    exp_54_ram[888] = 0;
    exp_54_ram[889] = 0;
    exp_54_ram[890] = 61;
    exp_54_ram[891] = 67;
    exp_54_ram[892] = 0;
    exp_54_ram[893] = 0;
    exp_54_ram[894] = 0;
    exp_54_ram[895] = 7;
    exp_54_ram[896] = 0;
    exp_54_ram[897] = 0;
    exp_54_ram[898] = 0;
    exp_54_ram[899] = 0;
    exp_54_ram[900] = 0;
    exp_54_ram[901] = 0;
    exp_54_ram[902] = 0;
    exp_54_ram[903] = 252;
    exp_54_ram[904] = 0;
    exp_54_ram[905] = 0;
    exp_54_ram[906] = 3;
    exp_54_ram[907] = 0;
    exp_54_ram[908] = 0;
    exp_54_ram[909] = 0;
    exp_54_ram[910] = 0;
    exp_54_ram[911] = 0;
    exp_54_ram[912] = 250;
    exp_54_ram[913] = 0;
    exp_54_ram[914] = 0;
    exp_54_ram[915] = 0;
    exp_54_ram[916] = 0;
    exp_54_ram[917] = 0;
    exp_54_ram[918] = 253;
    exp_54_ram[919] = 0;
    exp_54_ram[920] = 0;
    exp_54_ram[921] = 0;
    exp_54_ram[922] = 0;
    exp_54_ram[923] = 6;
    exp_54_ram[924] = 0;
    exp_54_ram[925] = 0;
    exp_54_ram[926] = 0;
    exp_54_ram[927] = 2;
    exp_54_ram[928] = 0;
    exp_54_ram[929] = 1;
    exp_54_ram[930] = 1;
    exp_54_ram[931] = 255;
    exp_54_ram[932] = 255;
    exp_54_ram[933] = 255;
    exp_54_ram[934] = 255;
    exp_54_ram[935] = 255;
    exp_54_ram[936] = 255;
    exp_54_ram[937] = 255;
    exp_54_ram[938] = 64;
    exp_54_ram[939] = 253;
    exp_54_ram[940] = 0;
    exp_54_ram[941] = 255;
    exp_54_ram[942] = 0;
    exp_54_ram[943] = 0;
    exp_54_ram[944] = 0;
    exp_54_ram[945] = 64;
    exp_54_ram[946] = 3;
    exp_54_ram[947] = 0;
    exp_54_ram[948] = 0;
    exp_54_ram[949] = 0;
    exp_54_ram[950] = 0;
    exp_54_ram[951] = 0;
    exp_54_ram[952] = 2;
    exp_54_ram[953] = 0;
    exp_54_ram[954] = 0;
    exp_54_ram[955] = 0;
    exp_54_ram[956] = 0;
    exp_54_ram[957] = 0;
    exp_54_ram[958] = 1;
    exp_54_ram[959] = 252;
    exp_54_ram[960] = 0;
    exp_54_ram[961] = 0;
    exp_54_ram[962] = 0;
    exp_54_ram[963] = 0;
    exp_54_ram[964] = 1;
    exp_54_ram[965] = 252;
    exp_54_ram[966] = 0;
    exp_54_ram[967] = 4;
    exp_54_ram[968] = 255;
    exp_54_ram[969] = 6;
    exp_54_ram[970] = 0;
    exp_54_ram[971] = 0;
    exp_54_ram[972] = 0;
    exp_54_ram[973] = 223;
    exp_54_ram[974] = 0;
    exp_54_ram[975] = 0;
    exp_54_ram[976] = 25;
    exp_54_ram[977] = 0;
    exp_54_ram[978] = 222;
    exp_54_ram[979] = 0;
    exp_54_ram[980] = 0;
    exp_54_ram[981] = 0;
    exp_54_ram[982] = 0;
    exp_54_ram[983] = 1;
    exp_54_ram[984] = 0;
    exp_54_ram[985] = 0;
    exp_54_ram[986] = 0;
    exp_54_ram[987] = 0;
    exp_54_ram[988] = 255;
    exp_54_ram[989] = 255;
    exp_54_ram[990] = 4;
    exp_54_ram[991] = 255;
    exp_54_ram[992] = 0;
    exp_54_ram[993] = 1;
    exp_54_ram[994] = 2;
    exp_54_ram[995] = 0;
    exp_54_ram[996] = 1;
    exp_54_ram[997] = 2;
    exp_54_ram[998] = 255;
    exp_54_ram[999] = 0;
    exp_54_ram[1000] = 247;
    exp_54_ram[1001] = 0;
    exp_54_ram[1002] = 0;
    exp_54_ram[1003] = 1;
    exp_54_ram[1004] = 0;
    exp_54_ram[1005] = 1;
    exp_54_ram[1006] = 0;
    exp_54_ram[1007] = 1;
    exp_54_ram[1008] = 0;
    exp_54_ram[1009] = 0;
    exp_54_ram[1010] = 128;
    exp_54_ram[1011] = 0;
    exp_54_ram[1012] = 0;
    exp_54_ram[1013] = 0;
    exp_54_ram[1014] = 0;
    exp_54_ram[1015] = 0;
    exp_54_ram[1016] = 0;
    exp_54_ram[1017] = 0;
    exp_54_ram[1018] = 254;
    exp_54_ram[1019] = 1;
    exp_54_ram[1020] = 1;
    exp_54_ram[1021] = 0;
    exp_54_ram[1022] = 0;
    exp_54_ram[1023] = 0;
    exp_54_ram[1024] = 1;
    exp_54_ram[1025] = 1;
    exp_54_ram[1026] = 1;
    exp_54_ram[1027] = 0;
    exp_54_ram[1028] = 1;
    exp_54_ram[1029] = 0;
    exp_54_ram[1030] = 123;
    exp_54_ram[1031] = 0;
    exp_54_ram[1032] = 0;
    exp_54_ram[1033] = 118;
    exp_54_ram[1034] = 24;
    exp_54_ram[1035] = 4;
    exp_54_ram[1036] = 1;
    exp_54_ram[1037] = 0;
    exp_54_ram[1038] = 0;
    exp_54_ram[1039] = 24;
    exp_54_ram[1040] = 6;
    exp_54_ram[1041] = 0;
    exp_54_ram[1042] = 0;
    exp_54_ram[1043] = 242;
    exp_54_ram[1044] = 0;
    exp_54_ram[1045] = 198;
    exp_54_ram[1046] = 0;
    exp_54_ram[1047] = 1;
    exp_54_ram[1048] = 1;
    exp_54_ram[1049] = 0;
    exp_54_ram[1050] = 0;
    exp_54_ram[1051] = 253;
    exp_54_ram[1052] = 0;
    exp_54_ram[1053] = 234;
    exp_54_ram[1054] = 0;
    exp_54_ram[1055] = 0;
    exp_54_ram[1056] = 22;
    exp_54_ram[1057] = 195;
    exp_54_ram[1058] = 0;
    exp_54_ram[1059] = 1;
    exp_54_ram[1060] = 1;
    exp_54_ram[1061] = 0;
    exp_54_ram[1062] = 0;
    exp_54_ram[1063] = 249;
    exp_54_ram[1064] = 0;
    exp_54_ram[1065] = 0;
    exp_54_ram[1066] = 0;
    exp_54_ram[1067] = 0;
    exp_54_ram[1068] = 64;
    exp_54_ram[1069] = 0;
    exp_54_ram[1070] = 0;
    exp_54_ram[1071] = 0;
    exp_54_ram[1072] = 64;
    exp_54_ram[1073] = 0;
    exp_54_ram[1074] = 0;
    exp_54_ram[1075] = 0;
    exp_54_ram[1076] = 65;
    exp_54_ram[1077] = 65;
    exp_54_ram[1078] = 0;
    exp_54_ram[1079] = 0;
    exp_54_ram[1080] = 0;
    exp_54_ram[1081] = 0;
    exp_54_ram[1082] = 0;
    exp_54_ram[1083] = 65;
    exp_54_ram[1084] = 0;
    exp_54_ram[1085] = 0;
    exp_54_ram[1086] = 0;
    exp_54_ram[1087] = 24;
    exp_54_ram[1088] = 255;
    exp_54_ram[1089] = 0;
    exp_54_ram[1090] = 187;
    exp_54_ram[1091] = 0;
    exp_54_ram[1092] = 65;
    exp_54_ram[1093] = 0;
    exp_54_ram[1094] = 0;
    exp_54_ram[1095] = 1;
    exp_54_ram[1096] = 0;
    exp_54_ram[1097] = 1;
    exp_54_ram[1098] = 0;
    exp_54_ram[1099] = 1;
    exp_54_ram[1100] = 0;
    exp_54_ram[1101] = 1;
    exp_54_ram[1102] = 1;
    exp_54_ram[1103] = 1;
    exp_54_ram[1104] = 0;
    exp_54_ram[1105] = 0;
    exp_54_ram[1106] = 0;
    exp_54_ram[1107] = 0;
    exp_54_ram[1108] = 2;
    exp_54_ram[1109] = 0;
    exp_54_ram[1110] = 255;
    exp_54_ram[1111] = 0;
    exp_54_ram[1112] = 0;
    exp_54_ram[1113] = 0;
    exp_54_ram[1114] = 230;
    exp_54_ram[1115] = 0;
    exp_54_ram[1116] = 61;
    exp_54_ram[1117] = 0;
    exp_54_ram[1118] = 241;
    exp_54_ram[1119] = 0;
    exp_54_ram[1120] = 135;
    exp_54_ram[1121] = 0;
    exp_54_ram[1122] = 0;
    exp_54_ram[1123] = 0;
    exp_54_ram[1124] = 0;
    exp_54_ram[1125] = 0;
    exp_54_ram[1126] = 0;
    exp_54_ram[1127] = 0;
    exp_54_ram[1128] = 1;
    exp_54_ram[1129] = 0;
    exp_54_ram[1130] = 255;
    exp_54_ram[1131] = 0;
    exp_54_ram[1132] = 0;
    exp_54_ram[1133] = 0;
    exp_54_ram[1134] = 0;
    exp_54_ram[1135] = 0;
    exp_54_ram[1136] = 0;
    exp_54_ram[1137] = 249;
    exp_54_ram[1138] = 64;
    exp_54_ram[1139] = 0;
    exp_54_ram[1140] = 0;
    exp_54_ram[1141] = 64;
    exp_54_ram[1142] = 64;
    exp_54_ram[1143] = 135;
    exp_54_ram[1144] = 0;
    exp_54_ram[1145] = 0;
    exp_54_ram[1146] = 0;
    exp_54_ram[1147] = 0;
    exp_54_ram[1148] = 0;
    exp_54_ram[1149] = 1;
    exp_54_ram[1150] = 0;
    exp_54_ram[1151] = 249;
    exp_54_ram[1152] = 0;
    exp_54_ram[1153] = 6;
    exp_54_ram[1154] = 1;
    exp_54_ram[1155] = 0;
    exp_54_ram[1156] = 62;
    exp_54_ram[1157] = 1;
    exp_54_ram[1158] = 6;
    exp_54_ram[1159] = 6;
    exp_54_ram[1160] = 7;
    exp_54_ram[1161] = 5;
    exp_54_ram[1162] = 5;
    exp_54_ram[1163] = 195;
    exp_54_ram[1164] = 0;
    exp_54_ram[1165] = 2;
    exp_54_ram[1166] = 63;
    exp_54_ram[1167] = 2;
    exp_54_ram[1168] = 194;
    exp_54_ram[1169] = 1;
    exp_54_ram[1170] = 0;
    exp_54_ram[1171] = 131;
    exp_54_ram[1172] = 0;
    exp_54_ram[1173] = 0;
    exp_54_ram[1174] = 1;
    exp_54_ram[1175] = 2;
    exp_54_ram[1176] = 0;
    exp_54_ram[1177] = 0;
    exp_54_ram[1178] = 131;
    exp_54_ram[1179] = 191;
    exp_54_ram[1180] = 1;
    exp_54_ram[1181] = 1;
    exp_54_ram[1182] = 0;
    exp_54_ram[1183] = 0;
    exp_54_ram[1184] = 0;
    exp_54_ram[1185] = 0;
    exp_54_ram[1186] = 2;
    exp_54_ram[1187] = 0;
    exp_54_ram[1188] = 189;
    exp_54_ram[1189] = 1;
    exp_54_ram[1190] = 0;
    exp_54_ram[1191] = 0;
    exp_54_ram[1192] = 3;
    exp_54_ram[1193] = 15;
    exp_54_ram[1194] = 0;
    exp_54_ram[1195] = 0;
    exp_54_ram[1196] = 0;
    exp_54_ram[1197] = 1;
    exp_54_ram[1198] = 3;
    exp_54_ram[1199] = 0;
    exp_54_ram[1200] = 0;
    exp_54_ram[1201] = 0;
    exp_54_ram[1202] = 3;
    exp_54_ram[1203] = 0;
    exp_54_ram[1204] = 0;
    exp_54_ram[1205] = 12;
    exp_54_ram[1206] = 0;
    exp_54_ram[1207] = 0;
    exp_54_ram[1208] = 0;
    exp_54_ram[1209] = 1;
    exp_54_ram[1210] = 3;
    exp_54_ram[1211] = 0;
    exp_54_ram[1212] = 0;
    exp_54_ram[1213] = 0;
    exp_54_ram[1214] = 3;
    exp_54_ram[1215] = 0;
    exp_54_ram[1216] = 0;
    exp_54_ram[1217] = 9;
    exp_54_ram[1218] = 0;
    exp_54_ram[1219] = 0;
    exp_54_ram[1220] = 0;
    exp_54_ram[1221] = 1;
    exp_54_ram[1222] = 3;
    exp_54_ram[1223] = 0;
    exp_54_ram[1224] = 0;
    exp_54_ram[1225] = 0;
    exp_54_ram[1226] = 3;
    exp_54_ram[1227] = 0;
    exp_54_ram[1228] = 0;
    exp_54_ram[1229] = 6;
    exp_54_ram[1230] = 0;
    exp_54_ram[1231] = 0;
    exp_54_ram[1232] = 0;
    exp_54_ram[1233] = 1;
    exp_54_ram[1234] = 3;
    exp_54_ram[1235] = 0;
    exp_54_ram[1236] = 0;
    exp_54_ram[1237] = 62;
    exp_54_ram[1238] = 3;
    exp_54_ram[1239] = 0;
    exp_54_ram[1240] = 1;
    exp_54_ram[1241] = 118;
    exp_54_ram[1242] = 2;
    exp_54_ram[1243] = 0;
    exp_54_ram[1244] = 0;
    exp_54_ram[1245] = 0;
    exp_54_ram[1246] = 0;
    exp_54_ram[1247] = 6;
    exp_54_ram[1248] = 3;
    exp_54_ram[1249] = 0;
    exp_54_ram[1250] = 0;
    exp_54_ram[1251] = 0;
    exp_54_ram[1252] = 0;
    exp_54_ram[1253] = 0;
    exp_54_ram[1254] = 0;
    exp_54_ram[1255] = 0;
    exp_54_ram[1256] = 3;
    exp_54_ram[1257] = 0;
    exp_54_ram[1258] = 126;
    exp_54_ram[1259] = 0;
    exp_54_ram[1260] = 0;
    exp_54_ram[1261] = 0;
    exp_54_ram[1262] = 6;
    exp_54_ram[1263] = 3;
    exp_54_ram[1264] = 0;
    exp_54_ram[1265] = 0;
    exp_54_ram[1266] = 6;
    exp_54_ram[1267] = 6;
    exp_54_ram[1268] = 3;
    exp_54_ram[1269] = 0;
    exp_54_ram[1270] = 0;
    exp_54_ram[1271] = 0;
    exp_54_ram[1272] = 6;
    exp_54_ram[1273] = 5;
    exp_54_ram[1274] = 131;
    exp_54_ram[1275] = 5;
    exp_54_ram[1276] = 7;
    exp_54_ram[1277] = 0;
    exp_54_ram[1278] = 252;
    exp_54_ram[1279] = 3;
    exp_54_ram[1280] = 0;
    exp_54_ram[1281] = 2;
    exp_54_ram[1282] = 2;
    exp_54_ram[1283] = 3;
    exp_54_ram[1284] = 3;
    exp_54_ram[1285] = 3;
    exp_54_ram[1286] = 2;
    exp_54_ram[1287] = 3;
    exp_54_ram[1288] = 1;
    exp_54_ram[1289] = 1;
    exp_54_ram[1290] = 1;
    exp_54_ram[1291] = 0;
    exp_54_ram[1292] = 0;
    exp_54_ram[1293] = 0;
    exp_54_ram[1294] = 123;
    exp_54_ram[1295] = 0;
    exp_54_ram[1296] = 24;
    exp_54_ram[1297] = 0;
    exp_54_ram[1298] = 173;
    exp_54_ram[1299] = 0;
    exp_54_ram[1300] = 0;
    exp_54_ram[1301] = 22;
    exp_54_ram[1302] = 134;
    exp_54_ram[1303] = 0;
    exp_54_ram[1304] = 0;
    exp_54_ram[1305] = 2;
    exp_54_ram[1306] = 0;
    exp_54_ram[1307] = 64;
    exp_54_ram[1308] = 0;
    exp_54_ram[1309] = 64;
    exp_54_ram[1310] = 0;
    exp_54_ram[1311] = 0;
    exp_54_ram[1312] = 252;
    exp_54_ram[1313] = 0;
    exp_54_ram[1314] = 0;
    exp_54_ram[1315] = 0;
    exp_54_ram[1316] = 24;
    exp_54_ram[1317] = 0;
    exp_54_ram[1318] = 0;
    exp_54_ram[1319] = 173;
    exp_54_ram[1320] = 0;
    exp_54_ram[1321] = 0;
    exp_54_ram[1322] = 0;
    exp_54_ram[1323] = 0;
    exp_54_ram[1324] = 128;
    exp_54_ram[1325] = 0;
    exp_54_ram[1326] = 2;
    exp_54_ram[1327] = 64;
    exp_54_ram[1328] = 0;
    exp_54_ram[1329] = 1;
    exp_54_ram[1330] = 1;
    exp_54_ram[1331] = 0;
    exp_54_ram[1332] = 64;
    exp_54_ram[1333] = 252;
    exp_54_ram[1334] = 0;
    exp_54_ram[1335] = 0;
    exp_54_ram[1336] = 24;
    exp_54_ram[1337] = 107;
    exp_54_ram[1338] = 0;
    exp_54_ram[1339] = 0;
    exp_54_ram[1340] = 0;
    exp_54_ram[1341] = 0;
    exp_54_ram[1342] = 0;
    exp_54_ram[1343] = 0;
    exp_54_ram[1344] = 225;
    exp_54_ram[1345] = 105;
    exp_54_ram[1346] = 0;
    exp_54_ram[1347] = 0;
    exp_54_ram[1348] = 0;
    exp_54_ram[1349] = 0;
    exp_54_ram[1350] = 3;
    exp_54_ram[1351] = 137;
    exp_54_ram[1352] = 103;
    exp_54_ram[1353] = 0;
    exp_54_ram[1354] = 0;
    exp_54_ram[1355] = 0;
    exp_54_ram[1356] = 0;
    exp_54_ram[1357] = 0;
    exp_54_ram[1358] = 1;
    exp_54_ram[1359] = 1;
    exp_54_ram[1360] = 1;
    exp_54_ram[1361] = 0;
    exp_54_ram[1362] = 0;
    exp_54_ram[1363] = 0;
    exp_54_ram[1364] = 129;
    exp_54_ram[1365] = 0;
    exp_54_ram[1366] = 1;
    exp_54_ram[1367] = 3;
    exp_54_ram[1368] = 0;
    exp_54_ram[1369] = 3;
    exp_54_ram[1370] = 3;
    exp_54_ram[1371] = 3;
    exp_54_ram[1372] = 2;
    exp_54_ram[1373] = 2;
    exp_54_ram[1374] = 2;
    exp_54_ram[1375] = 2;
    exp_54_ram[1376] = 1;
    exp_54_ram[1377] = 1;
    exp_54_ram[1378] = 1;
    exp_54_ram[1379] = 4;
    exp_54_ram[1380] = 0;
    exp_54_ram[1381] = 246;
    exp_54_ram[1382] = 9;
    exp_54_ram[1383] = 1;
    exp_54_ram[1384] = 2;
    exp_54_ram[1385] = 8;
    exp_54_ram[1386] = 9;
    exp_54_ram[1387] = 1;
    exp_54_ram[1388] = 9;
    exp_54_ram[1389] = 9;
    exp_54_ram[1390] = 0;
    exp_54_ram[1391] = 0;
    exp_54_ram[1392] = 0;
    exp_54_ram[1393] = 3;
    exp_54_ram[1394] = 0;
    exp_54_ram[1395] = 8;
    exp_54_ram[1396] = 8;
    exp_54_ram[1397] = 9;
    exp_54_ram[1398] = 5;
    exp_54_ram[1399] = 4;
    exp_54_ram[1400] = 5;
    exp_54_ram[1401] = 5;
    exp_54_ram[1402] = 2;
    exp_54_ram[1403] = 2;
    exp_54_ram[1404] = 4;
    exp_54_ram[1405] = 134;
    exp_54_ram[1406] = 0;
    exp_54_ram[1407] = 158;
    exp_54_ram[1408] = 0;
    exp_54_ram[1409] = 0;
    exp_54_ram[1410] = 3;
    exp_54_ram[1411] = 222;
    exp_54_ram[1412] = 5;
    exp_54_ram[1413] = 4;
    exp_54_ram[1414] = 2;
    exp_54_ram[1415] = 3;
    exp_54_ram[1416] = 64;
    exp_54_ram[1417] = 0;
    exp_54_ram[1418] = 4;
    exp_54_ram[1419] = 131;
    exp_54_ram[1420] = 0;
    exp_54_ram[1421] = 155;
    exp_54_ram[1422] = 2;
    exp_54_ram[1423] = 0;
    exp_54_ram[1424] = 0;
    exp_54_ram[1425] = 0;
    exp_54_ram[1426] = 5;
    exp_54_ram[1427] = 7;
    exp_54_ram[1428] = 6;
    exp_54_ram[1429] = 7;
    exp_54_ram[1430] = 7;
    exp_54_ram[1431] = 6;
    exp_54_ram[1432] = 4;
    exp_54_ram[1433] = 255;
    exp_54_ram[1434] = 0;
    exp_54_ram[1435] = 151;
    exp_54_ram[1436] = 0;
    exp_54_ram[1437] = 0;
    exp_54_ram[1438] = 3;
    exp_54_ram[1439] = 215;
    exp_54_ram[1440] = 2;
    exp_54_ram[1441] = 5;
    exp_54_ram[1442] = 0;
    exp_54_ram[1443] = 6;
    exp_54_ram[1444] = 253;
    exp_54_ram[1445] = 0;
    exp_54_ram[1446] = 149;
    exp_54_ram[1447] = 2;
    exp_54_ram[1448] = 0;
    exp_54_ram[1449] = 0;
    exp_54_ram[1450] = 0;
    exp_54_ram[1451] = 0;
    exp_54_ram[1452] = 251;
    exp_54_ram[1453] = 0;
    exp_54_ram[1454] = 147;
    exp_54_ram[1455] = 0;
    exp_54_ram[1456] = 0;
    exp_54_ram[1457] = 0;
    exp_54_ram[1458] = 0;
    exp_54_ram[1459] = 0;
    exp_54_ram[1460] = 0;
    exp_54_ram[1461] = 0;
    exp_54_ram[1462] = 0;
    exp_54_ram[1463] = 1;
    exp_54_ram[1464] = 0;
    exp_54_ram[1465] = 9;
    exp_54_ram[1466] = 9;
    exp_54_ram[1467] = 9;
    exp_54_ram[1468] = 9;
    exp_54_ram[1469] = 8;
    exp_54_ram[1470] = 8;
    exp_54_ram[1471] = 8;
    exp_54_ram[1472] = 8;
    exp_54_ram[1473] = 10;
    exp_54_ram[1474] = 0;
    exp_54_ram[1475] = 248;
    exp_54_ram[1476] = 0;
    exp_54_ram[1477] = 7;
    exp_54_ram[1478] = 2;
    exp_54_ram[1479] = 0;
    exp_54_ram[1480] = 3;
    exp_54_ram[1481] = 6;
    exp_54_ram[1482] = 6;
    exp_54_ram[1483] = 6;
    exp_54_ram[1484] = 7;
    exp_54_ram[1485] = 242;
    exp_54_ram[1486] = 2;
    exp_54_ram[1487] = 3;
    exp_54_ram[1488] = 0;
    exp_54_ram[1489] = 2;
    exp_54_ram[1490] = 241;
    exp_54_ram[1491] = 0;
    exp_54_ram[1492] = 137;
    exp_54_ram[1493] = 0;
    exp_54_ram[1494] = 0;
    exp_54_ram[1495] = 7;
    exp_54_ram[1496] = 0;
    exp_54_ram[1497] = 225;
    exp_54_ram[1498] = 0;
    exp_54_ram[1499] = 0;
    exp_54_ram[1500] = 0;
    exp_54_ram[1501] = 0;
    exp_54_ram[1502] = 0;
    exp_54_ram[1503] = 0;
    exp_54_ram[1504] = 0;
    exp_54_ram[1505] = 199;
    exp_54_ram[1506] = 2;
    exp_54_ram[1507] = 0;
    exp_54_ram[1508] = 0;
    exp_54_ram[1509] = 236;
    exp_54_ram[1510] = 7;
    exp_54_ram[1511] = 0;
    exp_54_ram[1512] = 2;
    exp_54_ram[1513] = 7;
    exp_54_ram[1514] = 0;
    exp_54_ram[1515] = 7;
    exp_54_ram[1516] = 7;
    exp_54_ram[1517] = 6;
    exp_54_ram[1518] = 0;
    exp_54_ram[1519] = 7;
    exp_54_ram[1520] = 8;
    exp_54_ram[1521] = 0;
    exp_54_ram[1522] = 250;
    exp_54_ram[1523] = 3;
    exp_54_ram[1524] = 2;
    exp_54_ram[1525] = 0;
    exp_54_ram[1526] = 232;
    exp_54_ram[1527] = 0;
    exp_54_ram[1528] = 219;
    exp_54_ram[1529] = 65;
    exp_54_ram[1530] = 0;
    exp_54_ram[1531] = 0;
    exp_54_ram[1532] = 0;
    exp_54_ram[1533] = 0;
    exp_54_ram[1534] = 0;
    exp_54_ram[1535] = 0;
    exp_54_ram[1536] = 246;
    exp_54_ram[1537] = 0;
    exp_54_ram[1538] = 225;
    exp_54_ram[1539] = 0;
    exp_54_ram[1540] = 246;
    exp_54_ram[1541] = 2;
    exp_54_ram[1542] = 2;
    exp_54_ram[1543] = 3;
    exp_54_ram[1544] = 0;
    exp_54_ram[1545] = 227;
    exp_54_ram[1546] = 0;
    exp_54_ram[1547] = 214;
    exp_54_ram[1548] = 0;
    exp_54_ram[1549] = 0;
    exp_54_ram[1550] = 225;
    exp_54_ram[1551] = 2;
    exp_54_ram[1552] = 246;
    exp_54_ram[1553] = 2;
    exp_54_ram[1554] = 245;
    exp_54_ram[1555] = 249;
    exp_54_ram[1556] = 0;
    exp_54_ram[1557] = 0;
    exp_54_ram[1558] = 3;
    exp_54_ram[1559] = 6;
    exp_54_ram[1560] = 185;
    exp_54_ram[1561] = 3;
    exp_54_ram[1562] = 2;
    exp_54_ram[1563] = 0;
    exp_54_ram[1564] = 223;
    exp_54_ram[1565] = 0;
    exp_54_ram[1566] = 209;
    exp_54_ram[1567] = 6;
    exp_54_ram[1568] = 7;
    exp_54_ram[1569] = 0;
    exp_54_ram[1570] = 251;
    exp_54_ram[1571] = 4;
    exp_54_ram[1572] = 5;
    exp_54_ram[1573] = 0;
    exp_54_ram[1574] = 0;
    exp_54_ram[1575] = 4;
    exp_54_ram[1576] = 0;
    exp_54_ram[1577] = 0;
    exp_54_ram[1578] = 4;
    exp_54_ram[1579] = 3;
    exp_54_ram[1580] = 249;
    exp_54_ram[1581] = 0;
    exp_54_ram[1582] = 0;
    exp_54_ram[1583] = 0;
    exp_54_ram[1584] = 225;
    exp_54_ram[1585] = 1;
    exp_54_ram[1586] = 0;
    exp_54_ram[1587] = 0;
    exp_54_ram[1588] = 0;
    exp_54_ram[1589] = 178;
    exp_54_ram[1590] = 0;
    exp_54_ram[1591] = 0;
    exp_54_ram[1592] = 2;
    exp_54_ram[1593] = 133;
    exp_54_ram[1594] = 215;
    exp_54_ram[1595] = 0;
    exp_54_ram[1596] = 0;
    exp_54_ram[1597] = 245;
    exp_54_ram[1598] = 133;
    exp_54_ram[1599] = 2;
    exp_54_ram[1600] = 4;
    exp_54_ram[1601] = 133;
    exp_54_ram[1602] = 4;
    exp_54_ram[1603] = 4;
    exp_54_ram[1604] = 4;
    exp_54_ram[1605] = 3;
    exp_54_ram[1606] = 5;
    exp_54_ram[1607] = 0;
    exp_54_ram[1608] = 253;
    exp_54_ram[1609] = 2;
    exp_54_ram[1610] = 2;
    exp_54_ram[1611] = 3;
    exp_54_ram[1612] = 3;
    exp_54_ram[1613] = 3;
    exp_54_ram[1614] = 252;
    exp_54_ram[1615] = 232;
    exp_54_ram[1616] = 254;
    exp_54_ram[1617] = 254;
    exp_54_ram[1618] = 0;
    exp_54_ram[1619] = 231;
    exp_54_ram[1620] = 0;
    exp_54_ram[1621] = 0;
    exp_54_ram[1622] = 254;
    exp_54_ram[1623] = 254;
    exp_54_ram[1624] = 64;
    exp_54_ram[1625] = 0;
    exp_54_ram[1626] = 1;
    exp_54_ram[1627] = 64;
    exp_54_ram[1628] = 65;
    exp_54_ram[1629] = 0;
    exp_54_ram[1630] = 253;
    exp_54_ram[1631] = 0;
    exp_54_ram[1632] = 0;
    exp_54_ram[1633] = 0;
    exp_54_ram[1634] = 0;
    exp_54_ram[1635] = 252;
    exp_54_ram[1636] = 0;
    exp_54_ram[1637] = 0;
    exp_54_ram[1638] = 0;
    exp_54_ram[1639] = 0;
    exp_54_ram[1640] = 0;
    exp_54_ram[1641] = 250;
    exp_54_ram[1642] = 0;
    exp_54_ram[1643] = 0;
    exp_54_ram[1644] = 2;
    exp_54_ram[1645] = 2;
    exp_54_ram[1646] = 2;
    exp_54_ram[1647] = 2;
    exp_54_ram[1648] = 3;
    exp_54_ram[1649] = 0;
    exp_54_ram[1650] = 255;
    exp_54_ram[1651] = 0;
    exp_54_ram[1652] = 0;
    exp_54_ram[1653] = 1;
    exp_54_ram[1654] = 89;
    exp_54_ram[1655] = 231;
    exp_54_ram[1656] = 0;
    exp_54_ram[1657] = 0;
    exp_54_ram[1658] = 0;
    exp_54_ram[1659] = 1;
    exp_54_ram[1660] = 0;
    exp_54_ram[1661] = 254;
    exp_54_ram[1662] = 0;
    exp_54_ram[1663] = 0;
    exp_54_ram[1664] = 2;
    exp_54_ram[1665] = 90;
    exp_54_ram[1666] = 228;
    exp_54_ram[1667] = 0;
    exp_54_ram[1668] = 254;
    exp_54_ram[1669] = 254;
    exp_54_ram[1670] = 10;
    exp_54_ram[1671] = 254;
    exp_54_ram[1672] = 92;
    exp_54_ram[1673] = 170;
    exp_54_ram[1674] = 3;
    exp_54_ram[1675] = 254;
    exp_54_ram[1676] = 0;
    exp_54_ram[1677] = 254;
    exp_54_ram[1678] = 0;
    exp_54_ram[1679] = 61;
    exp_54_ram[1680] = 0;
    exp_54_ram[1681] = 254;
    exp_54_ram[1682] = 220;
    exp_54_ram[1683] = 0;
    exp_54_ram[1684] = 61;
    exp_54_ram[1685] = 0;
    exp_54_ram[1686] = 2;
    exp_54_ram[1687] = 0;
    exp_54_ram[1688] = 236;
    exp_54_ram[1689] = 254;
    exp_54_ram[1690] = 7;
    exp_54_ram[1691] = 252;
    exp_54_ram[1692] = 3;
    exp_54_ram[1693] = 254;
    exp_54_ram[1694] = 64;
    exp_54_ram[1695] = 254;
    exp_54_ram[1696] = 0;
    exp_54_ram[1697] = 61;
    exp_54_ram[1698] = 0;
    exp_54_ram[1699] = 254;
    exp_54_ram[1700] = 216;
    exp_54_ram[1701] = 0;
    exp_54_ram[1702] = 61;
    exp_54_ram[1703] = 0;
    exp_54_ram[1704] = 2;
    exp_54_ram[1705] = 0;
    exp_54_ram[1706] = 231;
    exp_54_ram[1707] = 254;
    exp_54_ram[1708] = 0;
    exp_54_ram[1709] = 252;
    exp_54_ram[1710] = 254;
    exp_54_ram[1711] = 0;
    exp_54_ram[1712] = 254;
    exp_54_ram[1713] = 254;
    exp_54_ram[1714] = 0;
    exp_54_ram[1715] = 244;
    exp_54_ram[1716] = 0;
    exp_54_ram[1717] = 61;
    exp_54_ram[1718] = 0;
    exp_54_ram[1719] = 0;
    exp_54_ram[1720] = 211;
    exp_54_ram[1721] = 0;
    exp_54_ram[1722] = 1;
    exp_54_ram[1723] = 1;
    exp_54_ram[1724] = 2;
    exp_54_ram[1725] = 0;
    exp_54_ram[1726] = 254;
    exp_54_ram[1727] = 0;
    exp_54_ram[1728] = 0;
    exp_54_ram[1729] = 2;
    exp_54_ram[1730] = 254;
    exp_54_ram[1731] = 5;
    exp_54_ram[1732] = 0;
    exp_54_ram[1733] = 254;
    exp_54_ram[1734] = 0;
    exp_54_ram[1735] = 0;
    exp_54_ram[1736] = 254;
    exp_54_ram[1737] = 1;
    exp_54_ram[1738] = 0;
    exp_54_ram[1739] = 254;
    exp_54_ram[1740] = 0;
    exp_54_ram[1741] = 0;
    exp_54_ram[1742] = 254;
    exp_54_ram[1743] = 1;
    exp_54_ram[1744] = 0;
    exp_54_ram[1745] = 254;
    exp_54_ram[1746] = 0;
    exp_54_ram[1747] = 254;
    exp_54_ram[1748] = 255;
    exp_54_ram[1749] = 2;
    exp_54_ram[1750] = 254;
    exp_54_ram[1751] = 187;
    exp_54_ram[1752] = 0;
    exp_54_ram[1753] = 0;
    exp_54_ram[1754] = 0;
    exp_54_ram[1755] = 0;
    exp_54_ram[1756] = 227;
    exp_54_ram[1757] = 0;
    exp_54_ram[1758] = 222;
    exp_54_ram[1759] = 0;
    exp_54_ram[1760] = 0;
    exp_54_ram[1761] = 254;
    exp_54_ram[1762] = 254;
    exp_54_ram[1763] = 254;
    exp_54_ram[1764] = 0;
    exp_54_ram[1765] = 207;
    exp_54_ram[1766] = 254;
    exp_54_ram[1767] = 254;
    exp_54_ram[1768] = 229;
    exp_54_ram[1769] = 0;
    exp_54_ram[1770] = 0;
    exp_54_ram[1771] = 202;
    exp_54_ram[1772] = 0;
    exp_54_ram[1773] = 61;
    exp_54_ram[1774] = 0;
    exp_54_ram[1775] = 214;
    exp_54_ram[1776] = 251;
    exp_54_ram[1777] = 249;
    exp_54_ram[1778] = 6;
    exp_54_ram[1779] = 6;
    exp_54_ram[1780] = 7;
    exp_54_ram[1781] = 7;
    exp_54_ram[1782] = 5;
    exp_54_ram[1783] = 5;
    exp_54_ram[1784] = 5;
    exp_54_ram[1785] = 5;
    exp_54_ram[1786] = 5;
    exp_54_ram[1787] = 5;
    exp_54_ram[1788] = 5;
    exp_54_ram[1789] = 5;
    exp_54_ram[1790] = 7;
    exp_54_ram[1791] = 0;
    exp_54_ram[1792] = 250;
    exp_54_ram[1793] = 0;
    exp_54_ram[1794] = 0;
    exp_54_ram[1795] = 250;
    exp_54_ram[1796] = 250;
    exp_54_ram[1797] = 187;
    exp_54_ram[1798] = 252;
    exp_54_ram[1799] = 252;
    exp_54_ram[1800] = 252;
    exp_54_ram[1801] = 6;
    exp_54_ram[1802] = 251;
    exp_54_ram[1803] = 18;
    exp_54_ram[1804] = 103;
    exp_54_ram[1805] = 2;
    exp_54_ram[1806] = 250;
    exp_54_ram[1807] = 251;
    exp_54_ram[1808] = 18;
    exp_54_ram[1809] = 103;
    exp_54_ram[1810] = 2;
    exp_54_ram[1811] = 250;
    exp_54_ram[1812] = 251;
    exp_54_ram[1813] = 18;
    exp_54_ram[1814] = 103;
    exp_54_ram[1815] = 2;
    exp_54_ram[1816] = 250;
    exp_54_ram[1817] = 251;
    exp_54_ram[1818] = 18;
    exp_54_ram[1819] = 103;
    exp_54_ram[1820] = 2;
    exp_54_ram[1821] = 250;
    exp_54_ram[1822] = 252;
    exp_54_ram[1823] = 0;
    exp_54_ram[1824] = 252;
    exp_54_ram[1825] = 180;
    exp_54_ram[1826] = 0;
    exp_54_ram[1827] = 0;
    exp_54_ram[1828] = 252;
    exp_54_ram[1829] = 252;
    exp_54_ram[1830] = 64;
    exp_54_ram[1831] = 0;
    exp_54_ram[1832] = 1;
    exp_54_ram[1833] = 64;
    exp_54_ram[1834] = 65;
    exp_54_ram[1835] = 0;
    exp_54_ram[1836] = 0;
    exp_54_ram[1837] = 61;
    exp_54_ram[1838] = 250;
    exp_54_ram[1839] = 250;
    exp_54_ram[1840] = 250;
    exp_54_ram[1841] = 250;
    exp_54_ram[1842] = 0;
    exp_54_ram[1843] = 0;
    exp_54_ram[1844] = 244;
    exp_54_ram[1845] = 0;
    exp_54_ram[1846] = 0;
    exp_54_ram[1847] = 0;
    exp_54_ram[1848] = 0;
    exp_54_ram[1849] = 0;
    exp_54_ram[1850] = 244;
    exp_54_ram[1851] = 252;
    exp_54_ram[1852] = 92;
    exp_54_ram[1853] = 253;
    exp_54_ram[1854] = 173;
    exp_54_ram[1855] = 252;
    exp_54_ram[1856] = 252;
    exp_54_ram[1857] = 252;
    exp_54_ram[1858] = 18;
    exp_54_ram[1859] = 251;
    exp_54_ram[1860] = 251;
    exp_54_ram[1861] = 18;
    exp_54_ram[1862] = 103;
    exp_54_ram[1863] = 2;
    exp_54_ram[1864] = 0;
    exp_54_ram[1865] = 2;
    exp_54_ram[1866] = 0;
    exp_54_ram[1867] = 18;
    exp_54_ram[1868] = 103;
    exp_54_ram[1869] = 2;
    exp_54_ram[1870] = 2;
    exp_54_ram[1871] = 0;
    exp_54_ram[1872] = 1;
    exp_54_ram[1873] = 0;
    exp_54_ram[1874] = 251;
    exp_54_ram[1875] = 251;
    exp_54_ram[1876] = 251;
    exp_54_ram[1877] = 251;
    exp_54_ram[1878] = 18;
    exp_54_ram[1879] = 103;
    exp_54_ram[1880] = 2;
    exp_54_ram[1881] = 0;
    exp_54_ram[1882] = 2;
    exp_54_ram[1883] = 0;
    exp_54_ram[1884] = 18;
    exp_54_ram[1885] = 103;
    exp_54_ram[1886] = 2;
    exp_54_ram[1887] = 2;
    exp_54_ram[1888] = 0;
    exp_54_ram[1889] = 1;
    exp_54_ram[1890] = 0;
    exp_54_ram[1891] = 251;
    exp_54_ram[1892] = 251;
    exp_54_ram[1893] = 251;
    exp_54_ram[1894] = 251;
    exp_54_ram[1895] = 18;
    exp_54_ram[1896] = 103;
    exp_54_ram[1897] = 2;
    exp_54_ram[1898] = 0;
    exp_54_ram[1899] = 2;
    exp_54_ram[1900] = 0;
    exp_54_ram[1901] = 18;
    exp_54_ram[1902] = 103;
    exp_54_ram[1903] = 2;
    exp_54_ram[1904] = 2;
    exp_54_ram[1905] = 0;
    exp_54_ram[1906] = 1;
    exp_54_ram[1907] = 0;
    exp_54_ram[1908] = 251;
    exp_54_ram[1909] = 251;
    exp_54_ram[1910] = 251;
    exp_54_ram[1911] = 251;
    exp_54_ram[1912] = 18;
    exp_54_ram[1913] = 103;
    exp_54_ram[1914] = 2;
    exp_54_ram[1915] = 0;
    exp_54_ram[1916] = 2;
    exp_54_ram[1917] = 0;
    exp_54_ram[1918] = 18;
    exp_54_ram[1919] = 103;
    exp_54_ram[1920] = 2;
    exp_54_ram[1921] = 2;
    exp_54_ram[1922] = 0;
    exp_54_ram[1923] = 1;
    exp_54_ram[1924] = 0;
    exp_54_ram[1925] = 251;
    exp_54_ram[1926] = 251;
    exp_54_ram[1927] = 252;
    exp_54_ram[1928] = 0;
    exp_54_ram[1929] = 252;
    exp_54_ram[1930] = 154;
    exp_54_ram[1931] = 0;
    exp_54_ram[1932] = 0;
    exp_54_ram[1933] = 252;
    exp_54_ram[1934] = 252;
    exp_54_ram[1935] = 64;
    exp_54_ram[1936] = 0;
    exp_54_ram[1937] = 1;
    exp_54_ram[1938] = 64;
    exp_54_ram[1939] = 65;
    exp_54_ram[1940] = 0;
    exp_54_ram[1941] = 0;
    exp_54_ram[1942] = 61;
    exp_54_ram[1943] = 250;
    exp_54_ram[1944] = 250;
    exp_54_ram[1945] = 250;
    exp_54_ram[1946] = 250;
    exp_54_ram[1947] = 0;
    exp_54_ram[1948] = 0;
    exp_54_ram[1949] = 232;
    exp_54_ram[1950] = 0;
    exp_54_ram[1951] = 0;
    exp_54_ram[1952] = 0;
    exp_54_ram[1953] = 0;
    exp_54_ram[1954] = 0;
    exp_54_ram[1955] = 232;
    exp_54_ram[1956] = 252;
    exp_54_ram[1957] = 95;
    exp_54_ram[1958] = 226;
    exp_54_ram[1959] = 146;
    exp_54_ram[1960] = 252;
    exp_54_ram[1961] = 252;
    exp_54_ram[1962] = 252;
    exp_54_ram[1963] = 6;
    exp_54_ram[1964] = 251;
    exp_54_ram[1965] = 18;
    exp_54_ram[1966] = 103;
    exp_54_ram[1967] = 2;
    exp_54_ram[1968] = 250;
    exp_54_ram[1969] = 251;
    exp_54_ram[1970] = 18;
    exp_54_ram[1971] = 103;
    exp_54_ram[1972] = 2;
    exp_54_ram[1973] = 250;
    exp_54_ram[1974] = 251;
    exp_54_ram[1975] = 18;
    exp_54_ram[1976] = 103;
    exp_54_ram[1977] = 2;
    exp_54_ram[1978] = 250;
    exp_54_ram[1979] = 251;
    exp_54_ram[1980] = 18;
    exp_54_ram[1981] = 103;
    exp_54_ram[1982] = 2;
    exp_54_ram[1983] = 250;
    exp_54_ram[1984] = 252;
    exp_54_ram[1985] = 0;
    exp_54_ram[1986] = 252;
    exp_54_ram[1987] = 139;
    exp_54_ram[1988] = 0;
    exp_54_ram[1989] = 0;
    exp_54_ram[1990] = 252;
    exp_54_ram[1991] = 252;
    exp_54_ram[1992] = 64;
    exp_54_ram[1993] = 0;
    exp_54_ram[1994] = 1;
    exp_54_ram[1995] = 64;
    exp_54_ram[1996] = 65;
    exp_54_ram[1997] = 0;
    exp_54_ram[1998] = 0;
    exp_54_ram[1999] = 61;
    exp_54_ram[2000] = 248;
    exp_54_ram[2001] = 248;
    exp_54_ram[2002] = 249;
    exp_54_ram[2003] = 249;
    exp_54_ram[2004] = 0;
    exp_54_ram[2005] = 0;
    exp_54_ram[2006] = 244;
    exp_54_ram[2007] = 0;
    exp_54_ram[2008] = 0;
    exp_54_ram[2009] = 0;
    exp_54_ram[2010] = 0;
    exp_54_ram[2011] = 0;
    exp_54_ram[2012] = 244;
    exp_54_ram[2013] = 252;
    exp_54_ram[2014] = 97;
    exp_54_ram[2015] = 212;
    exp_54_ram[2016] = 132;
    exp_54_ram[2017] = 252;
    exp_54_ram[2018] = 252;
    exp_54_ram[2019] = 252;
    exp_54_ram[2020] = 13;
    exp_54_ram[2021] = 251;
    exp_54_ram[2022] = 251;
    exp_54_ram[2023] = 18;
    exp_54_ram[2024] = 103;
    exp_54_ram[2025] = 0;
    exp_54_ram[2026] = 0;
    exp_54_ram[2027] = 0;
    exp_54_ram[2028] = 141;
    exp_54_ram[2029] = 0;
    exp_54_ram[2030] = 0;
    exp_54_ram[2031] = 250;
    exp_54_ram[2032] = 250;
    exp_54_ram[2033] = 251;
    exp_54_ram[2034] = 251;
    exp_54_ram[2035] = 18;
    exp_54_ram[2036] = 103;
    exp_54_ram[2037] = 0;
    exp_54_ram[2038] = 0;
    exp_54_ram[2039] = 0;
    exp_54_ram[2040] = 138;
    exp_54_ram[2041] = 0;
    exp_54_ram[2042] = 0;
    exp_54_ram[2043] = 250;
    exp_54_ram[2044] = 250;
    exp_54_ram[2045] = 251;
    exp_54_ram[2046] = 251;
    exp_54_ram[2047] = 18;
    exp_54_ram[2048] = 103;
    exp_54_ram[2049] = 0;
    exp_54_ram[2050] = 0;
    exp_54_ram[2051] = 0;
    exp_54_ram[2052] = 135;
    exp_54_ram[2053] = 0;
    exp_54_ram[2054] = 0;
    exp_54_ram[2055] = 250;
    exp_54_ram[2056] = 250;
    exp_54_ram[2057] = 251;
    exp_54_ram[2058] = 251;
    exp_54_ram[2059] = 18;
    exp_54_ram[2060] = 103;
    exp_54_ram[2061] = 0;
    exp_54_ram[2062] = 0;
    exp_54_ram[2063] = 0;
    exp_54_ram[2064] = 132;
    exp_54_ram[2065] = 0;
    exp_54_ram[2066] = 0;
    exp_54_ram[2067] = 250;
    exp_54_ram[2068] = 250;
    exp_54_ram[2069] = 252;
    exp_54_ram[2070] = 0;
    exp_54_ram[2071] = 252;
    exp_54_ram[2072] = 246;
    exp_54_ram[2073] = 0;
    exp_54_ram[2074] = 0;
    exp_54_ram[2075] = 252;
    exp_54_ram[2076] = 252;
    exp_54_ram[2077] = 64;
    exp_54_ram[2078] = 0;
    exp_54_ram[2079] = 1;
    exp_54_ram[2080] = 64;
    exp_54_ram[2081] = 65;
    exp_54_ram[2082] = 0;
    exp_54_ram[2083] = 0;
    exp_54_ram[2084] = 61;
    exp_54_ram[2085] = 0;
    exp_54_ram[2086] = 0;
    exp_54_ram[2087] = 0;
    exp_54_ram[2088] = 0;
    exp_54_ram[2089] = 238;
    exp_54_ram[2090] = 0;
    exp_54_ram[2091] = 0;
    exp_54_ram[2092] = 0;
    exp_54_ram[2093] = 0;
    exp_54_ram[2094] = 0;
    exp_54_ram[2095] = 236;
    exp_54_ram[2096] = 252;
    exp_54_ram[2097] = 100;
    exp_54_ram[2098] = 191;
    exp_54_ram[2099] = 0;
    exp_54_ram[2100] = 6;
    exp_54_ram[2101] = 6;
    exp_54_ram[2102] = 6;
    exp_54_ram[2103] = 6;
    exp_54_ram[2104] = 5;
    exp_54_ram[2105] = 5;
    exp_54_ram[2106] = 5;
    exp_54_ram[2107] = 5;
    exp_54_ram[2108] = 4;
    exp_54_ram[2109] = 4;
    exp_54_ram[2110] = 4;
    exp_54_ram[2111] = 4;
    exp_54_ram[2112] = 7;
    exp_54_ram[2113] = 0;
    exp_54_ram[2114] = 240;
    exp_54_ram[2115] = 14;
    exp_54_ram[2116] = 14;
    exp_54_ram[2117] = 16;
    exp_54_ram[2118] = 254;
    exp_54_ram[2119] = 2;
    exp_54_ram[2120] = 254;
    exp_54_ram[2121] = 15;
    exp_54_ram[2122] = 254;
    exp_54_ram[2123] = 255;
    exp_54_ram[2124] = 0;
    exp_54_ram[2125] = 248;
    exp_54_ram[2126] = 254;
    exp_54_ram[2127] = 0;
    exp_54_ram[2128] = 254;
    exp_54_ram[2129] = 254;
    exp_54_ram[2130] = 6;
    exp_54_ram[2131] = 252;
    exp_54_ram[2132] = 254;
    exp_54_ram[2133] = 11;
    exp_54_ram[2134] = 254;
    exp_54_ram[2135] = 102;
    exp_54_ram[2136] = 182;
    exp_54_ram[2137] = 254;
    exp_54_ram[2138] = 240;
    exp_54_ram[2139] = 0;
    exp_54_ram[2140] = 6;
    exp_54_ram[2141] = 254;
    exp_54_ram[2142] = 64;
    exp_54_ram[2143] = 0;
    exp_54_ram[2144] = 247;
    exp_54_ram[2145] = 0;
    exp_54_ram[2146] = 0;
    exp_54_ram[2147] = 0;
    exp_54_ram[2148] = 205;
    exp_54_ram[2149] = 254;
    exp_54_ram[2150] = 254;
    exp_54_ram[2151] = 5;
    exp_54_ram[2152] = 254;
    exp_54_ram[2153] = 255;
    exp_54_ram[2154] = 0;
    exp_54_ram[2155] = 248;
    exp_54_ram[2156] = 0;
    exp_54_ram[2157] = 254;
    exp_54_ram[2158] = 255;
    exp_54_ram[2159] = 0;
    exp_54_ram[2160] = 241;
    exp_54_ram[2161] = 0;
    exp_54_ram[2162] = 254;
    exp_54_ram[2163] = 0;
    exp_54_ram[2164] = 0;
    exp_54_ram[2165] = 103;
    exp_54_ram[2166] = 231;
    exp_54_ram[2167] = 16;
    exp_54_ram[2168] = 254;
    exp_54_ram[2169] = 0;
    exp_54_ram[2170] = 254;
    exp_54_ram[2171] = 254;
    exp_54_ram[2172] = 6;
    exp_54_ram[2173] = 250;
    exp_54_ram[2174] = 104;
    exp_54_ram[2175] = 229;
    exp_54_ram[2176] = 254;
    exp_54_ram[2177] = 0;
    exp_54_ram[2178] = 254;
    exp_54_ram[2179] = 254;
    exp_54_ram[2180] = 0;
    exp_54_ram[2181] = 244;
    exp_54_ram[2182] = 1;
    exp_54_ram[2183] = 175;
    exp_54_ram[2184] = 0;
    exp_54_ram[2185] = 254;
    exp_54_ram[2186] = 2;
    exp_54_ram[2187] = 174;
    exp_54_ram[2188] = 0;
    exp_54_ram[2189] = 252;
    exp_54_ram[2190] = 4;
    exp_54_ram[2191] = 173;
    exp_54_ram[2192] = 0;
    exp_54_ram[2193] = 252;
    exp_54_ram[2194] = 252;
    exp_54_ram[2195] = 7;
    exp_54_ram[2196] = 254;
    exp_54_ram[2197] = 182;
    exp_54_ram[2198] = 4;
    exp_54_ram[2199] = 171;
    exp_54_ram[2200] = 0;
    exp_54_ram[2201] = 254;
    exp_54_ram[2202] = 253;
    exp_54_ram[2203] = 180;
    exp_54_ram[2204] = 2;
    exp_54_ram[2205] = 169;
    exp_54_ram[2206] = 0;
    exp_54_ram[2207] = 252;
    exp_54_ram[2208] = 253;
    exp_54_ram[2209] = 179;
    exp_54_ram[2210] = 1;
    exp_54_ram[2211] = 168;
    exp_54_ram[2212] = 0;
    exp_54_ram[2213] = 252;
    exp_54_ram[2214] = 254;
    exp_54_ram[2215] = 253;
    exp_54_ram[2216] = 253;
    exp_54_ram[2217] = 0;
    exp_54_ram[2218] = 0;
    exp_54_ram[2219] = 104;
    exp_54_ram[2220] = 161;
    exp_54_ram[2221] = 253;
    exp_54_ram[2222] = 0;
    exp_54_ram[2223] = 252;
    exp_54_ram[2224] = 253;
    exp_54_ram[2225] = 6;
    exp_54_ram[2226] = 248;
    exp_54_ram[2227] = 254;
    exp_54_ram[2228] = 174;
    exp_54_ram[2229] = 253;
    exp_54_ram[2230] = 174;
    exp_54_ram[2231] = 253;
    exp_54_ram[2232] = 173;
    exp_54_ram[2233] = 15;
    exp_54_ram[2234] = 15;
    exp_54_ram[2235] = 16;
    exp_54_ram[2236] = 0;
    exp_54_ram[2237] = 254;
    exp_54_ram[2238] = 0;
    exp_54_ram[2239] = 0;
    exp_54_ram[2240] = 2;
    exp_54_ram[2241] = 106;
    exp_54_ram[2242] = 212;
    exp_54_ram[2243] = 107;
    exp_54_ram[2244] = 211;
    exp_54_ram[2245] = 108;
    exp_54_ram[2246] = 211;
    exp_54_ram[2247] = 109;
    exp_54_ram[2248] = 210;
    exp_54_ram[2249] = 110;
    exp_54_ram[2250] = 210;
    exp_54_ram[2251] = 112;
    exp_54_ram[2252] = 209;
    exp_54_ram[2253] = 206;
    exp_54_ram[2254] = 0;
    exp_54_ram[2255] = 254;
    exp_54_ram[2256] = 254;
    exp_54_ram[2257] = 249;
    exp_54_ram[2258] = 0;
    exp_54_ram[2259] = 250;
    exp_54_ram[2260] = 0;
    exp_54_ram[2261] = 0;
    exp_54_ram[2262] = 66;
    exp_54_ram[2263] = 0;
    exp_54_ram[2264] = 0;
    exp_54_ram[2265] = 0;
    exp_54_ram[2266] = 230;
    exp_54_ram[2267] = 2;
    exp_54_ram[2268] = 232;
    exp_54_ram[2269] = 1;
    exp_54_ram[2270] = 248;
    exp_54_ram[2271] = 1;
    exp_54_ram[2272] = 132;
    exp_54_ram[2273] = 0;
    exp_54_ram[2274] = 216;
    exp_54_ram[2275] = 0;
    exp_54_ram[2276] = 247;
    exp_54_ram[2277] = 0;
    exp_54_ram[2278] = 0;
    exp_54_ram[2279] = 2;
    exp_54_ram[2280] = 255;
    exp_54_ram[2281] = 2;
    exp_54_ram[2282] = 0;
    exp_54_ram[2283] = 0;
    exp_54_ram[2284] = 0;
    exp_54_ram[2285] = 64;
    exp_54_ram[2286] = 1;
    exp_54_ram[2287] = 0;
    exp_54_ram[2288] = 254;
    exp_54_ram[2289] = 255;
    exp_54_ram[2290] = 0;
    exp_54_ram[2291] = 254;
    exp_54_ram[2292] = 2;
    exp_54_ram[2293] = 0;
    exp_54_ram[2294] = 128;
    exp_54_ram[2295] = 128;
    exp_54_ram[2296] = 128;
    exp_54_ram[2297] = 77;
    exp_54_ram[2298] = 117;
    exp_54_ram[2299] = 100;
    exp_54_ram[2300] = 70;
    exp_54_ram[2301] = 97;
    exp_54_ram[2302] = 0;
    exp_54_ram[2303] = 70;
    exp_54_ram[2304] = 97;
    exp_54_ram[2305] = 114;
    exp_54_ram[2306] = 74;
    exp_54_ram[2307] = 117;
    exp_54_ram[2308] = 103;
    exp_54_ram[2309] = 79;
    exp_54_ram[2310] = 111;
    exp_54_ram[2311] = 99;
    exp_54_ram[2312] = 0;
    exp_54_ram[2313] = 0;
    exp_54_ram[2314] = 0;
    exp_54_ram[2315] = 0;
    exp_54_ram[2316] = 0;
    exp_54_ram[2317] = 0;
    exp_54_ram[2318] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_252;
  assign exp_252 = exp_533;

  reg [3:0] exp_533_reg;
  always@(*) begin
    case (exp_385)
      0:exp_533_reg <= exp_520;
      1:exp_533_reg <= exp_525;
      2:exp_533_reg <= exp_526;
      3:exp_533_reg <= exp_527;
      4:exp_533_reg <= exp_528;
      5:exp_533_reg <= exp_529;
      6:exp_533_reg <= exp_530;
      7:exp_533_reg <= exp_531;
      default:exp_533_reg <= exp_532;
    endcase
  end
  assign exp_533 = exp_533_reg;
  assign exp_532 = 0;
  assign exp_520 = exp_516 << exp_519;
  assign exp_516 = 1;
  assign exp_519 = exp_518 + exp_517;
  assign exp_518 = 0;
  assign exp_517 = exp_453[1:0];
  assign exp_525 = exp_521 << exp_524;
  assign exp_521 = 3;
  assign exp_524 = exp_523 + exp_522;
  assign exp_523 = 0;
  assign exp_522 = exp_453[1:1];
  assign exp_526 = 15;
  assign exp_527 = 0;
  assign exp_528 = 0;
  assign exp_529 = 0;
  assign exp_530 = 0;
  assign exp_531 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_247;
  assign exp_247 = exp_515;

  reg [31:0] exp_515_reg;
  always@(*) begin
    case (exp_385)
      0:exp_515_reg <= exp_502;
      1:exp_515_reg <= exp_506;
      2:exp_515_reg <= exp_508;
      3:exp_515_reg <= exp_509;
      4:exp_515_reg <= exp_510;
      5:exp_515_reg <= exp_511;
      6:exp_515_reg <= exp_512;
      7:exp_515_reg <= exp_513;
      default:exp_515_reg <= exp_514;
    endcase
  end
  assign exp_515 = exp_515_reg;
  assign exp_514 = 0;

  reg [31:0] exp_502_reg;
  always@(*) begin
    case (exp_456)
      0:exp_502_reg <= exp_488;
      1:exp_502_reg <= exp_496;
      2:exp_502_reg <= exp_498;
      3:exp_502_reg <= exp_500;
      default:exp_502_reg <= exp_501;
    endcase
  end
  assign exp_502 = exp_502_reg;
  assign exp_501 = 0;
  assign exp_488 = exp_487;
  assign exp_487 = exp_486 + exp_485;
  assign exp_486 = 0;
  assign exp_485 = exp_375[7:0];

      reg [31:0] exp_375_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_375_reg <= exp_318;
        end
      end
      assign exp_375 = exp_375_reg;
      assign exp_496 = exp_488 << exp_495;
  assign exp_495 = 8;
  assign exp_498 = exp_488 << exp_497;
  assign exp_497 = 16;
  assign exp_500 = exp_488 << exp_499;
  assign exp_499 = 24;

  reg [31:0] exp_506_reg;
  always@(*) begin
    case (exp_459)
      0:exp_506_reg <= exp_492;
      1:exp_506_reg <= exp_504;
      default:exp_506_reg <= exp_505;
    endcase
  end
  assign exp_506 = exp_506_reg;
  assign exp_459 = exp_458 + exp_457;
  assign exp_458 = 0;
  assign exp_457 = exp_453[1:1];
  assign exp_505 = 0;
  assign exp_492 = exp_491;
  assign exp_491 = exp_490 + exp_489;
  assign exp_490 = 0;
  assign exp_489 = exp_375[15:0];
  assign exp_504 = exp_492 << exp_503;
  assign exp_503 = 16;
  assign exp_508 = exp_507 + exp_494;
  assign exp_507 = 0;
  assign exp_494 = exp_493 + exp_375;
  assign exp_493 = 0;
  assign exp_509 = 0;
  assign exp_510 = 0;
  assign exp_511 = 0;
  assign exp_512 = 0;
  assign exp_513 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 0;
    exp_47_ram[32] = 193;
    exp_47_ram[33] = 0;
    exp_47_ram[34] = 0;
    exp_47_ram[35] = 5;
    exp_47_ram[36] = 5;
    exp_47_ram[37] = 6;
    exp_47_ram[38] = 6;
    exp_47_ram[39] = 8;
    exp_47_ram[40] = 6;
    exp_47_ram[41] = 0;
    exp_47_ram[42] = 197;
    exp_47_ram[43] = 1;
    exp_47_ram[44] = 230;
    exp_47_ram[45] = 240;
    exp_47_ram[46] = 199;
    exp_47_ram[47] = 55;
    exp_47_ram[48] = 230;
    exp_47_ram[49] = 166;
    exp_47_ram[50] = 6;
    exp_47_ram[51] = 0;
    exp_47_ram[52] = 230;
    exp_47_ram[53] = 229;
    exp_47_ram[54] = 229;
    exp_47_ram[55] = 215;
    exp_47_ram[56] = 232;
    exp_47_ram[57] = 214;
    exp_47_ram[58] = 183;
    exp_47_ram[59] = 216;
    exp_47_ram[60] = 8;
    exp_47_ram[61] = 21;
    exp_47_ram[62] = 8;
    exp_47_ram[63] = 6;
    exp_47_ram[64] = 3;
    exp_47_ram[65] = 21;
    exp_47_ram[66] = 6;
    exp_47_ram[67] = 214;
    exp_47_ram[68] = 7;
    exp_47_ram[69] = 247;
    exp_47_ram[70] = 183;
    exp_47_ram[71] = 7;
    exp_47_ram[72] = 246;
    exp_47_ram[73] = 7;
    exp_47_ram[74] = 183;
    exp_47_ram[75] = 230;
    exp_47_ram[76] = 7;
    exp_47_ram[77] = 183;
    exp_47_ram[78] = 23;
    exp_47_ram[79] = 3;
    exp_47_ram[80] = 3;
    exp_47_ram[81] = 23;
    exp_47_ram[82] = 7;
    exp_47_ram[83] = 103;
    exp_47_ram[84] = 246;
    exp_47_ram[85] = 7;
    exp_47_ram[86] = 211;
    exp_47_ram[87] = 104;
    exp_47_ram[88] = 247;
    exp_47_ram[89] = 3;
    exp_47_ram[90] = 211;
    exp_47_ram[91] = 231;
    exp_47_ram[92] = 5;
    exp_47_ram[93] = 197;
    exp_47_ram[94] = 0;
    exp_47_ram[95] = 64;
    exp_47_ram[96] = 0;
    exp_47_ram[97] = 0;
    exp_47_ram[98] = 166;
    exp_47_ram[99] = 128;
    exp_47_ram[100] = 31;
    exp_47_ram[101] = 6;
    exp_47_ram[102] = 16;
    exp_47_ram[103] = 199;
    exp_47_ram[104] = 1;
    exp_47_ram[105] = 232;
    exp_47_ram[106] = 240;
    exp_47_ram[107] = 7;
    exp_47_ram[108] = 128;
    exp_47_ram[109] = 168;
    exp_47_ram[110] = 230;
    exp_47_ram[111] = 6;
    exp_47_ram[112] = 0;
    exp_47_ram[113] = 167;
    exp_47_ram[114] = 230;
    exp_47_ram[115] = 230;
    exp_47_ram[116] = 7;
    exp_47_ram[117] = 16;
    exp_47_ram[118] = 8;
    exp_47_ram[119] = 8;
    exp_47_ram[120] = 6;
    exp_47_ram[121] = 3;
    exp_47_ram[122] = 23;
    exp_47_ram[123] = 23;
    exp_47_ram[124] = 6;
    exp_47_ram[125] = 230;
    exp_47_ram[126] = 246;
    exp_47_ram[127] = 7;
    exp_47_ram[128] = 199;
    exp_47_ram[129] = 7;
    exp_47_ram[130] = 247;
    exp_47_ram[131] = 7;
    exp_47_ram[132] = 199;
    exp_47_ram[133] = 231;
    exp_47_ram[134] = 7;
    exp_47_ram[135] = 199;
    exp_47_ram[136] = 23;
    exp_47_ram[137] = 3;
    exp_47_ram[138] = 3;
    exp_47_ram[139] = 23;
    exp_47_ram[140] = 7;
    exp_47_ram[141] = 103;
    exp_47_ram[142] = 230;
    exp_47_ram[143] = 7;
    exp_47_ram[144] = 211;
    exp_47_ram[145] = 104;
    exp_47_ram[146] = 247;
    exp_47_ram[147] = 3;
    exp_47_ram[148] = 211;
    exp_47_ram[149] = 231;
    exp_47_ram[150] = 5;
    exp_47_ram[151] = 197;
    exp_47_ram[152] = 0;
    exp_47_ram[153] = 0;
    exp_47_ram[154] = 0;
    exp_47_ram[155] = 232;
    exp_47_ram[156] = 128;
    exp_47_ram[157] = 31;
    exp_47_ram[158] = 216;
    exp_47_ram[159] = 231;
    exp_47_ram[160] = 216;
    exp_47_ram[161] = 215;
    exp_47_ram[162] = 232;
    exp_47_ram[163] = 8;
    exp_47_ram[164] = 247;
    exp_47_ram[165] = 21;
    exp_47_ram[166] = 8;
    exp_47_ram[167] = 7;
    exp_47_ram[168] = 6;
    exp_47_ram[169] = 21;
    exp_47_ram[170] = 7;
    exp_47_ram[171] = 183;
    exp_47_ram[172] = 167;
    exp_47_ram[173] = 5;
    exp_47_ram[174] = 215;
    exp_47_ram[175] = 7;
    exp_47_ram[176] = 245;
    exp_47_ram[177] = 7;
    exp_47_ram[178] = 215;
    exp_47_ram[179] = 229;
    exp_47_ram[180] = 7;
    exp_47_ram[181] = 215;
    exp_47_ram[182] = 22;
    exp_47_ram[183] = 6;
    exp_47_ram[184] = 6;
    exp_47_ram[185] = 22;
    exp_47_ram[186] = 7;
    exp_47_ram[187] = 215;
    exp_47_ram[188] = 199;
    exp_47_ram[189] = 6;
    exp_47_ram[190] = 167;
    exp_47_ram[191] = 7;
    exp_47_ram[192] = 246;
    exp_47_ram[193] = 7;
    exp_47_ram[194] = 167;
    exp_47_ram[195] = 230;
    exp_47_ram[196] = 7;
    exp_47_ram[197] = 5;
    exp_47_ram[198] = 167;
    exp_47_ram[199] = 229;
    exp_47_ram[200] = 159;
    exp_47_ram[201] = 213;
    exp_47_ram[202] = 1;
    exp_47_ram[203] = 230;
    exp_47_ram[204] = 240;
    exp_47_ram[205] = 215;
    exp_47_ram[206] = 53;
    exp_47_ram[207] = 182;
    exp_47_ram[208] = 0;
    exp_47_ram[209] = 167;
    exp_47_ram[210] = 7;
    exp_47_ram[211] = 0;
    exp_47_ram[212] = 183;
    exp_47_ram[213] = 229;
    exp_47_ram[214] = 229;
    exp_47_ram[215] = 16;
    exp_47_ram[216] = 246;
    exp_47_ram[217] = 200;
    exp_47_ram[218] = 21;
    exp_47_ram[219] = 95;
    exp_47_ram[220] = 0;
    exp_47_ram[221] = 0;
    exp_47_ram[222] = 230;
    exp_47_ram[223] = 128;
    exp_47_ram[224] = 223;
    exp_47_ram[225] = 230;
    exp_47_ram[226] = 182;
    exp_47_ram[227] = 216;
    exp_47_ram[228] = 231;
    exp_47_ram[229] = 8;
    exp_47_ram[230] = 222;
    exp_47_ram[231] = 183;
    exp_47_ram[232] = 232;
    exp_47_ram[233] = 182;
    exp_47_ram[234] = 247;
    exp_47_ram[235] = 8;
    exp_47_ram[236] = 7;
    exp_47_ram[237] = 6;
    exp_47_ram[238] = 222;
    exp_47_ram[239] = 6;
    exp_47_ram[240] = 230;
    exp_47_ram[241] = 199;
    exp_47_ram[242] = 14;
    exp_47_ram[243] = 231;
    exp_47_ram[244] = 7;
    exp_47_ram[245] = 254;
    exp_47_ram[246] = 7;
    exp_47_ram[247] = 231;
    exp_47_ram[248] = 238;
    exp_47_ram[249] = 7;
    exp_47_ram[250] = 231;
    exp_47_ram[251] = 215;
    exp_47_ram[252] = 215;
    exp_47_ram[253] = 6;
    exp_47_ram[254] = 231;
    exp_47_ram[255] = 6;
    exp_47_ram[256] = 7;
    exp_47_ram[257] = 246;
    exp_47_ram[258] = 7;
    exp_47_ram[259] = 199;
    exp_47_ram[260] = 7;
    exp_47_ram[261] = 247;
    exp_47_ram[262] = 7;
    exp_47_ram[263] = 199;
    exp_47_ram[264] = 231;
    exp_47_ram[265] = 7;
    exp_47_ram[266] = 5;
    exp_47_ram[267] = 1;
    exp_47_ram[268] = 197;
    exp_47_ram[269] = 254;
    exp_47_ram[270] = 213;
    exp_47_ram[271] = 5;
    exp_47_ram[272] = 211;
    exp_47_ram[273] = 3;
    exp_47_ram[274] = 199;
    exp_47_ram[275] = 216;
    exp_47_ram[276] = 214;
    exp_47_ram[277] = 14;
    exp_47_ram[278] = 104;
    exp_47_ram[279] = 216;
    exp_47_ram[280] = 7;
    exp_47_ram[281] = 102;
    exp_47_ram[282] = 215;
    exp_47_ram[283] = 214;
    exp_47_ram[284] = 7;
    exp_47_ram[285] = 198;
    exp_47_ram[286] = 199;
    exp_47_ram[287] = 199;
    exp_47_ram[288] = 1;
    exp_47_ram[289] = 247;
    exp_47_ram[290] = 247;
    exp_47_ram[291] = 7;
    exp_47_ram[292] = 254;
    exp_47_ram[293] = 184;
    exp_47_ram[294] = 199;
    exp_47_ram[295] = 0;
    exp_47_ram[296] = 232;
    exp_47_ram[297] = 245;
    exp_47_ram[298] = 31;
    exp_47_ram[299] = 0;
    exp_47_ram[300] = 0;
    exp_47_ram[301] = 223;
    exp_47_ram[302] = 5;
    exp_47_ram[303] = 0;
    exp_47_ram[304] = 21;
    exp_47_ram[305] = 6;
    exp_47_ram[306] = 197;
    exp_47_ram[307] = 21;
    exp_47_ram[308] = 22;
    exp_47_ram[309] = 5;
    exp_47_ram[310] = 0;
    exp_47_ram[311] = 5;
    exp_47_ram[312] = 5;
    exp_47_ram[313] = 5;
    exp_47_ram[314] = 5;
    exp_47_ram[315] = 240;
    exp_47_ram[316] = 6;
    exp_47_ram[317] = 16;
    exp_47_ram[318] = 182;
    exp_47_ram[319] = 192;
    exp_47_ram[320] = 22;
    exp_47_ram[321] = 22;
    exp_47_ram[322] = 182;
    exp_47_ram[323] = 0;
    exp_47_ram[324] = 197;
    exp_47_ram[325] = 197;
    exp_47_ram[326] = 213;
    exp_47_ram[327] = 22;
    exp_47_ram[328] = 22;
    exp_47_ram[329] = 6;
    exp_47_ram[330] = 0;
    exp_47_ram[331] = 0;
    exp_47_ram[332] = 95;
    exp_47_ram[333] = 5;
    exp_47_ram[334] = 2;
    exp_47_ram[335] = 160;
    exp_47_ram[336] = 176;
    exp_47_ram[337] = 176;
    exp_47_ram[338] = 223;
    exp_47_ram[339] = 176;
    exp_47_ram[340] = 0;
    exp_47_ram[341] = 31;
    exp_47_ram[342] = 160;
    exp_47_ram[343] = 2;
    exp_47_ram[344] = 0;
    exp_47_ram[345] = 5;
    exp_47_ram[346] = 5;
    exp_47_ram[347] = 159;
    exp_47_ram[348] = 5;
    exp_47_ram[349] = 2;
    exp_47_ram[350] = 176;
    exp_47_ram[351] = 5;
    exp_47_ram[352] = 160;
    exp_47_ram[353] = 31;
    exp_47_ram[354] = 176;
    exp_47_ram[355] = 2;
    exp_47_ram[356] = 108;
    exp_47_ram[357] = 87;
    exp_47_ram[358] = 100;
    exp_47_ram[359] = 0;
    exp_47_ram[360] = 110;
    exp_47_ram[361] = 103;
    exp_47_ram[362] = 105;
    exp_47_ram[363] = 32;
    exp_47_ram[364] = 101;
    exp_47_ram[365] = 101;
    exp_47_ram[366] = 46;
    exp_47_ram[367] = 0;
    exp_47_ram[368] = 10;
    exp_47_ram[369] = 32;
    exp_47_ram[370] = 98;
    exp_47_ram[371] = 105;
    exp_47_ram[372] = 103;
    exp_47_ram[373] = 109;
    exp_47_ram[374] = 105;
    exp_47_ram[375] = 101;
    exp_47_ram[376] = 110;
    exp_47_ram[377] = 115;
    exp_47_ram[378] = 110;
    exp_47_ram[379] = 0;
    exp_47_ram[380] = 32;
    exp_47_ram[381] = 98;
    exp_47_ram[382] = 105;
    exp_47_ram[383] = 103;
    exp_47_ram[384] = 109;
    exp_47_ram[385] = 105;
    exp_47_ram[386] = 101;
    exp_47_ram[387] = 110;
    exp_47_ram[388] = 115;
    exp_47_ram[389] = 110;
    exp_47_ram[390] = 0;
    exp_47_ram[391] = 32;
    exp_47_ram[392] = 98;
    exp_47_ram[393] = 105;
    exp_47_ram[394] = 103;
    exp_47_ram[395] = 100;
    exp_47_ram[396] = 100;
    exp_47_ram[397] = 105;
    exp_47_ram[398] = 32;
    exp_47_ram[399] = 111;
    exp_47_ram[400] = 0;
    exp_47_ram[401] = 32;
    exp_47_ram[402] = 98;
    exp_47_ram[403] = 105;
    exp_47_ram[404] = 103;
    exp_47_ram[405] = 100;
    exp_47_ram[406] = 100;
    exp_47_ram[407] = 105;
    exp_47_ram[408] = 32;
    exp_47_ram[409] = 111;
    exp_47_ram[410] = 0;
    exp_47_ram[411] = 105;
    exp_47_ram[412] = 101;
    exp_47_ram[413] = 37;
    exp_47_ram[414] = 46;
    exp_47_ram[415] = 105;
    exp_47_ram[416] = 0;
    exp_47_ram[417] = 115;
    exp_47_ram[418] = 0;
    exp_47_ram[419] = 108;
    exp_47_ram[420] = 116;
    exp_47_ram[421] = 37;
    exp_47_ram[422] = 32;
    exp_47_ram[423] = 120;
    exp_47_ram[424] = 56;
    exp_47_ram[425] = 0;
    exp_47_ram[426] = 104;
    exp_47_ram[427] = 45;
    exp_47_ram[428] = 101;
    exp_47_ram[429] = 0;
    exp_47_ram[430] = 41;
    exp_47_ram[431] = 108;
    exp_47_ram[432] = 87;
    exp_47_ram[433] = 100;
    exp_47_ram[434] = 32;
    exp_47_ram[435] = 103;
    exp_47_ram[436] = 82;
    exp_47_ram[437] = 114;
    exp_47_ram[438] = 32;
    exp_47_ram[439] = 112;
    exp_47_ram[440] = 116;
    exp_47_ram[441] = 0;
    exp_47_ram[442] = 32;
    exp_47_ram[443] = 116;
    exp_47_ram[444] = 108;
    exp_47_ram[445] = 108;
    exp_47_ram[446] = 116;
    exp_47_ram[447] = 0;
    exp_47_ram[448] = 32;
    exp_47_ram[449] = 116;
    exp_47_ram[450] = 109;
    exp_47_ram[451] = 0;
    exp_47_ram[452] = 2;
    exp_47_ram[453] = 3;
    exp_47_ram[454] = 4;
    exp_47_ram[455] = 4;
    exp_47_ram[456] = 5;
    exp_47_ram[457] = 5;
    exp_47_ram[458] = 5;
    exp_47_ram[459] = 5;
    exp_47_ram[460] = 6;
    exp_47_ram[461] = 6;
    exp_47_ram[462] = 6;
    exp_47_ram[463] = 6;
    exp_47_ram[464] = 6;
    exp_47_ram[465] = 6;
    exp_47_ram[466] = 6;
    exp_47_ram[467] = 6;
    exp_47_ram[468] = 7;
    exp_47_ram[469] = 7;
    exp_47_ram[470] = 7;
    exp_47_ram[471] = 7;
    exp_47_ram[472] = 7;
    exp_47_ram[473] = 7;
    exp_47_ram[474] = 7;
    exp_47_ram[475] = 7;
    exp_47_ram[476] = 7;
    exp_47_ram[477] = 7;
    exp_47_ram[478] = 7;
    exp_47_ram[479] = 7;
    exp_47_ram[480] = 7;
    exp_47_ram[481] = 7;
    exp_47_ram[482] = 7;
    exp_47_ram[483] = 7;
    exp_47_ram[484] = 8;
    exp_47_ram[485] = 8;
    exp_47_ram[486] = 8;
    exp_47_ram[487] = 8;
    exp_47_ram[488] = 8;
    exp_47_ram[489] = 8;
    exp_47_ram[490] = 8;
    exp_47_ram[491] = 8;
    exp_47_ram[492] = 8;
    exp_47_ram[493] = 8;
    exp_47_ram[494] = 8;
    exp_47_ram[495] = 8;
    exp_47_ram[496] = 8;
    exp_47_ram[497] = 8;
    exp_47_ram[498] = 8;
    exp_47_ram[499] = 8;
    exp_47_ram[500] = 8;
    exp_47_ram[501] = 8;
    exp_47_ram[502] = 8;
    exp_47_ram[503] = 8;
    exp_47_ram[504] = 8;
    exp_47_ram[505] = 8;
    exp_47_ram[506] = 8;
    exp_47_ram[507] = 8;
    exp_47_ram[508] = 8;
    exp_47_ram[509] = 8;
    exp_47_ram[510] = 8;
    exp_47_ram[511] = 8;
    exp_47_ram[512] = 8;
    exp_47_ram[513] = 8;
    exp_47_ram[514] = 8;
    exp_47_ram[515] = 8;
    exp_47_ram[516] = 165;
    exp_47_ram[517] = 0;
    exp_47_ram[518] = 0;
    exp_47_ram[519] = 7;
    exp_47_ram[520] = 7;
    exp_47_ram[521] = 0;
    exp_47_ram[522] = 5;
    exp_47_ram[523] = 0;
    exp_47_ram[524] = 167;
    exp_47_ram[525] = 7;
    exp_47_ram[526] = 7;
    exp_47_ram[527] = 0;
    exp_47_ram[528] = 21;
    exp_47_ram[529] = 229;
    exp_47_ram[530] = 159;
    exp_47_ram[531] = 1;
    exp_47_ram[532] = 0;
    exp_47_ram[533] = 129;
    exp_47_ram[534] = 135;
    exp_47_ram[535] = 17;
    exp_47_ram[536] = 4;
    exp_47_ram[537] = 95;
    exp_47_ram[538] = 160;
    exp_47_ram[539] = 193;
    exp_47_ram[540] = 244;
    exp_47_ram[541] = 129;
    exp_47_ram[542] = 0;
    exp_47_ram[543] = 1;
    exp_47_ram[544] = 0;
    exp_47_ram[545] = 1;
    exp_47_ram[546] = 129;
    exp_47_ram[547] = 17;
    exp_47_ram[548] = 22;
    exp_47_ram[549] = 5;
    exp_47_ram[550] = 159;
    exp_47_ram[551] = 193;
    exp_47_ram[552] = 4;
    exp_47_ram[553] = 129;
    exp_47_ram[554] = 1;
    exp_47_ram[555] = 0;
    exp_47_ram[556] = 214;
    exp_47_ram[557] = 166;
    exp_47_ram[558] = 134;
    exp_47_ram[559] = 6;
    exp_47_ram[560] = 223;
    exp_47_ram[561] = 1;
    exp_47_ram[562] = 129;
    exp_47_ram[563] = 145;
    exp_47_ram[564] = 33;
    exp_47_ram[565] = 49;
    exp_47_ram[566] = 65;
    exp_47_ram[567] = 129;
    exp_47_ram[568] = 145;
    exp_47_ram[569] = 7;
    exp_47_ram[570] = 17;
    exp_47_ram[571] = 81;
    exp_47_ram[572] = 97;
    exp_47_ram[573] = 113;
    exp_47_ram[574] = 161;
    exp_47_ram[575] = 177;
    exp_47_ram[576] = 128;
    exp_47_ram[577] = 5;
    exp_47_ram[578] = 5;
    exp_47_ram[579] = 6;
    exp_47_ram[580] = 6;
    exp_47_ram[581] = 7;
    exp_47_ram[582] = 8;
    exp_47_ram[583] = 8;
    exp_47_ram[584] = 248;
    exp_47_ram[585] = 0;
    exp_47_ram[586] = 248;
    exp_47_ram[587] = 128;
    exp_47_ram[588] = 0;
    exp_47_ram[589] = 0;
    exp_47_ram[590] = 144;
    exp_47_ram[591] = 16;
    exp_47_ram[592] = 128;
    exp_47_ram[593] = 7;
    exp_47_ram[594] = 124;
    exp_47_ram[595] = 247;
    exp_47_ram[596] = 3;
    exp_47_ram[597] = 13;
    exp_47_ram[598] = 93;
    exp_47_ram[599] = 247;
    exp_47_ram[600] = 251;
    exp_47_ram[601] = 3;
    exp_47_ram[602] = 243;
    exp_47_ram[603] = 5;
    exp_47_ram[604] = 4;
    exp_47_ram[605] = 4;
    exp_47_ram[606] = 3;
    exp_47_ram[607] = 159;
    exp_47_ram[608] = 16;
    exp_47_ram[609] = 124;
    exp_47_ram[610] = 253;
    exp_47_ram[611] = 139;
    exp_47_ram[612] = 139;
    exp_47_ram[613] = 193;
    exp_47_ram[614] = 129;
    exp_47_ram[615] = 65;
    exp_47_ram[616] = 1;
    exp_47_ram[617] = 193;
    exp_47_ram[618] = 129;
    exp_47_ram[619] = 65;
    exp_47_ram[620] = 1;
    exp_47_ram[621] = 193;
    exp_47_ram[622] = 129;
    exp_47_ram[623] = 65;
    exp_47_ram[624] = 1;
    exp_47_ram[625] = 193;
    exp_47_ram[626] = 1;
    exp_47_ram[627] = 0;
    exp_47_ram[628] = 10;
    exp_47_ram[629] = 115;
    exp_47_ram[630] = 31;
    exp_47_ram[631] = 115;
    exp_47_ram[632] = 159;
    exp_47_ram[633] = 169;
    exp_47_ram[634] = 5;
    exp_47_ram[635] = 4;
    exp_47_ram[636] = 4;
    exp_47_ram[637] = 9;
    exp_47_ram[638] = 223;
    exp_47_ram[639] = 159;
    exp_47_ram[640] = 160;
    exp_47_ram[641] = 0;
    exp_47_ram[642] = 223;
    exp_47_ram[643] = 154;
    exp_47_ram[644] = 160;
    exp_47_ram[645] = 11;
    exp_47_ram[646] = 160;
    exp_47_ram[647] = 159;
    exp_47_ram[648] = 6;
    exp_47_ram[649] = 7;
    exp_47_ram[650] = 1;
    exp_47_ram[651] = 129;
    exp_47_ram[652] = 145;
    exp_47_ram[653] = 49;
    exp_47_ram[654] = 81;
    exp_47_ram[655] = 97;
    exp_47_ram[656] = 113;
    exp_47_ram[657] = 145;
    exp_47_ram[658] = 161;
    exp_47_ram[659] = 177;
    exp_47_ram[660] = 6;
    exp_47_ram[661] = 17;
    exp_47_ram[662] = 33;
    exp_47_ram[663] = 65;
    exp_47_ram[664] = 129;
    exp_47_ram[665] = 5;
    exp_47_ram[666] = 5;
    exp_47_ram[667] = 6;
    exp_47_ram[668] = 0;
    exp_47_ram[669] = 0;
    exp_47_ram[670] = 80;
    exp_47_ram[671] = 144;
    exp_47_ram[672] = 160;
    exp_47_ram[673] = 144;
    exp_47_ram[674] = 80;
    exp_47_ram[675] = 233;
    exp_47_ram[676] = 7;
    exp_47_ram[677] = 23;
    exp_47_ram[678] = 41;
    exp_47_ram[679] = 85;
    exp_47_ram[680] = 10;
    exp_47_ram[681] = 7;
    exp_47_ram[682] = 0;
    exp_47_ram[683] = 215;
    exp_47_ram[684] = 39;
    exp_47_ram[685] = 41;
    exp_47_ram[686] = 7;
    exp_47_ram[687] = 7;
    exp_47_ram[688] = 193;
    exp_47_ram[689] = 129;
    exp_47_ram[690] = 65;
    exp_47_ram[691] = 1;
    exp_47_ram[692] = 193;
    exp_47_ram[693] = 129;
    exp_47_ram[694] = 65;
    exp_47_ram[695] = 1;
    exp_47_ram[696] = 193;
    exp_47_ram[697] = 129;
    exp_47_ram[698] = 65;
    exp_47_ram[699] = 1;
    exp_47_ram[700] = 193;
    exp_47_ram[701] = 6;
    exp_47_ram[702] = 1;
    exp_47_ram[703] = 0;
    exp_47_ram[704] = 6;
    exp_47_ram[705] = 4;
    exp_47_ram[706] = 4;
    exp_47_ram[707] = 159;
    exp_47_ram[708] = 5;
    exp_47_ram[709] = 10;
    exp_47_ram[710] = 7;
    exp_47_ram[711] = 9;
    exp_47_ram[712] = 223;
    exp_47_ram[713] = 0;
    exp_47_ram[714] = 0;
    exp_47_ram[715] = 41;
    exp_47_ram[716] = 6;
    exp_47_ram[717] = 25;
    exp_47_ram[718] = 41;
    exp_47_ram[719] = 6;
    exp_47_ram[720] = 189;
    exp_47_ram[721] = 102;
    exp_47_ram[722] = 219;
    exp_47_ram[723] = 48;
    exp_47_ram[724] = 182;
    exp_47_ram[725] = 213;
    exp_47_ram[726] = 86;
    exp_47_ram[727] = 128;
    exp_47_ram[728] = 182;
    exp_47_ram[729] = 76;
    exp_47_ram[730] = 16;
    exp_47_ram[731] = 64;
    exp_47_ram[732] = 183;
    exp_47_ram[733] = 10;
    exp_47_ram[734] = 229;
    exp_47_ram[735] = 6;
    exp_47_ram[736] = 31;
    exp_47_ram[737] = 64;
    exp_47_ram[738] = 182;
    exp_47_ram[739] = 76;
    exp_47_ram[740] = 12;
    exp_47_ram[741] = 12;
    exp_47_ram[742] = 6;
    exp_47_ram[743] = 4;
    exp_47_ram[744] = 4;
    exp_47_ram[745] = 208;
    exp_47_ram[746] = 225;
    exp_47_ram[747] = 241;
    exp_47_ram[748] = 95;
    exp_47_ram[749] = 193;
    exp_47_ram[750] = 129;
    exp_47_ram[751] = 5;
    exp_47_ram[752] = 0;
    exp_47_ram[753] = 160;
    exp_47_ram[754] = 247;
    exp_47_ram[755] = 144;
    exp_47_ram[756] = 4;
    exp_47_ram[757] = 4;
    exp_47_ram[758] = 223;
    exp_47_ram[759] = 128;
    exp_47_ram[760] = 118;
    exp_47_ram[761] = 219;
    exp_47_ram[762] = 240;
    exp_47_ram[763] = 182;
    exp_47_ram[764] = 48;
    exp_47_ram[765] = 246;
    exp_47_ram[766] = 12;
    exp_47_ram[767] = 76;
    exp_47_ram[768] = 12;
    exp_47_ram[769] = 5;
    exp_47_ram[770] = 7;
    exp_47_ram[771] = 159;
    exp_47_ram[772] = 128;
    exp_47_ram[773] = 182;
    exp_47_ram[774] = 76;
    exp_47_ram[775] = 0;
    exp_47_ram[776] = 0;
    exp_47_ram[777] = 192;
    exp_47_ram[778] = 6;
    exp_47_ram[779] = 4;
    exp_47_ram[780] = 4;
    exp_47_ram[781] = 80;
    exp_47_ram[782] = 95;
    exp_47_ram[783] = 12;
    exp_47_ram[784] = 6;
    exp_47_ram[785] = 4;
    exp_47_ram[786] = 4;
    exp_47_ram[787] = 76;
    exp_47_ram[788] = 95;
    exp_47_ram[789] = 5;
    exp_47_ram[790] = 12;
    exp_47_ram[791] = 159;
    exp_47_ram[792] = 6;
    exp_47_ram[793] = 4;
    exp_47_ram[794] = 4;
    exp_47_ram[795] = 241;
    exp_47_ram[796] = 95;
    exp_47_ram[797] = 129;
    exp_47_ram[798] = 5;
    exp_47_ram[799] = 28;
    exp_47_ram[800] = 31;
    exp_47_ram[801] = 0;
    exp_47_ram[802] = 160;
    exp_47_ram[803] = 12;
    exp_47_ram[804] = 31;
    exp_47_ram[805] = 76;
    exp_47_ram[806] = 0;
    exp_47_ram[807] = 160;
    exp_47_ram[808] = 12;
    exp_47_ram[809] = 223;
    exp_47_ram[810] = 76;
    exp_47_ram[811] = 0;
    exp_47_ram[812] = 128;
    exp_47_ram[813] = 223;
    exp_47_ram[814] = 0;
    exp_47_ram[815] = 6;
    exp_47_ram[816] = 0;
    exp_47_ram[817] = 1;
    exp_47_ram[818] = 241;
    exp_47_ram[819] = 0;
    exp_47_ram[820] = 193;
    exp_47_ram[821] = 5;
    exp_47_ram[822] = 135;
    exp_47_ram[823] = 177;
    exp_47_ram[824] = 209;
    exp_47_ram[825] = 0;
    exp_47_ram[826] = 65;
    exp_47_ram[827] = 17;
    exp_47_ram[828] = 225;
    exp_47_ram[829] = 1;
    exp_47_ram[830] = 17;
    exp_47_ram[831] = 209;
    exp_47_ram[832] = 31;
    exp_47_ram[833] = 193;
    exp_47_ram[834] = 1;
    exp_47_ram[835] = 0;
    exp_47_ram[836] = 53;
    exp_47_ram[837] = 39;
    exp_47_ram[838] = 0;
    exp_47_ram[839] = 133;
    exp_47_ram[840] = 7;
    exp_47_ram[841] = 0;
    exp_47_ram[842] = 39;
    exp_47_ram[843] = 229;
    exp_47_ram[844] = 0;
    exp_47_ram[845] = 0;
    exp_47_ram[846] = 71;
    exp_47_ram[847] = 5;
    exp_47_ram[848] = 7;
    exp_47_ram[849] = 243;
    exp_47_ram[850] = 229;
    exp_47_ram[851] = 1;
    exp_47_ram[852] = 0;
    exp_47_ram[853] = 248;
    exp_47_ram[854] = 8;
    exp_47_ram[855] = 103;
    exp_47_ram[856] = 39;
    exp_47_ram[857] = 213;
    exp_47_ram[858] = 6;
    exp_47_ram[859] = 24;
    exp_47_ram[860] = 246;
    exp_47_ram[861] = 184;
    exp_47_ram[862] = 8;
    exp_47_ram[863] = 199;
    exp_47_ram[864] = 23;
    exp_47_ram[865] = 159;
    exp_47_ram[866] = 183;
    exp_47_ram[867] = 182;
    exp_47_ram[868] = 199;
    exp_47_ram[869] = 231;
    exp_47_ram[870] = 22;
    exp_47_ram[871] = 38;
    exp_47_ram[872] = 247;
    exp_47_ram[873] = 213;
    exp_47_ram[874] = 199;
    exp_47_ram[875] = 246;
    exp_47_ram[876] = 23;
    exp_47_ram[877] = 95;
    exp_47_ram[878] = 0;
    exp_47_ram[879] = 134;
    exp_47_ram[880] = 245;
    exp_47_ram[881] = 197;
    exp_47_ram[882] = 197;
    exp_47_ram[883] = 167;
    exp_47_ram[884] = 5;
    exp_47_ram[885] = 1;
    exp_47_ram[886] = 245;
    exp_47_ram[887] = 183;
    exp_47_ram[888] = 245;
    exp_47_ram[889] = 0;
    exp_47_ram[890] = 71;
    exp_47_ram[891] = 134;
    exp_47_ram[892] = 0;
    exp_47_ram[893] = 8;
    exp_47_ram[894] = 7;
    exp_47_ram[895] = 23;
    exp_47_ram[896] = 39;
    exp_47_ram[897] = 214;
    exp_47_ram[898] = 6;
    exp_47_ram[899] = 181;
    exp_47_ram[900] = 215;
    exp_47_ram[901] = 101;
    exp_47_ram[902] = 23;
    exp_47_ram[903] = 5;
    exp_47_ram[904] = 39;
    exp_47_ram[905] = 230;
    exp_47_ram[906] = 23;
    exp_47_ram[907] = 39;
    exp_47_ram[908] = 166;
    exp_47_ram[909] = 5;
    exp_47_ram[910] = 184;
    exp_47_ram[911] = 104;
    exp_47_ram[912] = 8;
    exp_47_ram[913] = 213;
    exp_47_ram[914] = 22;
    exp_47_ram[915] = 21;
    exp_47_ram[916] = 215;
    exp_47_ram[917] = 167;
    exp_47_ram[918] = 31;
    exp_47_ram[919] = 0;
    exp_47_ram[920] = 181;
    exp_47_ram[921] = 55;
    exp_47_ram[922] = 5;
    exp_47_ram[923] = 7;
    exp_47_ram[924] = 5;
    exp_47_ram[925] = 197;
    exp_47_ram[926] = 240;
    exp_47_ram[927] = 192;
    exp_47_ram[928] = 7;
    exp_47_ram[929] = 7;
    exp_47_ram[930] = 6;
    exp_47_ram[931] = 22;
    exp_47_ram[932] = 71;
    exp_47_ram[933] = 22;
    exp_47_ram[934] = 135;
    exp_47_ram[935] = 22;
    exp_47_ram[936] = 199;
    exp_47_ram[937] = 22;
    exp_47_ram[938] = 227;
    exp_47_ram[939] = 24;
    exp_47_ram[940] = 246;
    exp_47_ram[941] = 6;
    exp_47_ram[942] = 197;
    exp_47_ram[943] = 197;
    exp_47_ram[944] = 48;
    exp_47_ram[945] = 247;
    exp_47_ram[946] = 6;
    exp_47_ram[947] = 55;
    exp_47_ram[948] = 199;
    exp_47_ram[949] = 230;
    exp_47_ram[950] = 229;
    exp_47_ram[951] = 0;
    exp_47_ram[952] = 246;
    exp_47_ram[953] = 0;
    exp_47_ram[954] = 245;
    exp_47_ram[955] = 8;
    exp_47_ram[956] = 246;
    exp_47_ram[957] = 71;
    exp_47_ram[958] = 24;
    exp_47_ram[959] = 159;
    exp_47_ram[960] = 245;
    exp_47_ram[961] = 7;
    exp_47_ram[962] = 246;
    exp_47_ram[963] = 23;
    exp_47_ram[964] = 7;
    exp_47_ram[965] = 223;
    exp_47_ram[966] = 53;
    exp_47_ram[967] = 7;
    exp_47_ram[968] = 1;
    exp_47_ram[969] = 64;
    exp_47_ram[970] = 129;
    exp_47_ram[971] = 17;
    exp_47_ram[972] = 5;
    exp_47_ram[973] = 143;
    exp_47_ram[974] = 16;
    exp_47_ram[975] = 5;
    exp_47_ram[976] = 0;
    exp_47_ram[977] = 4;
    exp_47_ram[978] = 79;
    exp_47_ram[979] = 21;
    exp_47_ram[980] = 193;
    exp_47_ram[981] = 129;
    exp_47_ram[982] = 7;
    exp_47_ram[983] = 1;
    exp_47_ram[984] = 0;
    exp_47_ram[985] = 0;
    exp_47_ram[986] = 7;
    exp_47_ram[987] = 0;
    exp_47_ram[988] = 213;
    exp_47_ram[989] = 215;
    exp_47_ram[990] = 7;
    exp_47_ram[991] = 213;
    exp_47_ram[992] = 128;
    exp_47_ram[993] = 224;
    exp_47_ram[994] = 215;
    exp_47_ram[995] = 16;
    exp_47_ram[996] = 240;
    exp_47_ram[997] = 229;
    exp_47_ram[998] = 1;
    exp_47_ram[999] = 17;
    exp_47_ram[1000] = 159;
    exp_47_ram[1001] = 193;
    exp_47_ram[1002] = 160;
    exp_47_ram[1003] = 199;
    exp_47_ram[1004] = 7;
    exp_47_ram[1005] = 1;
    exp_47_ram[1006] = 0;
    exp_47_ram[1007] = 224;
    exp_47_ram[1008] = 7;
    exp_47_ram[1009] = 0;
    exp_47_ram[1010] = 0;
    exp_47_ram[1011] = 7;
    exp_47_ram[1012] = 71;
    exp_47_ram[1013] = 71;
    exp_47_ram[1014] = 6;
    exp_47_ram[1015] = 135;
    exp_47_ram[1016] = 213;
    exp_47_ram[1017] = 0;
    exp_47_ram[1018] = 1;
    exp_47_ram[1019] = 81;
    exp_47_ram[1020] = 69;
    exp_47_ram[1021] = 145;
    exp_47_ram[1022] = 1;
    exp_47_ram[1023] = 129;
    exp_47_ram[1024] = 33;
    exp_47_ram[1025] = 49;
    exp_47_ram[1026] = 65;
    exp_47_ram[1027] = 17;
    exp_47_ram[1028] = 97;
    exp_47_ram[1029] = 5;
    exp_47_ram[1030] = 32;
    exp_47_ram[1031] = 0;
    exp_47_ram[1032] = 0;
    exp_47_ram[1033] = 202;
    exp_47_ram[1034] = 4;
    exp_47_ram[1035] = 138;
    exp_47_ram[1036] = 10;
    exp_47_ram[1037] = 1;
    exp_47_ram[1038] = 0;
    exp_47_ram[1039] = 10;
    exp_47_ram[1040] = 155;
    exp_47_ram[1041] = 4;
    exp_47_ram[1042] = 4;
    exp_47_ram[1043] = 95;
    exp_47_ram[1044] = 10;
    exp_47_ram[1045] = 79;
    exp_47_ram[1046] = 169;
    exp_47_ram[1047] = 37;
    exp_47_ram[1048] = 55;
    exp_47_ram[1049] = 5;
    exp_47_ram[1050] = 20;
    exp_47_ram[1051] = 95;
    exp_47_ram[1052] = 4;
    exp_47_ram[1053] = 95;
    exp_47_ram[1054] = 160;
    exp_47_ram[1055] = 4;
    exp_47_ram[1056] = 213;
    exp_47_ram[1057] = 79;
    exp_47_ram[1058] = 169;
    exp_47_ram[1059] = 37;
    exp_47_ram[1060] = 55;
    exp_47_ram[1061] = 5;
    exp_47_ram[1062] = 20;
    exp_47_ram[1063] = 31;
    exp_47_ram[1064] = 138;
    exp_47_ram[1065] = 74;
    exp_47_ram[1066] = 10;
    exp_47_ram[1067] = 55;
    exp_47_ram[1068] = 231;
    exp_47_ram[1069] = 87;
    exp_47_ram[1070] = 231;
    exp_47_ram[1071] = 70;
    exp_47_ram[1072] = 199;
    exp_47_ram[1073] = 71;
    exp_47_ram[1074] = 39;
    exp_47_ram[1075] = 202;
    exp_47_ram[1076] = 247;
    exp_47_ram[1077] = 247;
    exp_47_ram[1078] = 231;
    exp_47_ram[1079] = 198;
    exp_47_ram[1080] = 247;
    exp_47_ram[1081] = 215;
    exp_47_ram[1082] = 1;
    exp_47_ram[1083] = 244;
    exp_47_ram[1084] = 151;
    exp_47_ram[1085] = 228;
    exp_47_ram[1086] = 215;
    exp_47_ram[1087] = 5;
    exp_47_ram[1088] = 245;
    exp_47_ram[1089] = 247;
    exp_47_ram[1090] = 15;
    exp_47_ram[1091] = 164;
    exp_47_ram[1092] = 245;
    exp_47_ram[1093] = 149;
    exp_47_ram[1094] = 244;
    exp_47_ram[1095] = 37;
    exp_47_ram[1096] = 244;
    exp_47_ram[1097] = 52;
    exp_47_ram[1098] = 181;
    exp_47_ram[1099] = 193;
    exp_47_ram[1100] = 133;
    exp_47_ram[1101] = 129;
    exp_47_ram[1102] = 65;
    exp_47_ram[1103] = 1;
    exp_47_ram[1104] = 193;
    exp_47_ram[1105] = 129;
    exp_47_ram[1106] = 65;
    exp_47_ram[1107] = 1;
    exp_47_ram[1108] = 1;
    exp_47_ram[1109] = 0;
    exp_47_ram[1110] = 1;
    exp_47_ram[1111] = 17;
    exp_47_ram[1112] = 129;
    exp_47_ram[1113] = 5;
    exp_47_ram[1114] = 31;
    exp_47_ram[1115] = 0;
    exp_47_ram[1116] = 7;
    exp_47_ram[1117] = 0;
    exp_47_ram[1118] = 95;
    exp_47_ram[1119] = 0;
    exp_47_ram[1120] = 135;
    exp_47_ram[1121] = 245;
    exp_47_ram[1122] = 4;
    exp_47_ram[1123] = 164;
    exp_47_ram[1124] = 4;
    exp_47_ram[1125] = 193;
    exp_47_ram[1126] = 129;
    exp_47_ram[1127] = 0;
    exp_47_ram[1128] = 1;
    exp_47_ram[1129] = 0;
    exp_47_ram[1130] = 1;
    exp_47_ram[1131] = 145;
    exp_47_ram[1132] = 5;
    exp_47_ram[1133] = 0;
    exp_47_ram[1134] = 129;
    exp_47_ram[1135] = 17;
    exp_47_ram[1136] = 5;
    exp_47_ram[1137] = 95;
    exp_47_ram[1138] = 164;
    exp_47_ram[1139] = 164;
    exp_47_ram[1140] = 0;
    exp_47_ram[1141] = 180;
    exp_47_ram[1142] = 148;
    exp_47_ram[1143] = 135;
    exp_47_ram[1144] = 193;
    exp_47_ram[1145] = 135;
    exp_47_ram[1146] = 129;
    exp_47_ram[1147] = 167;
    exp_47_ram[1148] = 65;
    exp_47_ram[1149] = 1;
    exp_47_ram[1150] = 0;
    exp_47_ram[1151] = 1;
    exp_47_ram[1152] = 0;
    exp_47_ram[1153] = 145;
    exp_47_ram[1154] = 96;
    exp_47_ram[1155] = 5;
    exp_47_ram[1156] = 69;
    exp_47_ram[1157] = 1;
    exp_47_ram[1158] = 17;
    exp_47_ram[1159] = 129;
    exp_47_ram[1160] = 33;
    exp_47_ram[1161] = 49;
    exp_47_ram[1162] = 65;
    exp_47_ram[1163] = 95;
    exp_47_ram[1164] = 0;
    exp_47_ram[1165] = 80;
    exp_47_ram[1166] = 197;
    exp_47_ram[1167] = 129;
    exp_47_ram[1168] = 31;
    exp_47_ram[1169] = 132;
    exp_47_ram[1170] = 0;
    exp_47_ram[1171] = 137;
    exp_47_ram[1172] = 23;
    exp_47_ram[1173] = 245;
    exp_47_ram[1174] = 1;
    exp_47_ram[1175] = 0;
    exp_47_ram[1176] = 183;
    exp_47_ram[1177] = 48;
    exp_47_ram[1178] = 137;
    exp_47_ram[1179] = 95;
    exp_47_ram[1180] = 36;
    exp_47_ram[1181] = 4;
    exp_47_ram[1182] = 48;
    exp_47_ram[1183] = 68;
    exp_47_ram[1184] = 23;
    exp_47_ram[1185] = 245;
    exp_47_ram[1186] = 129;
    exp_47_ram[1187] = 183;
    exp_47_ram[1188] = 31;
    exp_47_ram[1189] = 36;
    exp_47_ram[1190] = 196;
    exp_47_ram[1191] = 160;
    exp_47_ram[1192] = 160;
    exp_47_ram[1193] = 0;
    exp_47_ram[1194] = 161;
    exp_47_ram[1195] = 129;
    exp_47_ram[1196] = 177;
    exp_47_ram[1197] = 36;
    exp_47_ram[1198] = 7;
    exp_47_ram[1199] = 244;
    exp_47_ram[1200] = 193;
    exp_47_ram[1201] = 160;
    exp_47_ram[1202] = 7;
    exp_47_ram[1203] = 244;
    exp_47_ram[1204] = 132;
    exp_47_ram[1205] = 0;
    exp_47_ram[1206] = 161;
    exp_47_ram[1207] = 129;
    exp_47_ram[1208] = 177;
    exp_47_ram[1209] = 68;
    exp_47_ram[1210] = 7;
    exp_47_ram[1211] = 244;
    exp_47_ram[1212] = 193;
    exp_47_ram[1213] = 160;
    exp_47_ram[1214] = 7;
    exp_47_ram[1215] = 244;
    exp_47_ram[1216] = 68;
    exp_47_ram[1217] = 0;
    exp_47_ram[1218] = 161;
    exp_47_ram[1219] = 129;
    exp_47_ram[1220] = 177;
    exp_47_ram[1221] = 68;
    exp_47_ram[1222] = 7;
    exp_47_ram[1223] = 244;
    exp_47_ram[1224] = 193;
    exp_47_ram[1225] = 160;
    exp_47_ram[1226] = 7;
    exp_47_ram[1227] = 244;
    exp_47_ram[1228] = 4;
    exp_47_ram[1229] = 0;
    exp_47_ram[1230] = 161;
    exp_47_ram[1231] = 129;
    exp_47_ram[1232] = 177;
    exp_47_ram[1233] = 36;
    exp_47_ram[1234] = 7;
    exp_47_ram[1235] = 244;
    exp_47_ram[1236] = 193;
    exp_47_ram[1237] = 128;
    exp_47_ram[1238] = 7;
    exp_47_ram[1239] = 244;
    exp_47_ram[1240] = 68;
    exp_47_ram[1241] = 197;
    exp_47_ram[1242] = 192;
    exp_47_ram[1243] = 161;
    exp_47_ram[1244] = 177;
    exp_47_ram[1245] = 129;
    exp_47_ram[1246] = 193;
    exp_47_ram[1247] = 64;
    exp_47_ram[1248] = 7;
    exp_47_ram[1249] = 244;
    exp_47_ram[1250] = 192;
    exp_47_ram[1251] = 161;
    exp_47_ram[1252] = 177;
    exp_47_ram[1253] = 129;
    exp_47_ram[1254] = 193;
    exp_47_ram[1255] = 160;
    exp_47_ram[1256] = 7;
    exp_47_ram[1257] = 244;
    exp_47_ram[1258] = 208;
    exp_47_ram[1259] = 161;
    exp_47_ram[1260] = 129;
    exp_47_ram[1261] = 177;
    exp_47_ram[1262] = 193;
    exp_47_ram[1263] = 7;
    exp_47_ram[1264] = 244;
    exp_47_ram[1265] = 193;
    exp_47_ram[1266] = 65;
    exp_47_ram[1267] = 1;
    exp_47_ram[1268] = 7;
    exp_47_ram[1269] = 244;
    exp_47_ram[1270] = 160;
    exp_47_ram[1271] = 244;
    exp_47_ram[1272] = 129;
    exp_47_ram[1273] = 129;
    exp_47_ram[1274] = 137;
    exp_47_ram[1275] = 193;
    exp_47_ram[1276] = 1;
    exp_47_ram[1277] = 0;
    exp_47_ram[1278] = 1;
    exp_47_ram[1279] = 65;
    exp_47_ram[1280] = 1;
    exp_47_ram[1281] = 129;
    exp_47_ram[1282] = 145;
    exp_47_ram[1283] = 33;
    exp_47_ram[1284] = 49;
    exp_47_ram[1285] = 81;
    exp_47_ram[1286] = 17;
    exp_47_ram[1287] = 97;
    exp_47_ram[1288] = 113;
    exp_47_ram[1289] = 129;
    exp_47_ram[1290] = 145;
    exp_47_ram[1291] = 5;
    exp_47_ram[1292] = 5;
    exp_47_ram[1293] = 6;
    exp_47_ram[1294] = 32;
    exp_47_ram[1295] = 64;
    exp_47_ram[1296] = 10;
    exp_47_ram[1297] = 9;
    exp_47_ram[1298] = 31;
    exp_47_ram[1299] = 160;
    exp_47_ram[1300] = 10;
    exp_47_ram[1301] = 213;
    exp_47_ram[1302] = 15;
    exp_47_ram[1303] = 25;
    exp_47_ram[1304] = 9;
    exp_47_ram[1305] = 164;
    exp_47_ram[1306] = 170;
    exp_47_ram[1307] = 164;
    exp_47_ram[1308] = 164;
    exp_47_ram[1309] = 233;
    exp_47_ram[1310] = 5;
    exp_47_ram[1311] = 7;
    exp_47_ram[1312] = 95;
    exp_47_ram[1313] = 1;
    exp_47_ram[1314] = 0;
    exp_47_ram[1315] = 0;
    exp_47_ram[1316] = 12;
    exp_47_ram[1317] = 12;
    exp_47_ram[1318] = 9;
    exp_47_ram[1319] = 95;
    exp_47_ram[1320] = 12;
    exp_47_ram[1321] = 12;
    exp_47_ram[1322] = 5;
    exp_47_ram[1323] = 28;
    exp_47_ram[1324] = 143;
    exp_47_ram[1325] = 9;
    exp_47_ram[1326] = 164;
    exp_47_ram[1327] = 164;
    exp_47_ram[1328] = 164;
    exp_47_ram[1329] = 122;
    exp_47_ram[1330] = 122;
    exp_47_ram[1331] = 5;
    exp_47_ram[1332] = 249;
    exp_47_ram[1333] = 31;
    exp_47_ram[1334] = 1;
    exp_47_ram[1335] = 4;
    exp_47_ram[1336] = 5;
    exp_47_ram[1337] = 16;
    exp_47_ram[1338] = 177;
    exp_47_ram[1339] = 5;
    exp_47_ram[1340] = 161;
    exp_47_ram[1341] = 170;
    exp_47_ram[1342] = 193;
    exp_47_ram[1343] = 0;
    exp_47_ram[1344] = 5;
    exp_47_ram[1345] = 16;
    exp_47_ram[1346] = 177;
    exp_47_ram[1347] = 5;
    exp_47_ram[1348] = 161;
    exp_47_ram[1349] = 193;
    exp_47_ram[1350] = 192;
    exp_47_ram[1351] = 73;
    exp_47_ram[1352] = 80;
    exp_47_ram[1353] = 20;
    exp_47_ram[1354] = 161;
    exp_47_ram[1355] = 177;
    exp_47_ram[1356] = 180;
    exp_47_ram[1357] = 164;
    exp_47_ram[1358] = 36;
    exp_47_ram[1359] = 100;
    exp_47_ram[1360] = 52;
    exp_47_ram[1361] = 154;
    exp_47_ram[1362] = 244;
    exp_47_ram[1363] = 112;
    exp_47_ram[1364] = 15;
    exp_47_ram[1365] = 164;
    exp_47_ram[1366] = 68;
    exp_47_ram[1367] = 193;
    exp_47_ram[1368] = 4;
    exp_47_ram[1369] = 129;
    exp_47_ram[1370] = 65;
    exp_47_ram[1371] = 1;
    exp_47_ram[1372] = 193;
    exp_47_ram[1373] = 129;
    exp_47_ram[1374] = 65;
    exp_47_ram[1375] = 1;
    exp_47_ram[1376] = 193;
    exp_47_ram[1377] = 129;
    exp_47_ram[1378] = 65;
    exp_47_ram[1379] = 1;
    exp_47_ram[1380] = 0;
    exp_47_ram[1381] = 1;
    exp_47_ram[1382] = 97;
    exp_47_ram[1383] = 69;
    exp_47_ram[1384] = 64;
    exp_47_ram[1385] = 145;
    exp_47_ram[1386] = 33;
    exp_47_ram[1387] = 240;
    exp_47_ram[1388] = 65;
    exp_47_ram[1389] = 81;
    exp_47_ram[1390] = 16;
    exp_47_ram[1391] = 5;
    exp_47_ram[1392] = 144;
    exp_47_ram[1393] = 129;
    exp_47_ram[1394] = 1;
    exp_47_ram[1395] = 17;
    exp_47_ram[1396] = 129;
    exp_47_ram[1397] = 49;
    exp_47_ram[1398] = 65;
    exp_47_ram[1399] = 145;
    exp_47_ram[1400] = 97;
    exp_47_ram[1401] = 81;
    exp_47_ram[1402] = 1;
    exp_47_ram[1403] = 1;
    exp_47_ram[1404] = 1;
    exp_47_ram[1405] = 223;
    exp_47_ram[1406] = 1;
    exp_47_ram[1407] = 223;
    exp_47_ram[1408] = 5;
    exp_47_ram[1409] = 5;
    exp_47_ram[1410] = 129;
    exp_47_ram[1411] = 223;
    exp_47_ram[1412] = 1;
    exp_47_ram[1413] = 65;
    exp_47_ram[1414] = 64;
    exp_47_ram[1415] = 129;
    exp_47_ram[1416] = 231;
    exp_47_ram[1417] = 1;
    exp_47_ram[1418] = 241;
    exp_47_ram[1419] = 95;
    exp_47_ram[1420] = 1;
    exp_47_ram[1421] = 95;
    exp_47_ram[1422] = 64;
    exp_47_ram[1423] = 5;
    exp_47_ram[1424] = 5;
    exp_47_ram[1425] = 1;
    exp_47_ram[1426] = 193;
    exp_47_ram[1427] = 65;
    exp_47_ram[1428] = 145;
    exp_47_ram[1429] = 97;
    exp_47_ram[1430] = 81;
    exp_47_ram[1431] = 1;
    exp_47_ram[1432] = 1;
    exp_47_ram[1433] = 207;
    exp_47_ram[1434] = 1;
    exp_47_ram[1435] = 223;
    exp_47_ram[1436] = 5;
    exp_47_ram[1437] = 5;
    exp_47_ram[1438] = 129;
    exp_47_ram[1439] = 223;
    exp_47_ram[1440] = 64;
    exp_47_ram[1441] = 193;
    exp_47_ram[1442] = 1;
    exp_47_ram[1443] = 145;
    exp_47_ram[1444] = 15;
    exp_47_ram[1445] = 1;
    exp_47_ram[1446] = 31;
    exp_47_ram[1447] = 64;
    exp_47_ram[1448] = 5;
    exp_47_ram[1449] = 5;
    exp_47_ram[1450] = 1;
    exp_47_ram[1451] = 9;
    exp_47_ram[1452] = 15;
    exp_47_ram[1453] = 1;
    exp_47_ram[1454] = 31;
    exp_47_ram[1455] = 5;
    exp_47_ram[1456] = 5;
    exp_47_ram[1457] = 180;
    exp_47_ram[1458] = 149;
    exp_47_ram[1459] = 170;
    exp_47_ram[1460] = 16;
    exp_47_ram[1461] = 135;
    exp_47_ram[1462] = 244;
    exp_47_ram[1463] = 55;
    exp_47_ram[1464] = 0;
    exp_47_ram[1465] = 193;
    exp_47_ram[1466] = 129;
    exp_47_ram[1467] = 65;
    exp_47_ram[1468] = 1;
    exp_47_ram[1469] = 193;
    exp_47_ram[1470] = 129;
    exp_47_ram[1471] = 65;
    exp_47_ram[1472] = 1;
    exp_47_ram[1473] = 1;
    exp_47_ram[1474] = 0;
    exp_47_ram[1475] = 1;
    exp_47_ram[1476] = 5;
    exp_47_ram[1477] = 33;
    exp_47_ram[1478] = 64;
    exp_47_ram[1479] = 5;
    exp_47_ram[1480] = 193;
    exp_47_ram[1481] = 17;
    exp_47_ram[1482] = 129;
    exp_47_ram[1483] = 145;
    exp_47_ram[1484] = 49;
    exp_47_ram[1485] = 207;
    exp_47_ram[1486] = 64;
    exp_47_ram[1487] = 193;
    exp_47_ram[1488] = 1;
    exp_47_ram[1489] = 9;
    exp_47_ram[1490] = 143;
    exp_47_ram[1491] = 1;
    exp_47_ram[1492] = 159;
    exp_47_ram[1493] = 5;
    exp_47_ram[1494] = 5;
    exp_47_ram[1495] = 48;
    exp_47_ram[1496] = 0;
    exp_47_ram[1497] = 7;
    exp_47_ram[1498] = 245;
    exp_47_ram[1499] = 167;
    exp_47_ram[1500] = 7;
    exp_47_ram[1501] = 183;
    exp_47_ram[1502] = 4;
    exp_47_ram[1503] = 4;
    exp_47_ram[1504] = 1;
    exp_47_ram[1505] = 95;
    exp_47_ram[1506] = 64;
    exp_47_ram[1507] = 1;
    exp_47_ram[1508] = 9;
    exp_47_ram[1509] = 207;
    exp_47_ram[1510] = 48;
    exp_47_ram[1511] = 16;
    exp_47_ram[1512] = 249;
    exp_47_ram[1513] = 193;
    exp_47_ram[1514] = 4;
    exp_47_ram[1515] = 129;
    exp_47_ram[1516] = 1;
    exp_47_ram[1517] = 193;
    exp_47_ram[1518] = 4;
    exp_47_ram[1519] = 65;
    exp_47_ram[1520] = 1;
    exp_47_ram[1521] = 0;
    exp_47_ram[1522] = 9;
    exp_47_ram[1523] = 193;
    exp_47_ram[1524] = 64;
    exp_47_ram[1525] = 1;
    exp_47_ram[1526] = 143;
    exp_47_ram[1527] = 1;
    exp_47_ram[1528] = 95;
    exp_47_ram[1529] = 245;
    exp_47_ram[1530] = 164;
    exp_47_ram[1531] = 133;
    exp_47_ram[1532] = 180;
    exp_47_ram[1533] = 151;
    exp_47_ram[1534] = 149;
    exp_47_ram[1535] = 5;
    exp_47_ram[1536] = 7;
    exp_47_ram[1537] = 0;
    exp_47_ram[1538] = 4;
    exp_47_ram[1539] = 0;
    exp_47_ram[1540] = 159;
    exp_47_ram[1541] = 9;
    exp_47_ram[1542] = 64;
    exp_47_ram[1543] = 193;
    exp_47_ram[1544] = 1;
    exp_47_ram[1545] = 207;
    exp_47_ram[1546] = 1;
    exp_47_ram[1547] = 159;
    exp_47_ram[1548] = 5;
    exp_47_ram[1549] = 0;
    exp_47_ram[1550] = 5;
    exp_47_ram[1551] = 169;
    exp_47_ram[1552] = 95;
    exp_47_ram[1553] = 9;
    exp_47_ram[1554] = 223;
    exp_47_ram[1555] = 1;
    exp_47_ram[1556] = 5;
    exp_47_ram[1557] = 5;
    exp_47_ram[1558] = 193;
    exp_47_ram[1559] = 17;
    exp_47_ram[1560] = 159;
    exp_47_ram[1561] = 193;
    exp_47_ram[1562] = 64;
    exp_47_ram[1563] = 1;
    exp_47_ram[1564] = 15;
    exp_47_ram[1565] = 1;
    exp_47_ram[1566] = 223;
    exp_47_ram[1567] = 193;
    exp_47_ram[1568] = 1;
    exp_47_ram[1569] = 0;
    exp_47_ram[1570] = 1;
    exp_47_ram[1571] = 145;
    exp_47_ram[1572] = 33;
    exp_47_ram[1573] = 69;
    exp_47_ram[1574] = 5;
    exp_47_ram[1575] = 17;
    exp_47_ram[1576] = 4;
    exp_47_ram[1577] = 9;
    exp_47_ram[1578] = 129;
    exp_47_ram[1579] = 49;
    exp_47_ram[1580] = 223;
    exp_47_ram[1581] = 0;
    exp_47_ram[1582] = 5;
    exp_47_ram[1583] = 0;
    exp_47_ram[1584] = 6;
    exp_47_ram[1585] = 38;
    exp_47_ram[1586] = 197;
    exp_47_ram[1587] = 150;
    exp_47_ram[1588] = 1;
    exp_47_ram[1589] = 95;
    exp_47_ram[1590] = 0;
    exp_47_ram[1591] = 1;
    exp_47_ram[1592] = 64;
    exp_47_ram[1593] = 68;
    exp_47_ram[1594] = 143;
    exp_47_ram[1595] = 9;
    exp_47_ram[1596] = 4;
    exp_47_ram[1597] = 159;
    exp_47_ram[1598] = 68;
    exp_47_ram[1599] = 169;
    exp_47_ram[1600] = 193;
    exp_47_ram[1601] = 68;
    exp_47_ram[1602] = 129;
    exp_47_ram[1603] = 65;
    exp_47_ram[1604] = 1;
    exp_47_ram[1605] = 193;
    exp_47_ram[1606] = 1;
    exp_47_ram[1607] = 0;
    exp_47_ram[1608] = 1;
    exp_47_ram[1609] = 17;
    exp_47_ram[1610] = 129;
    exp_47_ram[1611] = 33;
    exp_47_ram[1612] = 49;
    exp_47_ram[1613] = 1;
    exp_47_ram[1614] = 164;
    exp_47_ram[1615] = 207;
    exp_47_ram[1616] = 164;
    exp_47_ram[1617] = 180;
    exp_47_ram[1618] = 0;
    exp_47_ram[1619] = 207;
    exp_47_ram[1620] = 5;
    exp_47_ram[1621] = 5;
    exp_47_ram[1622] = 132;
    exp_47_ram[1623] = 196;
    exp_47_ram[1624] = 166;
    exp_47_ram[1625] = 7;
    exp_47_ram[1626] = 6;
    exp_47_ram[1627] = 182;
    exp_47_ram[1628] = 7;
    exp_47_ram[1629] = 6;
    exp_47_ram[1630] = 196;
    exp_47_ram[1631] = 6;
    exp_47_ram[1632] = 0;
    exp_47_ram[1633] = 9;
    exp_47_ram[1634] = 7;
    exp_47_ram[1635] = 198;
    exp_47_ram[1636] = 9;
    exp_47_ram[1637] = 7;
    exp_47_ram[1638] = 214;
    exp_47_ram[1639] = 9;
    exp_47_ram[1640] = 7;
    exp_47_ram[1641] = 215;
    exp_47_ram[1642] = 0;
    exp_47_ram[1643] = 7;
    exp_47_ram[1644] = 193;
    exp_47_ram[1645] = 129;
    exp_47_ram[1646] = 65;
    exp_47_ram[1647] = 1;
    exp_47_ram[1648] = 1;
    exp_47_ram[1649] = 0;
    exp_47_ram[1650] = 1;
    exp_47_ram[1651] = 17;
    exp_47_ram[1652] = 129;
    exp_47_ram[1653] = 1;
    exp_47_ram[1654] = 0;
    exp_47_ram[1655] = 31;
    exp_47_ram[1656] = 0;
    exp_47_ram[1657] = 193;
    exp_47_ram[1658] = 129;
    exp_47_ram[1659] = 1;
    exp_47_ram[1660] = 0;
    exp_47_ram[1661] = 1;
    exp_47_ram[1662] = 17;
    exp_47_ram[1663] = 129;
    exp_47_ram[1664] = 1;
    exp_47_ram[1665] = 0;
    exp_47_ram[1666] = 95;
    exp_47_ram[1667] = 16;
    exp_47_ram[1668] = 244;
    exp_47_ram[1669] = 4;
    exp_47_ram[1670] = 192;
    exp_47_ram[1671] = 132;
    exp_47_ram[1672] = 0;
    exp_47_ram[1673] = 15;
    exp_47_ram[1674] = 192;
    exp_47_ram[1675] = 196;
    exp_47_ram[1676] = 23;
    exp_47_ram[1677] = 244;
    exp_47_ram[1678] = 0;
    exp_47_ram[1679] = 199;
    exp_47_ram[1680] = 7;
    exp_47_ram[1681] = 196;
    exp_47_ram[1682] = 159;
    exp_47_ram[1683] = 0;
    exp_47_ram[1684] = 7;
    exp_47_ram[1685] = 160;
    exp_47_ram[1686] = 247;
    exp_47_ram[1687] = 7;
    exp_47_ram[1688] = 31;
    exp_47_ram[1689] = 196;
    exp_47_ram[1690] = 240;
    exp_47_ram[1691] = 231;
    exp_47_ram[1692] = 192;
    exp_47_ram[1693] = 196;
    exp_47_ram[1694] = 23;
    exp_47_ram[1695] = 244;
    exp_47_ram[1696] = 0;
    exp_47_ram[1697] = 199;
    exp_47_ram[1698] = 7;
    exp_47_ram[1699] = 196;
    exp_47_ram[1700] = 31;
    exp_47_ram[1701] = 0;
    exp_47_ram[1702] = 7;
    exp_47_ram[1703] = 160;
    exp_47_ram[1704] = 247;
    exp_47_ram[1705] = 7;
    exp_47_ram[1706] = 159;
    exp_47_ram[1707] = 196;
    exp_47_ram[1708] = 16;
    exp_47_ram[1709] = 231;
    exp_47_ram[1710] = 132;
    exp_47_ram[1711] = 23;
    exp_47_ram[1712] = 244;
    exp_47_ram[1713] = 132;
    exp_47_ram[1714] = 144;
    exp_47_ram[1715] = 231;
    exp_47_ram[1716] = 0;
    exp_47_ram[1717] = 199;
    exp_47_ram[1718] = 7;
    exp_47_ram[1719] = 0;
    exp_47_ram[1720] = 31;
    exp_47_ram[1721] = 0;
    exp_47_ram[1722] = 193;
    exp_47_ram[1723] = 129;
    exp_47_ram[1724] = 1;
    exp_47_ram[1725] = 0;
    exp_47_ram[1726] = 1;
    exp_47_ram[1727] = 17;
    exp_47_ram[1728] = 129;
    exp_47_ram[1729] = 1;
    exp_47_ram[1730] = 196;
    exp_47_ram[1731] = 80;
    exp_47_ram[1732] = 231;
    exp_47_ram[1733] = 196;
    exp_47_ram[1734] = 144;
    exp_47_ram[1735] = 231;
    exp_47_ram[1736] = 196;
    exp_47_ram[1737] = 144;
    exp_47_ram[1738] = 231;
    exp_47_ram[1739] = 196;
    exp_47_ram[1740] = 16;
    exp_47_ram[1741] = 231;
    exp_47_ram[1742] = 196;
    exp_47_ram[1743] = 80;
    exp_47_ram[1744] = 231;
    exp_47_ram[1745] = 196;
    exp_47_ram[1746] = 7;
    exp_47_ram[1747] = 196;
    exp_47_ram[1748] = 240;
    exp_47_ram[1749] = 231;
    exp_47_ram[1750] = 196;
    exp_47_ram[1751] = 31;
    exp_47_ram[1752] = 5;
    exp_47_ram[1753] = 5;
    exp_47_ram[1754] = 7;
    exp_47_ram[1755] = 7;
    exp_47_ram[1756] = 143;
    exp_47_ram[1757] = 0;
    exp_47_ram[1758] = 15;
    exp_47_ram[1759] = 5;
    exp_47_ram[1760] = 5;
    exp_47_ram[1761] = 228;
    exp_47_ram[1762] = 244;
    exp_47_ram[1763] = 4;
    exp_47_ram[1764] = 7;
    exp_47_ram[1765] = 95;
    exp_47_ram[1766] = 164;
    exp_47_ram[1767] = 196;
    exp_47_ram[1768] = 207;
    exp_47_ram[1769] = 5;
    exp_47_ram[1770] = 7;
    exp_47_ram[1771] = 31;
    exp_47_ram[1772] = 0;
    exp_47_ram[1773] = 7;
    exp_47_ram[1774] = 7;
    exp_47_ram[1775] = 95;
    exp_47_ram[1776] = 95;
    exp_47_ram[1777] = 1;
    exp_47_ram[1778] = 17;
    exp_47_ram[1779] = 129;
    exp_47_ram[1780] = 33;
    exp_47_ram[1781] = 49;
    exp_47_ram[1782] = 65;
    exp_47_ram[1783] = 81;
    exp_47_ram[1784] = 97;
    exp_47_ram[1785] = 113;
    exp_47_ram[1786] = 129;
    exp_47_ram[1787] = 145;
    exp_47_ram[1788] = 161;
    exp_47_ram[1789] = 177;
    exp_47_ram[1790] = 1;
    exp_47_ram[1791] = 16;
    exp_47_ram[1792] = 244;
    exp_47_ram[1793] = 16;
    exp_47_ram[1794] = 0;
    exp_47_ram[1795] = 228;
    exp_47_ram[1796] = 244;
    exp_47_ram[1797] = 79;
    exp_47_ram[1798] = 164;
    exp_47_ram[1799] = 180;
    exp_47_ram[1800] = 4;
    exp_47_ram[1801] = 0;
    exp_47_ram[1802] = 196;
    exp_47_ram[1803] = 52;
    exp_47_ram[1804] = 135;
    exp_47_ram[1805] = 247;
    exp_47_ram[1806] = 244;
    exp_47_ram[1807] = 196;
    exp_47_ram[1808] = 52;
    exp_47_ram[1809] = 135;
    exp_47_ram[1810] = 247;
    exp_47_ram[1811] = 244;
    exp_47_ram[1812] = 196;
    exp_47_ram[1813] = 52;
    exp_47_ram[1814] = 135;
    exp_47_ram[1815] = 247;
    exp_47_ram[1816] = 244;
    exp_47_ram[1817] = 196;
    exp_47_ram[1818] = 52;
    exp_47_ram[1819] = 135;
    exp_47_ram[1820] = 247;
    exp_47_ram[1821] = 244;
    exp_47_ram[1822] = 196;
    exp_47_ram[1823] = 71;
    exp_47_ram[1824] = 244;
    exp_47_ram[1825] = 79;
    exp_47_ram[1826] = 5;
    exp_47_ram[1827] = 5;
    exp_47_ram[1828] = 4;
    exp_47_ram[1829] = 68;
    exp_47_ram[1830] = 166;
    exp_47_ram[1831] = 7;
    exp_47_ram[1832] = 6;
    exp_47_ram[1833] = 182;
    exp_47_ram[1834] = 7;
    exp_47_ram[1835] = 6;
    exp_47_ram[1836] = 0;
    exp_47_ram[1837] = 6;
    exp_47_ram[1838] = 212;
    exp_47_ram[1839] = 4;
    exp_47_ram[1840] = 132;
    exp_47_ram[1841] = 196;
    exp_47_ram[1842] = 5;
    exp_47_ram[1843] = 7;
    exp_47_ram[1844] = 198;
    exp_47_ram[1845] = 5;
    exp_47_ram[1846] = 7;
    exp_47_ram[1847] = 214;
    exp_47_ram[1848] = 5;
    exp_47_ram[1849] = 7;
    exp_47_ram[1850] = 215;
    exp_47_ram[1851] = 196;
    exp_47_ram[1852] = 64;
    exp_47_ram[1853] = 31;
    exp_47_ram[1854] = 15;
    exp_47_ram[1855] = 164;
    exp_47_ram[1856] = 180;
    exp_47_ram[1857] = 4;
    exp_47_ram[1858] = 0;
    exp_47_ram[1859] = 4;
    exp_47_ram[1860] = 68;
    exp_47_ram[1861] = 52;
    exp_47_ram[1862] = 134;
    exp_47_ram[1863] = 215;
    exp_47_ram[1864] = 0;
    exp_47_ram[1865] = 215;
    exp_47_ram[1866] = 214;
    exp_47_ram[1867] = 52;
    exp_47_ram[1868] = 134;
    exp_47_ram[1869] = 215;
    exp_47_ram[1870] = 215;
    exp_47_ram[1871] = 5;
    exp_47_ram[1872] = 54;
    exp_47_ram[1873] = 7;
    exp_47_ram[1874] = 36;
    exp_47_ram[1875] = 52;
    exp_47_ram[1876] = 4;
    exp_47_ram[1877] = 68;
    exp_47_ram[1878] = 52;
    exp_47_ram[1879] = 134;
    exp_47_ram[1880] = 215;
    exp_47_ram[1881] = 0;
    exp_47_ram[1882] = 215;
    exp_47_ram[1883] = 214;
    exp_47_ram[1884] = 52;
    exp_47_ram[1885] = 134;
    exp_47_ram[1886] = 215;
    exp_47_ram[1887] = 215;
    exp_47_ram[1888] = 5;
    exp_47_ram[1889] = 86;
    exp_47_ram[1890] = 7;
    exp_47_ram[1891] = 68;
    exp_47_ram[1892] = 84;
    exp_47_ram[1893] = 4;
    exp_47_ram[1894] = 68;
    exp_47_ram[1895] = 52;
    exp_47_ram[1896] = 134;
    exp_47_ram[1897] = 215;
    exp_47_ram[1898] = 0;
    exp_47_ram[1899] = 215;
    exp_47_ram[1900] = 214;
    exp_47_ram[1901] = 52;
    exp_47_ram[1902] = 134;
    exp_47_ram[1903] = 215;
    exp_47_ram[1904] = 215;
    exp_47_ram[1905] = 5;
    exp_47_ram[1906] = 118;
    exp_47_ram[1907] = 7;
    exp_47_ram[1908] = 100;
    exp_47_ram[1909] = 116;
    exp_47_ram[1910] = 4;
    exp_47_ram[1911] = 68;
    exp_47_ram[1912] = 52;
    exp_47_ram[1913] = 134;
    exp_47_ram[1914] = 215;
    exp_47_ram[1915] = 0;
    exp_47_ram[1916] = 215;
    exp_47_ram[1917] = 214;
    exp_47_ram[1918] = 52;
    exp_47_ram[1919] = 134;
    exp_47_ram[1920] = 215;
    exp_47_ram[1921] = 215;
    exp_47_ram[1922] = 5;
    exp_47_ram[1923] = 150;
    exp_47_ram[1924] = 7;
    exp_47_ram[1925] = 132;
    exp_47_ram[1926] = 148;
    exp_47_ram[1927] = 196;
    exp_47_ram[1928] = 71;
    exp_47_ram[1929] = 244;
    exp_47_ram[1930] = 15;
    exp_47_ram[1931] = 5;
    exp_47_ram[1932] = 5;
    exp_47_ram[1933] = 4;
    exp_47_ram[1934] = 68;
    exp_47_ram[1935] = 166;
    exp_47_ram[1936] = 7;
    exp_47_ram[1937] = 6;
    exp_47_ram[1938] = 182;
    exp_47_ram[1939] = 7;
    exp_47_ram[1940] = 6;
    exp_47_ram[1941] = 0;
    exp_47_ram[1942] = 6;
    exp_47_ram[1943] = 212;
    exp_47_ram[1944] = 4;
    exp_47_ram[1945] = 4;
    exp_47_ram[1946] = 68;
    exp_47_ram[1947] = 5;
    exp_47_ram[1948] = 7;
    exp_47_ram[1949] = 198;
    exp_47_ram[1950] = 5;
    exp_47_ram[1951] = 7;
    exp_47_ram[1952] = 214;
    exp_47_ram[1953] = 5;
    exp_47_ram[1954] = 7;
    exp_47_ram[1955] = 215;
    exp_47_ram[1956] = 196;
    exp_47_ram[1957] = 0;
    exp_47_ram[1958] = 223;
    exp_47_ram[1959] = 207;
    exp_47_ram[1960] = 164;
    exp_47_ram[1961] = 180;
    exp_47_ram[1962] = 4;
    exp_47_ram[1963] = 0;
    exp_47_ram[1964] = 196;
    exp_47_ram[1965] = 52;
    exp_47_ram[1966] = 135;
    exp_47_ram[1967] = 247;
    exp_47_ram[1968] = 244;
    exp_47_ram[1969] = 196;
    exp_47_ram[1970] = 52;
    exp_47_ram[1971] = 135;
    exp_47_ram[1972] = 247;
    exp_47_ram[1973] = 244;
    exp_47_ram[1974] = 196;
    exp_47_ram[1975] = 52;
    exp_47_ram[1976] = 135;
    exp_47_ram[1977] = 247;
    exp_47_ram[1978] = 244;
    exp_47_ram[1979] = 196;
    exp_47_ram[1980] = 52;
    exp_47_ram[1981] = 135;
    exp_47_ram[1982] = 247;
    exp_47_ram[1983] = 244;
    exp_47_ram[1984] = 196;
    exp_47_ram[1985] = 71;
    exp_47_ram[1986] = 244;
    exp_47_ram[1987] = 207;
    exp_47_ram[1988] = 5;
    exp_47_ram[1989] = 5;
    exp_47_ram[1990] = 4;
    exp_47_ram[1991] = 68;
    exp_47_ram[1992] = 166;
    exp_47_ram[1993] = 7;
    exp_47_ram[1994] = 6;
    exp_47_ram[1995] = 182;
    exp_47_ram[1996] = 7;
    exp_47_ram[1997] = 6;
    exp_47_ram[1998] = 0;
    exp_47_ram[1999] = 6;
    exp_47_ram[2000] = 212;
    exp_47_ram[2001] = 4;
    exp_47_ram[2002] = 132;
    exp_47_ram[2003] = 196;
    exp_47_ram[2004] = 5;
    exp_47_ram[2005] = 7;
    exp_47_ram[2006] = 198;
    exp_47_ram[2007] = 5;
    exp_47_ram[2008] = 7;
    exp_47_ram[2009] = 214;
    exp_47_ram[2010] = 5;
    exp_47_ram[2011] = 7;
    exp_47_ram[2012] = 215;
    exp_47_ram[2013] = 196;
    exp_47_ram[2014] = 192;
    exp_47_ram[2015] = 159;
    exp_47_ram[2016] = 143;
    exp_47_ram[2017] = 164;
    exp_47_ram[2018] = 180;
    exp_47_ram[2019] = 4;
    exp_47_ram[2020] = 0;
    exp_47_ram[2021] = 4;
    exp_47_ram[2022] = 68;
    exp_47_ram[2023] = 52;
    exp_47_ram[2024] = 134;
    exp_47_ram[2025] = 0;
    exp_47_ram[2026] = 7;
    exp_47_ram[2027] = 7;
    exp_47_ram[2028] = 207;
    exp_47_ram[2029] = 5;
    exp_47_ram[2030] = 5;
    exp_47_ram[2031] = 228;
    exp_47_ram[2032] = 244;
    exp_47_ram[2033] = 4;
    exp_47_ram[2034] = 68;
    exp_47_ram[2035] = 52;
    exp_47_ram[2036] = 134;
    exp_47_ram[2037] = 0;
    exp_47_ram[2038] = 7;
    exp_47_ram[2039] = 7;
    exp_47_ram[2040] = 207;
    exp_47_ram[2041] = 5;
    exp_47_ram[2042] = 5;
    exp_47_ram[2043] = 228;
    exp_47_ram[2044] = 244;
    exp_47_ram[2045] = 4;
    exp_47_ram[2046] = 68;
    exp_47_ram[2047] = 52;
    exp_47_ram[2048] = 134;
    exp_47_ram[2049] = 0;
    exp_47_ram[2050] = 7;
    exp_47_ram[2051] = 7;
    exp_47_ram[2052] = 207;
    exp_47_ram[2053] = 5;
    exp_47_ram[2054] = 5;
    exp_47_ram[2055] = 228;
    exp_47_ram[2056] = 244;
    exp_47_ram[2057] = 4;
    exp_47_ram[2058] = 68;
    exp_47_ram[2059] = 52;
    exp_47_ram[2060] = 134;
    exp_47_ram[2061] = 0;
    exp_47_ram[2062] = 7;
    exp_47_ram[2063] = 7;
    exp_47_ram[2064] = 207;
    exp_47_ram[2065] = 5;
    exp_47_ram[2066] = 5;
    exp_47_ram[2067] = 228;
    exp_47_ram[2068] = 244;
    exp_47_ram[2069] = 196;
    exp_47_ram[2070] = 71;
    exp_47_ram[2071] = 244;
    exp_47_ram[2072] = 159;
    exp_47_ram[2073] = 5;
    exp_47_ram[2074] = 5;
    exp_47_ram[2075] = 4;
    exp_47_ram[2076] = 68;
    exp_47_ram[2077] = 166;
    exp_47_ram[2078] = 7;
    exp_47_ram[2079] = 6;
    exp_47_ram[2080] = 182;
    exp_47_ram[2081] = 7;
    exp_47_ram[2082] = 6;
    exp_47_ram[2083] = 0;
    exp_47_ram[2084] = 6;
    exp_47_ram[2085] = 6;
    exp_47_ram[2086] = 0;
    exp_47_ram[2087] = 13;
    exp_47_ram[2088] = 7;
    exp_47_ram[2089] = 198;
    exp_47_ram[2090] = 13;
    exp_47_ram[2091] = 7;
    exp_47_ram[2092] = 214;
    exp_47_ram[2093] = 13;
    exp_47_ram[2094] = 7;
    exp_47_ram[2095] = 215;
    exp_47_ram[2096] = 196;
    exp_47_ram[2097] = 64;
    exp_47_ram[2098] = 223;
    exp_47_ram[2099] = 0;
    exp_47_ram[2100] = 193;
    exp_47_ram[2101] = 129;
    exp_47_ram[2102] = 65;
    exp_47_ram[2103] = 1;
    exp_47_ram[2104] = 193;
    exp_47_ram[2105] = 129;
    exp_47_ram[2106] = 65;
    exp_47_ram[2107] = 1;
    exp_47_ram[2108] = 193;
    exp_47_ram[2109] = 129;
    exp_47_ram[2110] = 65;
    exp_47_ram[2111] = 1;
    exp_47_ram[2112] = 1;
    exp_47_ram[2113] = 0;
    exp_47_ram[2114] = 1;
    exp_47_ram[2115] = 17;
    exp_47_ram[2116] = 129;
    exp_47_ram[2117] = 1;
    exp_47_ram[2118] = 4;
    exp_47_ram[2119] = 128;
    exp_47_ram[2120] = 196;
    exp_47_ram[2121] = 247;
    exp_47_ram[2122] = 196;
    exp_47_ram[2123] = 4;
    exp_47_ram[2124] = 246;
    exp_47_ram[2125] = 231;
    exp_47_ram[2126] = 196;
    exp_47_ram[2127] = 23;
    exp_47_ram[2128] = 244;
    exp_47_ram[2129] = 196;
    exp_47_ram[2130] = 48;
    exp_47_ram[2131] = 231;
    exp_47_ram[2132] = 4;
    exp_47_ram[2133] = 128;
    exp_47_ram[2134] = 132;
    exp_47_ram[2135] = 192;
    exp_47_ram[2136] = 95;
    exp_47_ram[2137] = 132;
    exp_47_ram[2138] = 196;
    exp_47_ram[2139] = 247;
    exp_47_ram[2140] = 64;
    exp_47_ram[2141] = 132;
    exp_47_ram[2142] = 247;
    exp_47_ram[2143] = 7;
    exp_47_ram[2144] = 4;
    exp_47_ram[2145] = 7;
    exp_47_ram[2146] = 7;
    exp_47_ram[2147] = 6;
    exp_47_ram[2148] = 31;
    exp_47_ram[2149] = 132;
    exp_47_ram[2150] = 244;
    exp_47_ram[2151] = 0;
    exp_47_ram[2152] = 68;
    exp_47_ram[2153] = 4;
    exp_47_ram[2154] = 247;
    exp_47_ram[2155] = 7;
    exp_47_ram[2156] = 7;
    exp_47_ram[2157] = 68;
    exp_47_ram[2158] = 4;
    exp_47_ram[2159] = 246;
    exp_47_ram[2160] = 199;
    exp_47_ram[2161] = 7;
    exp_47_ram[2162] = 132;
    exp_47_ram[2163] = 246;
    exp_47_ram[2164] = 247;
    exp_47_ram[2165] = 192;
    exp_47_ram[2166] = 79;
    exp_47_ram[2167] = 128;
    exp_47_ram[2168] = 68;
    exp_47_ram[2169] = 23;
    exp_47_ram[2170] = 244;
    exp_47_ram[2171] = 68;
    exp_47_ram[2172] = 48;
    exp_47_ram[2173] = 231;
    exp_47_ram[2174] = 64;
    exp_47_ram[2175] = 15;
    exp_47_ram[2176] = 132;
    exp_47_ram[2177] = 23;
    exp_47_ram[2178] = 244;
    exp_47_ram[2179] = 132;
    exp_47_ram[2180] = 48;
    exp_47_ram[2181] = 231;
    exp_47_ram[2182] = 0;
    exp_47_ram[2183] = 95;
    exp_47_ram[2184] = 5;
    exp_47_ram[2185] = 244;
    exp_47_ram[2186] = 0;
    exp_47_ram[2187] = 95;
    exp_47_ram[2188] = 5;
    exp_47_ram[2189] = 244;
    exp_47_ram[2190] = 0;
    exp_47_ram[2191] = 95;
    exp_47_ram[2192] = 5;
    exp_47_ram[2193] = 244;
    exp_47_ram[2194] = 4;
    exp_47_ram[2195] = 64;
    exp_47_ram[2196] = 4;
    exp_47_ram[2197] = 95;
    exp_47_ram[2198] = 0;
    exp_47_ram[2199] = 95;
    exp_47_ram[2200] = 5;
    exp_47_ram[2201] = 244;
    exp_47_ram[2202] = 196;
    exp_47_ram[2203] = 223;
    exp_47_ram[2204] = 0;
    exp_47_ram[2205] = 223;
    exp_47_ram[2206] = 5;
    exp_47_ram[2207] = 244;
    exp_47_ram[2208] = 132;
    exp_47_ram[2209] = 95;
    exp_47_ram[2210] = 0;
    exp_47_ram[2211] = 95;
    exp_47_ram[2212] = 5;
    exp_47_ram[2213] = 244;
    exp_47_ram[2214] = 4;
    exp_47_ram[2215] = 196;
    exp_47_ram[2216] = 132;
    exp_47_ram[2217] = 7;
    exp_47_ram[2218] = 7;
    exp_47_ram[2219] = 192;
    exp_47_ram[2220] = 95;
    exp_47_ram[2221] = 68;
    exp_47_ram[2222] = 23;
    exp_47_ram[2223] = 244;
    exp_47_ram[2224] = 68;
    exp_47_ram[2225] = 48;
    exp_47_ram[2226] = 231;
    exp_47_ram[2227] = 4;
    exp_47_ram[2228] = 159;
    exp_47_ram[2229] = 196;
    exp_47_ram[2230] = 31;
    exp_47_ram[2231] = 132;
    exp_47_ram[2232] = 159;
    exp_47_ram[2233] = 193;
    exp_47_ram[2234] = 129;
    exp_47_ram[2235] = 1;
    exp_47_ram[2236] = 0;
    exp_47_ram[2237] = 1;
    exp_47_ram[2238] = 17;
    exp_47_ram[2239] = 129;
    exp_47_ram[2240] = 1;
    exp_47_ram[2241] = 128;
    exp_47_ram[2242] = 79;
    exp_47_ram[2243] = 128;
    exp_47_ram[2244] = 207;
    exp_47_ram[2245] = 128;
    exp_47_ram[2246] = 79;
    exp_47_ram[2247] = 128;
    exp_47_ram[2248] = 207;
    exp_47_ram[2249] = 128;
    exp_47_ram[2250] = 79;
    exp_47_ram[2251] = 0;
    exp_47_ram[2252] = 207;
    exp_47_ram[2253] = 79;
    exp_47_ram[2254] = 5;
    exp_47_ram[2255] = 244;
    exp_47_ram[2256] = 244;
    exp_47_ram[2257] = 247;
    exp_47_ram[2258] = 64;
    exp_47_ram[2259] = 247;
    exp_47_ram[2260] = 39;
    exp_47_ram[2261] = 0;
    exp_47_ram[2262] = 71;
    exp_47_ram[2263] = 247;
    exp_47_ram[2264] = 7;
    exp_47_ram[2265] = 7;
    exp_47_ram[2266] = 15;
    exp_47_ram[2267] = 64;
    exp_47_ram[2268] = 79;
    exp_47_ram[2269] = 192;
    exp_47_ram[2270] = 15;
    exp_47_ram[2271] = 64;
    exp_47_ram[2272] = 95;
    exp_47_ram[2273] = 192;
    exp_47_ram[2274] = 31;
    exp_47_ram[2275] = 0;
    exp_47_ram[2276] = 95;
    exp_47_ram[2277] = 5;
    exp_47_ram[2278] = 5;
    exp_47_ram[2279] = 181;
    exp_47_ram[2280] = 1;
    exp_47_ram[2281] = 183;
    exp_47_ram[2282] = 7;
    exp_47_ram[2283] = 5;
    exp_47_ram[2284] = 21;
    exp_47_ram[2285] = 245;
    exp_47_ram[2286] = 1;
    exp_47_ram[2287] = 0;
    exp_47_ram[2288] = 176;
    exp_47_ram[2289] = 245;
    exp_47_ram[2290] = 245;
    exp_47_ram[2291] = 223;
    exp_47_ram[2292] = 250;
    exp_47_ram[2293] = 0;
    exp_47_ram[2294] = 0;
    exp_47_ram[2295] = 0;
    exp_47_ram[2296] = 0;
    exp_47_ram[2297] = 110;
    exp_47_ram[2298] = 84;
    exp_47_ram[2299] = 101;
    exp_47_ram[2300] = 117;
    exp_47_ram[2301] = 83;
    exp_47_ram[2302] = 0;
    exp_47_ram[2303] = 110;
    exp_47_ram[2304] = 77;
    exp_47_ram[2305] = 112;
    exp_47_ram[2306] = 121;
    exp_47_ram[2307] = 74;
    exp_47_ram[2308] = 117;
    exp_47_ram[2309] = 112;
    exp_47_ram[2310] = 78;
    exp_47_ram[2311] = 101;
    exp_47_ram[2312] = 0;
    exp_47_ram[2313] = 0;
    exp_47_ram[2314] = 0;
    exp_47_ram[2315] = 0;
    exp_47_ram[2316] = 0;
    exp_47_ram[2317] = 0;
    exp_47_ram[2318] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 65;
    exp_40_ram[32] = 1;
    exp_40_ram[33] = 32;
    exp_40_ram[34] = 0;
    exp_40_ram[35] = 8;
    exp_40_ram[36] = 135;
    exp_40_ram[37] = 8;
    exp_40_ram[38] = 133;
    exp_40_ram[39] = 131;
    exp_40_ram[40] = 146;
    exp_40_ram[41] = 6;
    exp_40_ram[42] = 246;
    exp_40_ram[43] = 7;
    exp_40_ram[44] = 120;
    exp_40_ram[45] = 7;
    exp_40_ram[46] = 55;
    exp_40_ram[47] = 23;
    exp_40_ram[48] = 85;
    exp_40_ram[49] = 134;
    exp_40_ram[50] = 198;
    exp_40_ram[51] = 5;
    exp_40_ram[52] = 135;
    exp_40_ram[53] = 6;
    exp_40_ram[54] = 12;
    exp_40_ram[55] = 149;
    exp_40_ram[56] = 215;
    exp_40_ram[57] = 24;
    exp_40_ram[58] = 101;
    exp_40_ram[59] = 147;
    exp_40_ram[60] = 88;
    exp_40_ram[61] = 214;
    exp_40_ram[62] = 22;
    exp_40_ram[63] = 86;
    exp_40_ram[64] = 87;
    exp_40_ram[65] = 247;
    exp_40_ram[66] = 133;
    exp_40_ram[67] = 5;
    exp_40_ram[68] = 23;
    exp_40_ram[69] = 103;
    exp_40_ram[70] = 254;
    exp_40_ram[71] = 135;
    exp_40_ram[72] = 133;
    exp_40_ram[73] = 232;
    exp_40_ram[74] = 246;
    exp_40_ram[75] = 133;
    exp_40_ram[76] = 135;
    exp_40_ram[77] = 135;
    exp_40_ram[78] = 247;
    exp_40_ram[79] = 19;
    exp_40_ram[80] = 83;
    exp_40_ram[81] = 215;
    exp_40_ram[82] = 23;
    exp_40_ram[83] = 99;
    exp_40_ram[84] = 6;
    exp_40_ram[85] = 134;
    exp_40_ram[86] = 124;
    exp_40_ram[87] = 3;
    exp_40_ram[88] = 134;
    exp_40_ram[89] = 102;
    exp_40_ram[90] = 116;
    exp_40_ram[91] = 134;
    exp_40_ram[92] = 21;
    exp_40_ram[93] = 101;
    exp_40_ram[94] = 5;
    exp_40_ram[95] = 0;
    exp_40_ram[96] = 5;
    exp_40_ram[97] = 7;
    exp_40_ram[98] = 108;
    exp_40_ram[99] = 7;
    exp_40_ram[100] = 240;
    exp_40_ram[101] = 22;
    exp_40_ram[102] = 7;
    exp_40_ram[103] = 88;
    exp_40_ram[104] = 7;
    exp_40_ram[105] = 112;
    exp_40_ram[106] = 7;
    exp_40_ram[107] = 116;
    exp_40_ram[108] = 5;
    exp_40_ram[109] = 87;
    exp_40_ram[110] = 134;
    exp_40_ram[111] = 199;
    exp_40_ram[112] = 6;
    exp_40_ram[113] = 7;
    exp_40_ram[114] = 6;
    exp_40_ram[115] = 22;
    exp_40_ram[116] = 135;
    exp_40_ram[117] = 5;
    exp_40_ram[118] = 88;
    exp_40_ram[119] = 22;
    exp_40_ram[120] = 86;
    exp_40_ram[121] = 87;
    exp_40_ram[122] = 246;
    exp_40_ram[123] = 215;
    exp_40_ram[124] = 150;
    exp_40_ram[125] = 231;
    exp_40_ram[126] = 14;
    exp_40_ram[127] = 133;
    exp_40_ram[128] = 126;
    exp_40_ram[129] = 7;
    exp_40_ram[130] = 133;
    exp_40_ram[131] = 104;
    exp_40_ram[132] = 118;
    exp_40_ram[133] = 133;
    exp_40_ram[134] = 7;
    exp_40_ram[135] = 7;
    exp_40_ram[136] = 119;
    exp_40_ram[137] = 19;
    exp_40_ram[138] = 83;
    exp_40_ram[139] = 87;
    exp_40_ram[140] = 151;
    exp_40_ram[141] = 227;
    exp_40_ram[142] = 6;
    exp_40_ram[143] = 6;
    exp_40_ram[144] = 124;
    exp_40_ram[145] = 3;
    exp_40_ram[146] = 6;
    exp_40_ram[147] = 102;
    exp_40_ram[148] = 116;
    exp_40_ram[149] = 6;
    exp_40_ram[150] = 21;
    exp_40_ram[151] = 101;
    exp_40_ram[152] = 128;
    exp_40_ram[153] = 7;
    exp_40_ram[154] = 5;
    exp_40_ram[155] = 100;
    exp_40_ram[156] = 5;
    exp_40_ram[157] = 240;
    exp_40_ram[158] = 24;
    exp_40_ram[159] = 213;
    exp_40_ram[160] = 147;
    exp_40_ram[161] = 151;
    exp_40_ram[162] = 215;
    exp_40_ram[163] = 88;
    exp_40_ram[164] = 102;
    exp_40_ram[165] = 119;
    exp_40_ram[166] = 23;
    exp_40_ram[167] = 215;
    exp_40_ram[168] = 85;
    exp_40_ram[169] = 85;
    exp_40_ram[170] = 23;
    exp_40_ram[171] = 103;
    exp_40_ram[172] = 134;
    exp_40_ram[173] = 5;
    exp_40_ram[174] = 126;
    exp_40_ram[175] = 7;
    exp_40_ram[176] = 5;
    exp_40_ram[177] = 104;
    exp_40_ram[178] = 118;
    exp_40_ram[179] = 5;
    exp_40_ram[180] = 7;
    exp_40_ram[181] = 6;
    exp_40_ram[182] = 247;
    exp_40_ram[183] = 22;
    exp_40_ram[184] = 86;
    exp_40_ram[185] = 214;
    exp_40_ram[186] = 23;
    exp_40_ram[187] = 133;
    exp_40_ram[188] = 103;
    exp_40_ram[189] = 135;
    exp_40_ram[190] = 254;
    exp_40_ram[191] = 135;
    exp_40_ram[192] = 135;
    exp_40_ram[193] = 232;
    exp_40_ram[194] = 246;
    exp_40_ram[195] = 135;
    exp_40_ram[196] = 135;
    exp_40_ram[197] = 149;
    exp_40_ram[198] = 135;
    exp_40_ram[199] = 229;
    exp_40_ram[200] = 240;
    exp_40_ram[201] = 228;
    exp_40_ram[202] = 7;
    exp_40_ram[203] = 242;
    exp_40_ram[204] = 7;
    exp_40_ram[205] = 53;
    exp_40_ram[206] = 149;
    exp_40_ram[207] = 213;
    exp_40_ram[208] = 7;
    exp_40_ram[209] = 7;
    exp_40_ram[210] = 71;
    exp_40_ram[211] = 5;
    exp_40_ram[212] = 7;
    exp_40_ram[213] = 5;
    exp_40_ram[214] = 22;
    exp_40_ram[215] = 5;
    exp_40_ram[216] = 224;
    exp_40_ram[217] = 181;
    exp_40_ram[218] = 69;
    exp_40_ram[219] = 240;
    exp_40_ram[220] = 7;
    exp_40_ram[221] = 5;
    exp_40_ram[222] = 226;
    exp_40_ram[223] = 5;
    exp_40_ram[224] = 240;
    exp_40_ram[225] = 88;
    exp_40_ram[226] = 150;
    exp_40_ram[227] = 104;
    exp_40_ram[228] = 222;
    exp_40_ram[229] = 94;
    exp_40_ram[230] = 118;
    exp_40_ram[231] = 151;
    exp_40_ram[232] = 215;
    exp_40_ram[233] = 19;
    exp_40_ram[234] = 102;
    exp_40_ram[235] = 23;
    exp_40_ram[236] = 215;
    exp_40_ram[237] = 87;
    exp_40_ram[238] = 94;
    exp_40_ram[239] = 150;
    exp_40_ram[240] = 231;
    exp_40_ram[241] = 143;
    exp_40_ram[242] = 5;
    exp_40_ram[243] = 126;
    exp_40_ram[244] = 7;
    exp_40_ram[245] = 5;
    exp_40_ram[246] = 104;
    exp_40_ram[247] = 118;
    exp_40_ram[248] = 5;
    exp_40_ram[249] = 7;
    exp_40_ram[250] = 7;
    exp_40_ram[251] = 118;
    exp_40_ram[252] = 87;
    exp_40_ram[253] = 150;
    exp_40_ram[254] = 142;
    exp_40_ram[255] = 23;
    exp_40_ram[256] = 215;
    exp_40_ram[257] = 231;
    exp_40_ram[258] = 6;
    exp_40_ram[259] = 254;
    exp_40_ram[260] = 135;
    exp_40_ram[261] = 6;
    exp_40_ram[262] = 232;
    exp_40_ram[263] = 246;
    exp_40_ram[264] = 6;
    exp_40_ram[265] = 135;
    exp_40_ram[266] = 21;
    exp_40_ram[267] = 14;
    exp_40_ram[268] = 101;
    exp_40_ram[269] = 134;
    exp_40_ram[270] = 120;
    exp_40_ram[271] = 86;
    exp_40_ram[272] = 118;
    exp_40_ram[273] = 83;
    exp_40_ram[274] = 135;
    exp_40_ram[275] = 14;
    exp_40_ram[276] = 6;
    exp_40_ram[277] = 87;
    exp_40_ram[278] = 8;
    exp_40_ram[279] = 8;
    exp_40_ram[280] = 7;
    exp_40_ram[281] = 6;
    exp_40_ram[282] = 116;
    exp_40_ram[283] = 6;
    exp_40_ram[284] = 86;
    exp_40_ram[285] = 134;
    exp_40_ram[286] = 230;
    exp_40_ram[287] = 158;
    exp_40_ram[288] = 7;
    exp_40_ram[289] = 135;
    exp_40_ram[290] = 119;
    exp_40_ram[291] = 23;
    exp_40_ram[292] = 126;
    exp_40_ram[293] = 152;
    exp_40_ram[294] = 7;
    exp_40_ram[295] = 5;
    exp_40_ram[296] = 240;
    exp_40_ram[297] = 5;
    exp_40_ram[298] = 240;
    exp_40_ram[299] = 5;
    exp_40_ram[300] = 5;
    exp_40_ram[301] = 240;
    exp_40_ram[302] = 6;
    exp_40_ram[303] = 5;
    exp_40_ram[304] = 246;
    exp_40_ram[305] = 132;
    exp_40_ram[306] = 5;
    exp_40_ram[307] = 213;
    exp_40_ram[308] = 22;
    exp_40_ram[309] = 150;
    exp_40_ram[310] = 128;
    exp_40_ram[311] = 64;
    exp_40_ram[312] = 198;
    exp_40_ram[313] = 134;
    exp_40_ram[314] = 5;
    exp_40_ram[315] = 5;
    exp_40_ram[316] = 12;
    exp_40_ram[317] = 6;
    exp_40_ram[318] = 122;
    exp_40_ram[319] = 88;
    exp_40_ram[320] = 22;
    exp_40_ram[321] = 150;
    exp_40_ram[322] = 106;
    exp_40_ram[323] = 5;
    exp_40_ram[324] = 230;
    exp_40_ram[325] = 133;
    exp_40_ram[326] = 101;
    exp_40_ram[327] = 214;
    exp_40_ram[328] = 86;
    exp_40_ram[329] = 150;
    exp_40_ram[330] = 128;
    exp_40_ram[331] = 130;
    exp_40_ram[332] = 240;
    exp_40_ram[333] = 133;
    exp_40_ram[334] = 128;
    exp_40_ram[335] = 5;
    exp_40_ram[336] = 72;
    exp_40_ram[337] = 5;
    exp_40_ram[338] = 240;
    exp_40_ram[339] = 5;
    exp_40_ram[340] = 130;
    exp_40_ram[341] = 240;
    exp_40_ram[342] = 5;
    exp_40_ram[343] = 128;
    exp_40_ram[344] = 130;
    exp_40_ram[345] = 202;
    exp_40_ram[346] = 76;
    exp_40_ram[347] = 240;
    exp_40_ram[348] = 133;
    exp_40_ram[349] = 128;
    exp_40_ram[350] = 5;
    exp_40_ram[351] = 88;
    exp_40_ram[352] = 5;
    exp_40_ram[353] = 240;
    exp_40_ram[354] = 5;
    exp_40_ram[355] = 128;
    exp_40_ram[356] = 101;
    exp_40_ram[357] = 32;
    exp_40_ram[358] = 108;
    exp_40_ram[359] = 0;
    exp_40_ram[360] = 117;
    exp_40_ram[361] = 110;
    exp_40_ram[362] = 110;
    exp_40_ram[363] = 116;
    exp_40_ram[364] = 100;
    exp_40_ram[365] = 100;
    exp_40_ram[366] = 46;
    exp_40_ram[367] = 0;
    exp_40_ram[368] = 117;
    exp_40_ram[369] = 117;
    exp_40_ram[370] = 45;
    exp_40_ram[371] = 32;
    exp_40_ram[372] = 101;
    exp_40_ram[373] = 32;
    exp_40_ram[374] = 116;
    exp_40_ram[375] = 105;
    exp_40_ram[376] = 105;
    exp_40_ram[377] = 32;
    exp_40_ram[378] = 111;
    exp_40_ram[379] = 0;
    exp_40_ram[380] = 117;
    exp_40_ram[381] = 45;
    exp_40_ram[382] = 32;
    exp_40_ram[383] = 101;
    exp_40_ram[384] = 32;
    exp_40_ram[385] = 116;
    exp_40_ram[386] = 105;
    exp_40_ram[387] = 105;
    exp_40_ram[388] = 32;
    exp_40_ram[389] = 111;
    exp_40_ram[390] = 0;
    exp_40_ram[391] = 117;
    exp_40_ram[392] = 45;
    exp_40_ram[393] = 32;
    exp_40_ram[394] = 101;
    exp_40_ram[395] = 32;
    exp_40_ram[396] = 105;
    exp_40_ram[397] = 32;
    exp_40_ram[398] = 49;
    exp_40_ram[399] = 99;
    exp_40_ram[400] = 10;
    exp_40_ram[401] = 117;
    exp_40_ram[402] = 45;
    exp_40_ram[403] = 32;
    exp_40_ram[404] = 101;
    exp_40_ram[405] = 32;
    exp_40_ram[406] = 105;
    exp_40_ram[407] = 32;
    exp_40_ram[408] = 49;
    exp_40_ram[409] = 99;
    exp_40_ram[410] = 10;
    exp_40_ram[411] = 108;
    exp_40_ram[412] = 109;
    exp_40_ram[413] = 32;
    exp_40_ram[414] = 46;
    exp_40_ram[415] = 97;
    exp_40_ram[416] = 0;
    exp_40_ram[417] = 97;
    exp_40_ram[418] = 0;
    exp_40_ram[419] = 108;
    exp_40_ram[420] = 97;
    exp_40_ram[421] = 32;
    exp_40_ram[422] = 120;
    exp_40_ram[423] = 56;
    exp_40_ram[424] = 48;
    exp_40_ram[425] = 0;
    exp_40_ram[426] = 67;
    exp_40_ram[427] = 115;
    exp_40_ram[428] = 68;
    exp_40_ram[429] = 0;
    exp_40_ram[430] = 97;
    exp_40_ram[431] = 101;
    exp_40_ram[432] = 32;
    exp_40_ram[433] = 108;
    exp_40_ram[434] = 41;
    exp_40_ram[435] = 105;
    exp_40_ram[436] = 32;
    exp_40_ram[437] = 101;
    exp_40_ram[438] = 41;
    exp_40_ram[439] = 111;
    exp_40_ram[440] = 97;
    exp_40_ram[441] = 0;
    exp_40_ram[442] = 41;
    exp_40_ram[443] = 115;
    exp_40_ram[444] = 117;
    exp_40_ram[445] = 112;
    exp_40_ram[446] = 97;
    exp_40_ram[447] = 110;
    exp_40_ram[448] = 41;
    exp_40_ram[449] = 115;
    exp_40_ram[450] = 101;
    exp_40_ram[451] = 121;
    exp_40_ram[452] = 1;
    exp_40_ram[453] = 3;
    exp_40_ram[454] = 4;
    exp_40_ram[455] = 4;
    exp_40_ram[456] = 5;
    exp_40_ram[457] = 5;
    exp_40_ram[458] = 5;
    exp_40_ram[459] = 5;
    exp_40_ram[460] = 6;
    exp_40_ram[461] = 6;
    exp_40_ram[462] = 6;
    exp_40_ram[463] = 6;
    exp_40_ram[464] = 6;
    exp_40_ram[465] = 6;
    exp_40_ram[466] = 6;
    exp_40_ram[467] = 6;
    exp_40_ram[468] = 7;
    exp_40_ram[469] = 7;
    exp_40_ram[470] = 7;
    exp_40_ram[471] = 7;
    exp_40_ram[472] = 7;
    exp_40_ram[473] = 7;
    exp_40_ram[474] = 7;
    exp_40_ram[475] = 7;
    exp_40_ram[476] = 7;
    exp_40_ram[477] = 7;
    exp_40_ram[478] = 7;
    exp_40_ram[479] = 7;
    exp_40_ram[480] = 7;
    exp_40_ram[481] = 7;
    exp_40_ram[482] = 7;
    exp_40_ram[483] = 7;
    exp_40_ram[484] = 8;
    exp_40_ram[485] = 8;
    exp_40_ram[486] = 8;
    exp_40_ram[487] = 8;
    exp_40_ram[488] = 8;
    exp_40_ram[489] = 8;
    exp_40_ram[490] = 8;
    exp_40_ram[491] = 8;
    exp_40_ram[492] = 8;
    exp_40_ram[493] = 8;
    exp_40_ram[494] = 8;
    exp_40_ram[495] = 8;
    exp_40_ram[496] = 8;
    exp_40_ram[497] = 8;
    exp_40_ram[498] = 8;
    exp_40_ram[499] = 8;
    exp_40_ram[500] = 8;
    exp_40_ram[501] = 8;
    exp_40_ram[502] = 8;
    exp_40_ram[503] = 8;
    exp_40_ram[504] = 8;
    exp_40_ram[505] = 8;
    exp_40_ram[506] = 8;
    exp_40_ram[507] = 8;
    exp_40_ram[508] = 8;
    exp_40_ram[509] = 8;
    exp_40_ram[510] = 8;
    exp_40_ram[511] = 8;
    exp_40_ram[512] = 8;
    exp_40_ram[513] = 8;
    exp_40_ram[514] = 8;
    exp_40_ram[515] = 8;
    exp_40_ram[516] = 160;
    exp_40_ram[517] = 128;
    exp_40_ram[518] = 39;
    exp_40_ram[519] = 167;
    exp_40_ram[520] = 165;
    exp_40_ram[521] = 128;
    exp_40_ram[522] = 7;
    exp_40_ram[523] = 5;
    exp_40_ram[524] = 135;
    exp_40_ram[525] = 71;
    exp_40_ram[526] = 20;
    exp_40_ram[527] = 128;
    exp_40_ram[528] = 5;
    exp_40_ram[529] = 160;
    exp_40_ram[530] = 240;
    exp_40_ram[531] = 1;
    exp_40_ram[532] = 39;
    exp_40_ram[533] = 36;
    exp_40_ram[534] = 164;
    exp_40_ram[535] = 38;
    exp_40_ram[536] = 5;
    exp_40_ram[537] = 240;
    exp_40_ram[538] = 7;
    exp_40_ram[539] = 32;
    exp_40_ram[540] = 32;
    exp_40_ram[541] = 36;
    exp_40_ram[542] = 5;
    exp_40_ram[543] = 1;
    exp_40_ram[544] = 128;
    exp_40_ram[545] = 1;
    exp_40_ram[546] = 36;
    exp_40_ram[547] = 38;
    exp_40_ram[548] = 132;
    exp_40_ram[549] = 142;
    exp_40_ram[550] = 240;
    exp_40_ram[551] = 32;
    exp_40_ram[552] = 5;
    exp_40_ram[553] = 36;
    exp_40_ram[554] = 1;
    exp_40_ram[555] = 128;
    exp_40_ram[556] = 6;
    exp_40_ram[557] = 128;
    exp_40_ram[558] = 6;
    exp_40_ram[559] = 0;
    exp_40_ram[560] = 240;
    exp_40_ram[561] = 1;
    exp_40_ram[562] = 44;
    exp_40_ram[563] = 42;
    exp_40_ram[564] = 40;
    exp_40_ram[565] = 38;
    exp_40_ram[566] = 36;
    exp_40_ram[567] = 44;
    exp_40_ram[568] = 42;
    exp_40_ram[569] = 137;
    exp_40_ram[570] = 46;
    exp_40_ram[571] = 34;
    exp_40_ram[572] = 32;
    exp_40_ram[573] = 46;
    exp_40_ram[574] = 40;
    exp_40_ram[575] = 38;
    exp_40_ram[576] = 7;
    exp_40_ram[577] = 4;
    exp_40_ram[578] = 132;
    exp_40_ram[579] = 5;
    exp_40_ram[580] = 140;
    exp_40_ram[581] = 9;
    exp_40_ram[582] = 12;
    exp_40_ram[583] = 138;
    exp_40_ram[584] = 0;
    exp_40_ram[585] = 7;
    exp_40_ram[586] = 18;
    exp_40_ram[587] = 13;
    exp_40_ram[588] = 11;
    exp_40_ram[589] = 13;
    exp_40_ram[590] = 11;
    exp_40_ram[591] = 10;
    exp_40_ram[592] = 0;
    exp_40_ram[593] = 139;
    exp_40_ram[594] = 215;
    exp_40_ram[595] = 243;
    exp_40_ram[596] = 22;
    exp_40_ram[597] = 148;
    exp_40_ram[598] = 22;
    exp_40_ram[599] = 247;
    exp_40_ram[600] = 104;
    exp_40_ram[601] = 3;
    exp_40_ram[602] = 115;
    exp_40_ram[603] = 6;
    exp_40_ram[604] = 134;
    exp_40_ram[605] = 5;
    exp_40_ram[606] = 5;
    exp_40_ram[607] = 240;
    exp_40_ram[608] = 13;
    exp_40_ram[609] = 252;
    exp_40_ram[610] = 13;
    exp_40_ram[611] = 215;
    exp_40_ram[612] = 250;
    exp_40_ram[613] = 32;
    exp_40_ram[614] = 36;
    exp_40_ram[615] = 36;
    exp_40_ram[616] = 41;
    exp_40_ram[617] = 41;
    exp_40_ram[618] = 42;
    exp_40_ram[619] = 42;
    exp_40_ram[620] = 43;
    exp_40_ram[621] = 43;
    exp_40_ram[622] = 44;
    exp_40_ram[623] = 44;
    exp_40_ram[624] = 45;
    exp_40_ram[625] = 45;
    exp_40_ram[626] = 1;
    exp_40_ram[627] = 128;
    exp_40_ram[628] = 6;
    exp_40_ram[629] = 3;
    exp_40_ram[630] = 240;
    exp_40_ram[631] = 3;
    exp_40_ram[632] = 240;
    exp_40_ram[633] = 96;
    exp_40_ram[634] = 6;
    exp_40_ram[635] = 134;
    exp_40_ram[636] = 5;
    exp_40_ram[637] = 133;
    exp_40_ram[638] = 240;
    exp_40_ram[639] = 240;
    exp_40_ram[640] = 13;
    exp_40_ram[641] = 11;
    exp_40_ram[642] = 240;
    exp_40_ram[643] = 219;
    exp_40_ram[644] = 13;
    exp_40_ram[645] = 139;
    exp_40_ram[646] = 12;
    exp_40_ram[647] = 240;
    exp_40_ram[648] = 71;
    exp_40_ram[649] = 138;
    exp_40_ram[650] = 1;
    exp_40_ram[651] = 36;
    exp_40_ram[652] = 34;
    exp_40_ram[653] = 46;
    exp_40_ram[654] = 42;
    exp_40_ram[655] = 40;
    exp_40_ram[656] = 38;
    exp_40_ram[657] = 34;
    exp_40_ram[658] = 32;
    exp_40_ram[659] = 46;
    exp_40_ram[660] = 9;
    exp_40_ram[661] = 38;
    exp_40_ram[662] = 32;
    exp_40_ram[663] = 44;
    exp_40_ram[664] = 36;
    exp_40_ram[665] = 4;
    exp_40_ram[666] = 132;
    exp_40_ram[667] = 140;
    exp_40_ram[668] = 6;
    exp_40_ram[669] = 7;
    exp_40_ram[670] = 10;
    exp_40_ram[671] = 13;
    exp_40_ram[672] = 13;
    exp_40_ram[673] = 11;
    exp_40_ram[674] = 11;
    exp_40_ram[675] = 135;
    exp_40_ram[676] = 197;
    exp_40_ram[677] = 9;
    exp_40_ram[678] = 138;
    exp_40_ram[679] = 18;
    exp_40_ram[680] = 71;
    exp_40_ram[681] = 142;
    exp_40_ram[682] = 6;
    exp_40_ram[683] = 156;
    exp_40_ram[684] = 9;
    exp_40_ram[685] = 135;
    exp_40_ram[686] = 71;
    exp_40_ram[687] = 22;
    exp_40_ram[688] = 32;
    exp_40_ram[689] = 36;
    exp_40_ram[690] = 36;
    exp_40_ram[691] = 41;
    exp_40_ram[692] = 41;
    exp_40_ram[693] = 42;
    exp_40_ram[694] = 42;
    exp_40_ram[695] = 43;
    exp_40_ram[696] = 43;
    exp_40_ram[697] = 44;
    exp_40_ram[698] = 44;
    exp_40_ram[699] = 45;
    exp_40_ram[700] = 45;
    exp_40_ram[701] = 5;
    exp_40_ram[702] = 1;
    exp_40_ram[703] = 128;
    exp_40_ram[704] = 6;
    exp_40_ram[705] = 5;
    exp_40_ram[706] = 134;
    exp_40_ram[707] = 240;
    exp_40_ram[708] = 6;
    exp_40_ram[709] = 71;
    exp_40_ram[710] = 132;
    exp_40_ram[711] = 7;
    exp_40_ram[712] = 240;
    exp_40_ram[713] = 7;
    exp_40_ram[714] = 7;
    exp_40_ram[715] = 134;
    exp_40_ram[716] = 198;
    exp_40_ram[717] = 9;
    exp_40_ram[718] = 138;
    exp_40_ram[719] = 133;
    exp_40_ram[720] = 120;
    exp_40_ram[721] = 132;
    exp_40_ram[722] = 108;
    exp_40_ram[723] = 5;
    exp_40_ram[724] = 134;
    exp_40_ram[725] = 232;
    exp_40_ram[726] = 136;
    exp_40_ram[727] = 5;
    exp_40_ram[728] = 154;
    exp_40_ram[729] = 140;
    exp_40_ram[730] = 8;
    exp_40_ram[731] = 0;
    exp_40_ram[732] = 7;
    exp_40_ram[733] = 70;
    exp_40_ram[734] = 135;
    exp_40_ram[735] = 152;
    exp_40_ram[736] = 240;
    exp_40_ram[737] = 5;
    exp_40_ram[738] = 150;
    exp_40_ram[739] = 140;
    exp_40_ram[740] = 172;
    exp_40_ram[741] = 216;
    exp_40_ram[742] = 6;
    exp_40_ram[743] = 5;
    exp_40_ram[744] = 134;
    exp_40_ram[745] = 5;
    exp_40_ram[746] = 38;
    exp_40_ram[747] = 36;
    exp_40_ram[748] = 240;
    exp_40_ram[749] = 39;
    exp_40_ram[750] = 39;
    exp_40_ram[751] = 6;
    exp_40_ram[752] = 8;
    exp_40_ram[753] = 8;
    exp_40_ram[754] = 7;
    exp_40_ram[755] = 6;
    exp_40_ram[756] = 133;
    exp_40_ram[757] = 5;
    exp_40_ram[758] = 240;
    exp_40_ram[759] = 0;
    exp_40_ram[760] = 138;
    exp_40_ram[761] = 230;
    exp_40_ram[762] = 5;
    exp_40_ram[763] = 142;
    exp_40_ram[764] = 7;
    exp_40_ram[765] = 144;
    exp_40_ram[766] = 172;
    exp_40_ram[767] = 135;
    exp_40_ram[768] = 69;
    exp_40_ram[769] = 30;
    exp_40_ram[770] = 140;
    exp_40_ram[771] = 240;
    exp_40_ram[772] = 5;
    exp_40_ram[773] = 144;
    exp_40_ram[774] = 140;
    exp_40_ram[775] = 8;
    exp_40_ram[776] = 8;
    exp_40_ram[777] = 0;
    exp_40_ram[778] = 6;
    exp_40_ram[779] = 5;
    exp_40_ram[780] = 134;
    exp_40_ram[781] = 5;
    exp_40_ram[782] = 240;
    exp_40_ram[783] = 197;
    exp_40_ram[784] = 6;
    exp_40_ram[785] = 5;
    exp_40_ram[786] = 134;
    exp_40_ram[787] = 140;
    exp_40_ram[788] = 240;
    exp_40_ram[789] = 6;
    exp_40_ram[790] = 12;
    exp_40_ram[791] = 240;
    exp_40_ram[792] = 6;
    exp_40_ram[793] = 5;
    exp_40_ram[794] = 134;
    exp_40_ram[795] = 36;
    exp_40_ram[796] = 240;
    exp_40_ram[797] = 39;
    exp_40_ram[798] = 6;
    exp_40_ram[799] = 12;
    exp_40_ram[800] = 240;
    exp_40_ram[801] = 8;
    exp_40_ram[802] = 8;
    exp_40_ram[803] = 134;
    exp_40_ram[804] = 240;
    exp_40_ram[805] = 140;
    exp_40_ram[806] = 8;
    exp_40_ram[807] = 8;
    exp_40_ram[808] = 166;
    exp_40_ram[809] = 240;
    exp_40_ram[810] = 140;
    exp_40_ram[811] = 8;
    exp_40_ram[812] = 8;
    exp_40_ram[813] = 240;
    exp_40_ram[814] = 6;
    exp_40_ram[815] = 5;
    exp_40_ram[816] = 128;
    exp_40_ram[817] = 1;
    exp_40_ram[818] = 42;
    exp_40_ram[819] = 39;
    exp_40_ram[820] = 36;
    exp_40_ram[821] = 6;
    exp_40_ram[822] = 165;
    exp_40_ram[823] = 34;
    exp_40_ram[824] = 38;
    exp_40_ram[825] = 5;
    exp_40_ram[826] = 6;
    exp_40_ram[827] = 46;
    exp_40_ram[828] = 40;
    exp_40_ram[829] = 44;
    exp_40_ram[830] = 46;
    exp_40_ram[831] = 38;
    exp_40_ram[832] = 240;
    exp_40_ram[833] = 32;
    exp_40_ram[834] = 1;
    exp_40_ram[835] = 128;
    exp_40_ram[836] = 7;
    exp_40_ram[837] = 215;
    exp_40_ram[838] = 37;
    exp_40_ram[839] = 5;
    exp_40_ram[840] = 154;
    exp_40_ram[841] = 7;
    exp_40_ram[842] = 23;
    exp_40_ram[843] = 5;
    exp_40_ram[844] = 128;
    exp_40_ram[845] = 39;
    exp_40_ram[846] = 35;
    exp_40_ram[847] = 39;
    exp_40_ram[848] = 22;
    exp_40_ram[849] = 7;
    exp_40_ram[850] = 32;
    exp_40_ram[851] = 8;
    exp_40_ram[852] = 7;
    exp_40_ram[853] = 136;
    exp_40_ram[854] = 5;
    exp_40_ram[855] = 84;
    exp_40_ram[856] = 22;
    exp_40_ram[857] = 6;
    exp_40_ram[858] = 168;
    exp_40_ram[859] = 118;
    exp_40_ram[860] = 102;
    exp_40_ram[861] = 120;
    exp_40_ram[862] = 8;
    exp_40_ram[863] = 7;
    exp_40_ram[864] = 7;
    exp_40_ram[865] = 240;
    exp_40_ram[866] = 229;
    exp_40_ram[867] = 160;
    exp_40_ram[868] = 240;
    exp_40_ram[869] = 134;
    exp_40_ram[870] = 134;
    exp_40_ram[871] = 150;
    exp_40_ram[872] = 199;
    exp_40_ram[873] = 6;
    exp_40_ram[874] = 135;
    exp_40_ram[875] = 160;
    exp_40_ram[876] = 7;
    exp_40_ram[877] = 240;
    exp_40_ram[878] = 38;
    exp_40_ram[879] = 7;
    exp_40_ram[880] = 5;
    exp_40_ram[881] = 117;
    exp_40_ram[882] = 5;
    exp_40_ram[883] = 133;
    exp_40_ram[884] = 39;
    exp_40_ram[885] = 5;
    exp_40_ram[886] = 133;
    exp_40_ram[887] = 247;
    exp_40_ram[888] = 32;
    exp_40_ram[889] = 39;
    exp_40_ram[890] = 168;
    exp_40_ram[891] = 6;
    exp_40_ram[892] = 7;
    exp_40_ram[893] = 3;
    exp_40_ram[894] = 135;
    exp_40_ram[895] = 208;
    exp_40_ram[896] = 150;
    exp_40_ram[897] = 6;
    exp_40_ram[898] = 165;
    exp_40_ram[899] = 118;
    exp_40_ram[900] = 135;
    exp_40_ram[901] = 117;
    exp_40_ram[902] = 135;
    exp_40_ram[903] = 30;
    exp_40_ram[904] = 23;
    exp_40_ram[905] = 7;
    exp_40_ram[906] = 218;
    exp_40_ram[907] = 149;
    exp_40_ram[908] = 5;
    exp_40_ram[909] = 40;
    exp_40_ram[910] = 117;
    exp_40_ram[911] = 120;
    exp_40_ram[912] = 28;
    exp_40_ram[913] = 6;
    exp_40_ram[914] = 134;
    exp_40_ram[915] = 5;
    exp_40_ram[916] = 32;
    exp_40_ram[917] = 135;
    exp_40_ram[918] = 240;
    exp_40_ram[919] = 128;
    exp_40_ram[920] = 103;
    exp_40_ram[921] = 247;
    exp_40_ram[922] = 6;
    exp_40_ram[923] = 152;
    exp_40_ram[924] = 135;
    exp_40_ram[925] = 131;
    exp_40_ram[926] = 8;
    exp_40_ram[927] = 0;
    exp_40_ram[928] = 40;
    exp_40_ram[929] = 7;
    exp_40_ram[930] = 134;
    exp_40_ram[931] = 168;
    exp_40_ram[932] = 40;
    exp_40_ram[933] = 170;
    exp_40_ram[934] = 40;
    exp_40_ram[935] = 172;
    exp_40_ram[936] = 40;
    exp_40_ram[937] = 174;
    exp_40_ram[938] = 8;
    exp_40_ram[939] = 106;
    exp_40_ram[940] = 119;
    exp_40_ram[941] = 118;
    exp_40_ram[942] = 6;
    exp_40_ram[943] = 133;
    exp_40_ram[944] = 6;
    exp_40_ram[945] = 8;
    exp_40_ram[946] = 96;
    exp_40_ram[947] = 118;
    exp_40_ram[948] = 119;
    exp_40_ram[949] = 134;
    exp_40_ram[950] = 133;
    exp_40_ram[951] = 7;
    exp_40_ram[952] = 16;
    exp_40_ram[953] = 128;
    exp_40_ram[954] = 136;
    exp_40_ram[955] = 40;
    exp_40_ram[956] = 136;
    exp_40_ram[957] = 135;
    exp_40_ram[958] = 32;
    exp_40_ram[959] = 240;
    exp_40_ram[960] = 135;
    exp_40_ram[961] = 72;
    exp_40_ram[962] = 135;
    exp_40_ram[963] = 135;
    exp_40_ram[964] = 0;
    exp_40_ram[965] = 240;
    exp_40_ram[966] = 119;
    exp_40_ram[967] = 148;
    exp_40_ram[968] = 1;
    exp_40_ram[969] = 5;
    exp_40_ram[970] = 36;
    exp_40_ram[971] = 38;
    exp_40_ram[972] = 4;
    exp_40_ram[973] = 240;
    exp_40_ram[974] = 7;
    exp_40_ram[975] = 26;
    exp_40_ram[976] = 5;
    exp_40_ram[977] = 5;
    exp_40_ram[978] = 240;
    exp_40_ram[979] = 55;
    exp_40_ram[980] = 32;
    exp_40_ram[981] = 36;
    exp_40_ram[982] = 133;
    exp_40_ram[983] = 1;
    exp_40_ram[984] = 128;
    exp_40_ram[985] = 7;
    exp_40_ram[986] = 133;
    exp_40_ram[987] = 128;
    exp_40_ram[988] = 135;
    exp_40_ram[989] = 247;
    exp_40_ram[990] = 130;
    exp_40_ram[991] = 247;
    exp_40_ram[992] = 6;
    exp_40_ram[993] = 7;
    exp_40_ram[994] = 12;
    exp_40_ram[995] = 7;
    exp_40_ram[996] = 7;
    exp_40_ram[997] = 150;
    exp_40_ram[998] = 1;
    exp_40_ram[999] = 38;
    exp_40_ram[1000] = 240;
    exp_40_ram[1001] = 32;
    exp_40_ram[1002] = 55;
    exp_40_ram[1003] = 135;
    exp_40_ram[1004] = 133;
    exp_40_ram[1005] = 1;
    exp_40_ram[1006] = 128;
    exp_40_ram[1007] = 7;
    exp_40_ram[1008] = 133;
    exp_40_ram[1009] = 128;
    exp_40_ram[1010] = 7;
    exp_40_ram[1011] = 166;
    exp_40_ram[1012] = 166;
    exp_40_ram[1013] = 165;
    exp_40_ram[1014] = 5;
    exp_40_ram[1015] = 167;
    exp_40_ram[1016] = 229;
    exp_40_ram[1017] = 128;
    exp_40_ram[1018] = 1;
    exp_40_ram[1019] = 34;
    exp_40_ram[1020] = 42;
    exp_40_ram[1021] = 42;
    exp_40_ram[1022] = 84;
    exp_40_ram[1023] = 44;
    exp_40_ram[1024] = 40;
    exp_40_ram[1025] = 38;
    exp_40_ram[1026] = 36;
    exp_40_ram[1027] = 46;
    exp_40_ram[1028] = 32;
    exp_40_ram[1029] = 10;
    exp_40_ram[1030] = 4;
    exp_40_ram[1031] = 9;
    exp_40_ram[1032] = 9;
    exp_40_ram[1033] = 138;
    exp_40_ram[1034] = 132;
    exp_40_ram[1035] = 146;
    exp_40_ram[1036] = 43;
    exp_40_ram[1037] = 90;
    exp_40_ram[1038] = 4;
    exp_40_ram[1039] = 138;
    exp_40_ram[1040] = 0;
    exp_40_ram[1041] = 133;
    exp_40_ram[1042] = 5;
    exp_40_ram[1043] = 240;
    exp_40_ram[1044] = 133;
    exp_40_ram[1045] = 240;
    exp_40_ram[1046] = 5;
    exp_40_ram[1047] = 55;
    exp_40_ram[1048] = 137;
    exp_40_ram[1049] = 9;
    exp_40_ram[1050] = 132;
    exp_40_ram[1051] = 240;
    exp_40_ram[1052] = 5;
    exp_40_ram[1053] = 240;
    exp_40_ram[1054] = 53;
    exp_40_ram[1055] = 133;
    exp_40_ram[1056] = 5;
    exp_40_ram[1057] = 240;
    exp_40_ram[1058] = 5;
    exp_40_ram[1059] = 55;
    exp_40_ram[1060] = 137;
    exp_40_ram[1061] = 9;
    exp_40_ram[1062] = 4;
    exp_40_ram[1063] = 240;
    exp_40_ram[1064] = 39;
    exp_40_ram[1065] = 38;
    exp_40_ram[1066] = 36;
    exp_40_ram[1067] = 23;
    exp_40_ram[1068] = 135;
    exp_40_ram[1069] = 151;
    exp_40_ram[1070] = 135;
    exp_40_ram[1071] = 23;
    exp_40_ram[1072] = 7;
    exp_40_ram[1073] = 151;
    exp_40_ram[1074] = 23;
    exp_40_ram[1075] = 37;
    exp_40_ram[1076] = 86;
    exp_40_ram[1077] = 214;
    exp_40_ram[1078] = 135;
    exp_40_ram[1079] = 134;
    exp_40_ram[1080] = 55;
    exp_40_ram[1081] = 135;
    exp_40_ram[1082] = 85;
    exp_40_ram[1083] = 214;
    exp_40_ram[1084] = 4;
    exp_40_ram[1085] = 183;
    exp_40_ram[1086] = 135;
    exp_40_ram[1087] = 133;
    exp_40_ram[1088] = 5;
    exp_40_ram[1089] = 4;
    exp_40_ram[1090] = 240;
    exp_40_ram[1091] = 133;
    exp_40_ram[1092] = 87;
    exp_40_ram[1093] = 180;
    exp_40_ram[1094] = 7;
    exp_40_ram[1095] = 133;
    exp_40_ram[1096] = 132;
    exp_40_ram[1097] = 4;
    exp_40_ram[1098] = 53;
    exp_40_ram[1099] = 32;
    exp_40_ram[1100] = 133;
    exp_40_ram[1101] = 36;
    exp_40_ram[1102] = 36;
    exp_40_ram[1103] = 41;
    exp_40_ram[1104] = 41;
    exp_40_ram[1105] = 42;
    exp_40_ram[1106] = 42;
    exp_40_ram[1107] = 43;
    exp_40_ram[1108] = 1;
    exp_40_ram[1109] = 128;
    exp_40_ram[1110] = 1;
    exp_40_ram[1111] = 38;
    exp_40_ram[1112] = 36;
    exp_40_ram[1113] = 4;
    exp_40_ram[1114] = 240;
    exp_40_ram[1115] = 39;
    exp_40_ram[1116] = 166;
    exp_40_ram[1117] = 6;
    exp_40_ram[1118] = 224;
    exp_40_ram[1119] = 55;
    exp_40_ram[1120] = 167;
    exp_40_ram[1121] = 5;
    exp_40_ram[1122] = 6;
    exp_40_ram[1123] = 32;
    exp_40_ram[1124] = 34;
    exp_40_ram[1125] = 32;
    exp_40_ram[1126] = 36;
    exp_40_ram[1127] = 5;
    exp_40_ram[1128] = 1;
    exp_40_ram[1129] = 128;
    exp_40_ram[1130] = 1;
    exp_40_ram[1131] = 34;
    exp_40_ram[1132] = 4;
    exp_40_ram[1133] = 5;
    exp_40_ram[1134] = 36;
    exp_40_ram[1135] = 38;
    exp_40_ram[1136] = 132;
    exp_40_ram[1137] = 240;
    exp_40_ram[1138] = 133;
    exp_40_ram[1139] = 180;
    exp_40_ram[1140] = 55;
    exp_40_ram[1141] = 4;
    exp_40_ram[1142] = 4;
    exp_40_ram[1143] = 135;
    exp_40_ram[1144] = 32;
    exp_40_ram[1145] = 162;
    exp_40_ram[1146] = 36;
    exp_40_ram[1147] = 160;
    exp_40_ram[1148] = 36;
    exp_40_ram[1149] = 1;
    exp_40_ram[1150] = 128;
    exp_40_ram[1151] = 1;
    exp_40_ram[1152] = 37;
    exp_40_ram[1153] = 34;
    exp_40_ram[1154] = 6;
    exp_40_ram[1155] = 4;
    exp_40_ram[1156] = 133;
    exp_40_ram[1157] = 5;
    exp_40_ram[1158] = 38;
    exp_40_ram[1159] = 36;
    exp_40_ram[1160] = 32;
    exp_40_ram[1161] = 46;
    exp_40_ram[1162] = 44;
    exp_40_ram[1163] = 240;
    exp_40_ram[1164] = 37;
    exp_40_ram[1165] = 6;
    exp_40_ram[1166] = 133;
    exp_40_ram[1167] = 5;
    exp_40_ram[1168] = 240;
    exp_40_ram[1169] = 167;
    exp_40_ram[1170] = 57;
    exp_40_ram[1171] = 132;
    exp_40_ram[1172] = 149;
    exp_40_ram[1173] = 133;
    exp_40_ram[1174] = 7;
    exp_40_ram[1175] = 9;
    exp_40_ram[1176] = 133;
    exp_40_ram[1177] = 6;
    exp_40_ram[1178] = 133;
    exp_40_ram[1179] = 240;
    exp_40_ram[1180] = 1;
    exp_40_ram[1181] = 167;
    exp_40_ram[1182] = 6;
    exp_40_ram[1183] = 5;
    exp_40_ram[1184] = 149;
    exp_40_ram[1185] = 133;
    exp_40_ram[1186] = 7;
    exp_40_ram[1187] = 133;
    exp_40_ram[1188] = 240;
    exp_40_ram[1189] = 3;
    exp_40_ram[1190] = 165;
    exp_40_ram[1191] = 5;
    exp_40_ram[1192] = 10;
    exp_40_ram[1193] = 16;
    exp_40_ram[1194] = 36;
    exp_40_ram[1195] = 39;
    exp_40_ram[1196] = 38;
    exp_40_ram[1197] = 5;
    exp_40_ram[1198] = 135;
    exp_40_ram[1199] = 4;
    exp_40_ram[1200] = 39;
    exp_40_ram[1201] = 5;
    exp_40_ram[1202] = 135;
    exp_40_ram[1203] = 4;
    exp_40_ram[1204] = 165;
    exp_40_ram[1205] = 16;
    exp_40_ram[1206] = 36;
    exp_40_ram[1207] = 39;
    exp_40_ram[1208] = 38;
    exp_40_ram[1209] = 6;
    exp_40_ram[1210] = 135;
    exp_40_ram[1211] = 5;
    exp_40_ram[1212] = 39;
    exp_40_ram[1213] = 5;
    exp_40_ram[1214] = 135;
    exp_40_ram[1215] = 6;
    exp_40_ram[1216] = 165;
    exp_40_ram[1217] = 16;
    exp_40_ram[1218] = 36;
    exp_40_ram[1219] = 39;
    exp_40_ram[1220] = 38;
    exp_40_ram[1221] = 8;
    exp_40_ram[1222] = 135;
    exp_40_ram[1223] = 7;
    exp_40_ram[1224] = 39;
    exp_40_ram[1225] = 5;
    exp_40_ram[1226] = 135;
    exp_40_ram[1227] = 7;
    exp_40_ram[1228] = 165;
    exp_40_ram[1229] = 16;
    exp_40_ram[1230] = 36;
    exp_40_ram[1231] = 39;
    exp_40_ram[1232] = 38;
    exp_40_ram[1233] = 9;
    exp_40_ram[1234] = 135;
    exp_40_ram[1235] = 8;
    exp_40_ram[1236] = 39;
    exp_40_ram[1237] = 5;
    exp_40_ram[1238] = 135;
    exp_40_ram[1239] = 9;
    exp_40_ram[1240] = 165;
    exp_40_ram[1241] = 5;
    exp_40_ram[1242] = 16;
    exp_40_ram[1243] = 36;
    exp_40_ram[1244] = 38;
    exp_40_ram[1245] = 39;
    exp_40_ram[1246] = 37;
    exp_40_ram[1247] = 5;
    exp_40_ram[1248] = 135;
    exp_40_ram[1249] = 10;
    exp_40_ram[1250] = 16;
    exp_40_ram[1251] = 36;
    exp_40_ram[1252] = 38;
    exp_40_ram[1253] = 39;
    exp_40_ram[1254] = 37;
    exp_40_ram[1255] = 5;
    exp_40_ram[1256] = 135;
    exp_40_ram[1257] = 10;
    exp_40_ram[1258] = 0;
    exp_40_ram[1259] = 36;
    exp_40_ram[1260] = 39;
    exp_40_ram[1261] = 38;
    exp_40_ram[1262] = 32;
    exp_40_ram[1263] = 135;
    exp_40_ram[1264] = 11;
    exp_40_ram[1265] = 39;
    exp_40_ram[1266] = 36;
    exp_40_ram[1267] = 41;
    exp_40_ram[1268] = 135;
    exp_40_ram[1269] = 11;
    exp_40_ram[1270] = 7;
    exp_40_ram[1271] = 28;
    exp_40_ram[1272] = 36;
    exp_40_ram[1273] = 42;
    exp_40_ram[1274] = 133;
    exp_40_ram[1275] = 41;
    exp_40_ram[1276] = 1;
    exp_40_ram[1277] = 128;
    exp_40_ram[1278] = 1;
    exp_40_ram[1279] = 36;
    exp_40_ram[1280] = 90;
    exp_40_ram[1281] = 44;
    exp_40_ram[1282] = 42;
    exp_40_ram[1283] = 40;
    exp_40_ram[1284] = 38;
    exp_40_ram[1285] = 34;
    exp_40_ram[1286] = 46;
    exp_40_ram[1287] = 32;
    exp_40_ram[1288] = 46;
    exp_40_ram[1289] = 44;
    exp_40_ram[1290] = 42;
    exp_40_ram[1291] = 4;
    exp_40_ram[1292] = 132;
    exp_40_ram[1293] = 9;
    exp_40_ram[1294] = 9;
    exp_40_ram[1295] = 10;
    exp_40_ram[1296] = 10;
    exp_40_ram[1297] = 133;
    exp_40_ram[1298] = 240;
    exp_40_ram[1299] = 53;
    exp_40_ram[1300] = 5;
    exp_40_ram[1301] = 5;
    exp_40_ram[1302] = 240;
    exp_40_ram[1303] = 135;
    exp_40_ram[1304] = 20;
    exp_40_ram[1305] = 224;
    exp_40_ram[1306] = 138;
    exp_40_ram[1307] = 133;
    exp_40_ram[1308] = 183;
    exp_40_ram[1309] = 9;
    exp_40_ram[1310] = 4;
    exp_40_ram[1311] = 137;
    exp_40_ram[1312] = 240;
    exp_40_ram[1313] = 92;
    exp_40_ram[1314] = 12;
    exp_40_ram[1315] = 10;
    exp_40_ram[1316] = 12;
    exp_40_ram[1317] = 133;
    exp_40_ram[1318] = 133;
    exp_40_ram[1319] = 240;
    exp_40_ram[1320] = 5;
    exp_40_ram[1321] = 139;
    exp_40_ram[1322] = 11;
    exp_40_ram[1323] = 140;
    exp_40_ram[1324] = 240;
    exp_40_ram[1325] = 20;
    exp_40_ram[1326] = 224;
    exp_40_ram[1327] = 133;
    exp_40_ram[1328] = 183;
    exp_40_ram[1329] = 138;
    exp_40_ram[1330] = 10;
    exp_40_ram[1331] = 4;
    exp_40_ram[1332] = 9;
    exp_40_ram[1333] = 240;
    exp_40_ram[1334] = 85;
    exp_40_ram[1335] = 133;
    exp_40_ram[1336] = 133;
    exp_40_ram[1337] = 0;
    exp_40_ram[1338] = 38;
    exp_40_ram[1339] = 4;
    exp_40_ram[1340] = 36;
    exp_40_ram[1341] = 10;
    exp_40_ram[1342] = 37;
    exp_40_ram[1343] = 21;
    exp_40_ram[1344] = 133;
    exp_40_ram[1345] = 0;
    exp_40_ram[1346] = 38;
    exp_40_ram[1347] = 9;
    exp_40_ram[1348] = 36;
    exp_40_ram[1349] = 37;
    exp_40_ram[1350] = 5;
    exp_40_ram[1351] = 137;
    exp_40_ram[1352] = 0;
    exp_40_ram[1353] = 135;
    exp_40_ram[1354] = 36;
    exp_40_ram[1355] = 38;
    exp_40_ram[1356] = 32;
    exp_40_ram[1357] = 34;
    exp_40_ram[1358] = 36;
    exp_40_ram[1359] = 40;
    exp_40_ram[1360] = 42;
    exp_40_ram[1361] = 133;
    exp_40_ram[1362] = 38;
    exp_40_ram[1363] = 5;
    exp_40_ram[1364] = 240;
    exp_40_ram[1365] = 44;
    exp_40_ram[1366] = 46;
    exp_40_ram[1367] = 32;
    exp_40_ram[1368] = 5;
    exp_40_ram[1369] = 36;
    exp_40_ram[1370] = 36;
    exp_40_ram[1371] = 41;
    exp_40_ram[1372] = 41;
    exp_40_ram[1373] = 42;
    exp_40_ram[1374] = 42;
    exp_40_ram[1375] = 43;
    exp_40_ram[1376] = 43;
    exp_40_ram[1377] = 44;
    exp_40_ram[1378] = 44;
    exp_40_ram[1379] = 1;
    exp_40_ram[1380] = 128;
    exp_40_ram[1381] = 1;
    exp_40_ram[1382] = 32;
    exp_40_ram[1383] = 43;
    exp_40_ram[1384] = 6;
    exp_40_ram[1385] = 42;
    exp_40_ram[1386] = 40;
    exp_40_ram[1387] = 4;
    exp_40_ram[1388] = 36;
    exp_40_ram[1389] = 34;
    exp_40_ram[1390] = 10;
    exp_40_ram[1391] = 9;
    exp_40_ram[1392] = 10;
    exp_40_ram[1393] = 5;
    exp_40_ram[1394] = 5;
    exp_40_ram[1395] = 46;
    exp_40_ram[1396] = 44;
    exp_40_ram[1397] = 38;
    exp_40_ram[1398] = 32;
    exp_40_ram[1399] = 34;
    exp_40_ram[1400] = 38;
    exp_40_ram[1401] = 36;
    exp_40_ram[1402] = 46;
    exp_40_ram[1403] = 44;
    exp_40_ram[1404] = 44;
    exp_40_ram[1405] = 240;
    exp_40_ram[1406] = 5;
    exp_40_ram[1407] = 240;
    exp_40_ram[1408] = 134;
    exp_40_ram[1409] = 5;
    exp_40_ram[1410] = 5;
    exp_40_ram[1411] = 240;
    exp_40_ram[1412] = 39;
    exp_40_ram[1413] = 39;
    exp_40_ram[1414] = 6;
    exp_40_ram[1415] = 5;
    exp_40_ram[1416] = 135;
    exp_40_ram[1417] = 5;
    exp_40_ram[1418] = 34;
    exp_40_ram[1419] = 240;
    exp_40_ram[1420] = 5;
    exp_40_ram[1421] = 240;
    exp_40_ram[1422] = 6;
    exp_40_ram[1423] = 9;
    exp_40_ram[1424] = 132;
    exp_40_ram[1425] = 5;
    exp_40_ram[1426] = 5;
    exp_40_ram[1427] = 34;
    exp_40_ram[1428] = 36;
    exp_40_ram[1429] = 40;
    exp_40_ram[1430] = 38;
    exp_40_ram[1431] = 32;
    exp_40_ram[1432] = 46;
    exp_40_ram[1433] = 240;
    exp_40_ram[1434] = 5;
    exp_40_ram[1435] = 240;
    exp_40_ram[1436] = 134;
    exp_40_ram[1437] = 5;
    exp_40_ram[1438] = 5;
    exp_40_ram[1439] = 240;
    exp_40_ram[1440] = 6;
    exp_40_ram[1441] = 5;
    exp_40_ram[1442] = 5;
    exp_40_ram[1443] = 36;
    exp_40_ram[1444] = 240;
    exp_40_ram[1445] = 5;
    exp_40_ram[1446] = 240;
    exp_40_ram[1447] = 6;
    exp_40_ram[1448] = 10;
    exp_40_ram[1449] = 132;
    exp_40_ram[1450] = 5;
    exp_40_ram[1451] = 5;
    exp_40_ram[1452] = 240;
    exp_40_ram[1453] = 5;
    exp_40_ram[1454] = 240;
    exp_40_ram[1455] = 7;
    exp_40_ram[1456] = 135;
    exp_40_ram[1457] = 230;
    exp_40_ram[1458] = 156;
    exp_40_ram[1459] = 122;
    exp_40_ram[1460] = 5;
    exp_40_ram[1461] = 232;
    exp_40_ram[1462] = 20;
    exp_40_ram[1463] = 100;
    exp_40_ram[1464] = 5;
    exp_40_ram[1465] = 32;
    exp_40_ram[1466] = 36;
    exp_40_ram[1467] = 36;
    exp_40_ram[1468] = 41;
    exp_40_ram[1469] = 41;
    exp_40_ram[1470] = 42;
    exp_40_ram[1471] = 42;
    exp_40_ram[1472] = 43;
    exp_40_ram[1473] = 1;
    exp_40_ram[1474] = 128;
    exp_40_ram[1475] = 1;
    exp_40_ram[1476] = 5;
    exp_40_ram[1477] = 40;
    exp_40_ram[1478] = 6;
    exp_40_ram[1479] = 9;
    exp_40_ram[1480] = 5;
    exp_40_ram[1481] = 46;
    exp_40_ram[1482] = 44;
    exp_40_ram[1483] = 42;
    exp_40_ram[1484] = 38;
    exp_40_ram[1485] = 240;
    exp_40_ram[1486] = 6;
    exp_40_ram[1487] = 5;
    exp_40_ram[1488] = 5;
    exp_40_ram[1489] = 41;
    exp_40_ram[1490] = 240;
    exp_40_ram[1491] = 5;
    exp_40_ram[1492] = 240;
    exp_40_ram[1493] = 4;
    exp_40_ram[1494] = 132;
    exp_40_ram[1495] = 86;
    exp_40_ram[1496] = 23;
    exp_40_ram[1497] = 135;
    exp_40_ram[1498] = 7;
    exp_40_ram[1499] = 183;
    exp_40_ram[1500] = 132;
    exp_40_ram[1501] = 4;
    exp_40_ram[1502] = 5;
    exp_40_ram[1503] = 134;
    exp_40_ram[1504] = 5;
    exp_40_ram[1505] = 240;
    exp_40_ram[1506] = 6;
    exp_40_ram[1507] = 5;
    exp_40_ram[1508] = 5;
    exp_40_ram[1509] = 240;
    exp_40_ram[1510] = 94;
    exp_40_ram[1511] = 7;
    exp_40_ram[1512] = 32;
    exp_40_ram[1513] = 32;
    exp_40_ram[1514] = 5;
    exp_40_ram[1515] = 36;
    exp_40_ram[1516] = 41;
    exp_40_ram[1517] = 41;
    exp_40_ram[1518] = 133;
    exp_40_ram[1519] = 36;
    exp_40_ram[1520] = 1;
    exp_40_ram[1521] = 128;
    exp_40_ram[1522] = 136;
    exp_40_ram[1523] = 5;
    exp_40_ram[1524] = 6;
    exp_40_ram[1525] = 5;
    exp_40_ram[1526] = 240;
    exp_40_ram[1527] = 5;
    exp_40_ram[1528] = 240;
    exp_40_ram[1529] = 85;
    exp_40_ram[1530] = 5;
    exp_40_ram[1531] = 55;
    exp_40_ram[1532] = 132;
    exp_40_ram[1533] = 132;
    exp_40_ram[1534] = 103;
    exp_40_ram[1535] = 4;
    exp_40_ram[1536] = 140;
    exp_40_ram[1537] = 20;
    exp_40_ram[1538] = 4;
    exp_40_ram[1539] = 4;
    exp_40_ram[1540] = 240;
    exp_40_ram[1541] = 136;
    exp_40_ram[1542] = 6;
    exp_40_ram[1543] = 5;
    exp_40_ram[1544] = 5;
    exp_40_ram[1545] = 240;
    exp_40_ram[1546] = 5;
    exp_40_ram[1547] = 240;
    exp_40_ram[1548] = 6;
    exp_40_ram[1549] = 21;
    exp_40_ram[1550] = 5;
    exp_40_ram[1551] = 32;
    exp_40_ram[1552] = 240;
    exp_40_ram[1553] = 32;
    exp_40_ram[1554] = 240;
    exp_40_ram[1555] = 1;
    exp_40_ram[1556] = 134;
    exp_40_ram[1557] = 5;
    exp_40_ram[1558] = 5;
    exp_40_ram[1559] = 38;
    exp_40_ram[1560] = 240;
    exp_40_ram[1561] = 5;
    exp_40_ram[1562] = 6;
    exp_40_ram[1563] = 5;
    exp_40_ram[1564] = 240;
    exp_40_ram[1565] = 5;
    exp_40_ram[1566] = 240;
    exp_40_ram[1567] = 32;
    exp_40_ram[1568] = 1;
    exp_40_ram[1569] = 128;
    exp_40_ram[1570] = 1;
    exp_40_ram[1571] = 34;
    exp_40_ram[1572] = 32;
    exp_40_ram[1573] = 36;
    exp_40_ram[1574] = 41;
    exp_40_ram[1575] = 38;
    exp_40_ram[1576] = 133;
    exp_40_ram[1577] = 5;
    exp_40_ram[1578] = 36;
    exp_40_ram[1579] = 46;
    exp_40_ram[1580] = 240;
    exp_40_ram[1581] = 6;
    exp_40_ram[1582] = 6;
    exp_40_ram[1583] = 22;
    exp_40_ram[1584] = 6;
    exp_40_ram[1585] = 5;
    exp_40_ram[1586] = 182;
    exp_40_ram[1587] = 6;
    exp_40_ram[1588] = 5;
    exp_40_ram[1589] = 240;
    exp_40_ram[1590] = 52;
    exp_40_ram[1591] = 5;
    exp_40_ram[1592] = 6;
    exp_40_ram[1593] = 5;
    exp_40_ram[1594] = 240;
    exp_40_ram[1595] = 5;
    exp_40_ram[1596] = 133;
    exp_40_ram[1597] = 240;
    exp_40_ram[1598] = 9;
    exp_40_ram[1599] = 160;
    exp_40_ram[1600] = 32;
    exp_40_ram[1601] = 5;
    exp_40_ram[1602] = 36;
    exp_40_ram[1603] = 36;
    exp_40_ram[1604] = 41;
    exp_40_ram[1605] = 41;
    exp_40_ram[1606] = 1;
    exp_40_ram[1607] = 128;
    exp_40_ram[1608] = 1;
    exp_40_ram[1609] = 38;
    exp_40_ram[1610] = 36;
    exp_40_ram[1611] = 34;
    exp_40_ram[1612] = 32;
    exp_40_ram[1613] = 4;
    exp_40_ram[1614] = 46;
    exp_40_ram[1615] = 240;
    exp_40_ram[1616] = 36;
    exp_40_ram[1617] = 38;
    exp_40_ram[1618] = 0;
    exp_40_ram[1619] = 240;
    exp_40_ram[1620] = 6;
    exp_40_ram[1621] = 134;
    exp_40_ram[1622] = 37;
    exp_40_ram[1623] = 37;
    exp_40_ram[1624] = 7;
    exp_40_ram[1625] = 8;
    exp_40_ram[1626] = 56;
    exp_40_ram[1627] = 135;
    exp_40_ram[1628] = 134;
    exp_40_ram[1629] = 135;
    exp_40_ram[1630] = 38;
    exp_40_ram[1631] = 137;
    exp_40_ram[1632] = 9;
    exp_40_ram[1633] = 134;
    exp_40_ram[1634] = 134;
    exp_40_ram[1635] = 224;
    exp_40_ram[1636] = 134;
    exp_40_ram[1637] = 134;
    exp_40_ram[1638] = 24;
    exp_40_ram[1639] = 6;
    exp_40_ram[1640] = 7;
    exp_40_ram[1641] = 228;
    exp_40_ram[1642] = 0;
    exp_40_ram[1643] = 133;
    exp_40_ram[1644] = 32;
    exp_40_ram[1645] = 36;
    exp_40_ram[1646] = 41;
    exp_40_ram[1647] = 41;
    exp_40_ram[1648] = 1;
    exp_40_ram[1649] = 128;
    exp_40_ram[1650] = 1;
    exp_40_ram[1651] = 38;
    exp_40_ram[1652] = 36;
    exp_40_ram[1653] = 4;
    exp_40_ram[1654] = 5;
    exp_40_ram[1655] = 224;
    exp_40_ram[1656] = 0;
    exp_40_ram[1657] = 32;
    exp_40_ram[1658] = 36;
    exp_40_ram[1659] = 1;
    exp_40_ram[1660] = 128;
    exp_40_ram[1661] = 1;
    exp_40_ram[1662] = 46;
    exp_40_ram[1663] = 44;
    exp_40_ram[1664] = 4;
    exp_40_ram[1665] = 5;
    exp_40_ram[1666] = 224;
    exp_40_ram[1667] = 7;
    exp_40_ram[1668] = 38;
    exp_40_ram[1669] = 36;
    exp_40_ram[1670] = 0;
    exp_40_ram[1671] = 37;
    exp_40_ram[1672] = 5;
    exp_40_ram[1673] = 240;
    exp_40_ram[1674] = 0;
    exp_40_ram[1675] = 39;
    exp_40_ram[1676] = 151;
    exp_40_ram[1677] = 38;
    exp_40_ram[1678] = 39;
    exp_40_ram[1679] = 167;
    exp_40_ram[1680] = 133;
    exp_40_ram[1681] = 37;
    exp_40_ram[1682] = 224;
    exp_40_ram[1683] = 39;
    exp_40_ram[1684] = 167;
    exp_40_ram[1685] = 7;
    exp_40_ram[1686] = 87;
    exp_40_ram[1687] = 133;
    exp_40_ram[1688] = 240;
    exp_40_ram[1689] = 39;
    exp_40_ram[1690] = 7;
    exp_40_ram[1691] = 208;
    exp_40_ram[1692] = 0;
    exp_40_ram[1693] = 39;
    exp_40_ram[1694] = 215;
    exp_40_ram[1695] = 38;
    exp_40_ram[1696] = 39;
    exp_40_ram[1697] = 167;
    exp_40_ram[1698] = 133;
    exp_40_ram[1699] = 37;
    exp_40_ram[1700] = 224;
    exp_40_ram[1701] = 39;
    exp_40_ram[1702] = 167;
    exp_40_ram[1703] = 7;
    exp_40_ram[1704] = 87;
    exp_40_ram[1705] = 133;
    exp_40_ram[1706] = 240;
    exp_40_ram[1707] = 39;
    exp_40_ram[1708] = 7;
    exp_40_ram[1709] = 192;
    exp_40_ram[1710] = 39;
    exp_40_ram[1711] = 135;
    exp_40_ram[1712] = 36;
    exp_40_ram[1713] = 39;
    exp_40_ram[1714] = 7;
    exp_40_ram[1715] = 216;
    exp_40_ram[1716] = 39;
    exp_40_ram[1717] = 167;
    exp_40_ram[1718] = 133;
    exp_40_ram[1719] = 5;
    exp_40_ram[1720] = 224;
    exp_40_ram[1721] = 0;
    exp_40_ram[1722] = 32;
    exp_40_ram[1723] = 36;
    exp_40_ram[1724] = 1;
    exp_40_ram[1725] = 128;
    exp_40_ram[1726] = 1;
    exp_40_ram[1727] = 46;
    exp_40_ram[1728] = 44;
    exp_40_ram[1729] = 4;
    exp_40_ram[1730] = 39;
    exp_40_ram[1731] = 7;
    exp_40_ram[1732] = 170;
    exp_40_ram[1733] = 39;
    exp_40_ram[1734] = 7;
    exp_40_ram[1735] = 168;
    exp_40_ram[1736] = 39;
    exp_40_ram[1737] = 7;
    exp_40_ram[1738] = 166;
    exp_40_ram[1739] = 39;
    exp_40_ram[1740] = 7;
    exp_40_ram[1741] = 164;
    exp_40_ram[1742] = 39;
    exp_40_ram[1743] = 7;
    exp_40_ram[1744] = 162;
    exp_40_ram[1745] = 39;
    exp_40_ram[1746] = 160;
    exp_40_ram[1747] = 39;
    exp_40_ram[1748] = 7;
    exp_40_ram[1749] = 160;
    exp_40_ram[1750] = 37;
    exp_40_ram[1751] = 240;
    exp_40_ram[1752] = 7;
    exp_40_ram[1753] = 135;
    exp_40_ram[1754] = 5;
    exp_40_ram[1755] = 133;
    exp_40_ram[1756] = 240;
    exp_40_ram[1757] = 5;
    exp_40_ram[1758] = 240;
    exp_40_ram[1759] = 7;
    exp_40_ram[1760] = 135;
    exp_40_ram[1761] = 32;
    exp_40_ram[1762] = 34;
    exp_40_ram[1763] = 7;
    exp_40_ram[1764] = 133;
    exp_40_ram[1765] = 240;
    exp_40_ram[1766] = 38;
    exp_40_ram[1767] = 37;
    exp_40_ram[1768] = 240;
    exp_40_ram[1769] = 7;
    exp_40_ram[1770] = 133;
    exp_40_ram[1771] = 224;
    exp_40_ram[1772] = 39;
    exp_40_ram[1773] = 167;
    exp_40_ram[1774] = 133;
    exp_40_ram[1775] = 240;
    exp_40_ram[1776] = 240;
    exp_40_ram[1777] = 1;
    exp_40_ram[1778] = 38;
    exp_40_ram[1779] = 36;
    exp_40_ram[1780] = 34;
    exp_40_ram[1781] = 32;
    exp_40_ram[1782] = 46;
    exp_40_ram[1783] = 44;
    exp_40_ram[1784] = 42;
    exp_40_ram[1785] = 40;
    exp_40_ram[1786] = 38;
    exp_40_ram[1787] = 36;
    exp_40_ram[1788] = 34;
    exp_40_ram[1789] = 32;
    exp_40_ram[1790] = 4;
    exp_40_ram[1791] = 7;
    exp_40_ram[1792] = 46;
    exp_40_ram[1793] = 7;
    exp_40_ram[1794] = 7;
    exp_40_ram[1795] = 40;
    exp_40_ram[1796] = 42;
    exp_40_ram[1797] = 240;
    exp_40_ram[1798] = 32;
    exp_40_ram[1799] = 34;
    exp_40_ram[1800] = 38;
    exp_40_ram[1801] = 0;
    exp_40_ram[1802] = 39;
    exp_40_ram[1803] = 87;
    exp_40_ram[1804] = 135;
    exp_40_ram[1805] = 7;
    exp_40_ram[1806] = 46;
    exp_40_ram[1807] = 39;
    exp_40_ram[1808] = 87;
    exp_40_ram[1809] = 135;
    exp_40_ram[1810] = 7;
    exp_40_ram[1811] = 46;
    exp_40_ram[1812] = 39;
    exp_40_ram[1813] = 87;
    exp_40_ram[1814] = 135;
    exp_40_ram[1815] = 7;
    exp_40_ram[1816] = 46;
    exp_40_ram[1817] = 39;
    exp_40_ram[1818] = 87;
    exp_40_ram[1819] = 135;
    exp_40_ram[1820] = 7;
    exp_40_ram[1821] = 46;
    exp_40_ram[1822] = 39;
    exp_40_ram[1823] = 135;
    exp_40_ram[1824] = 38;
    exp_40_ram[1825] = 240;
    exp_40_ram[1826] = 6;
    exp_40_ram[1827] = 134;
    exp_40_ram[1828] = 37;
    exp_40_ram[1829] = 37;
    exp_40_ram[1830] = 7;
    exp_40_ram[1831] = 8;
    exp_40_ram[1832] = 56;
    exp_40_ram[1833] = 135;
    exp_40_ram[1834] = 134;
    exp_40_ram[1835] = 135;
    exp_40_ram[1836] = 38;
    exp_40_ram[1837] = 166;
    exp_40_ram[1838] = 36;
    exp_40_ram[1839] = 38;
    exp_40_ram[1840] = 37;
    exp_40_ram[1841] = 37;
    exp_40_ram[1842] = 134;
    exp_40_ram[1843] = 134;
    exp_40_ram[1844] = 236;
    exp_40_ram[1845] = 134;
    exp_40_ram[1846] = 134;
    exp_40_ram[1847] = 24;
    exp_40_ram[1848] = 6;
    exp_40_ram[1849] = 7;
    exp_40_ram[1850] = 224;
    exp_40_ram[1851] = 37;
    exp_40_ram[1852] = 5;
    exp_40_ram[1853] = 224;
    exp_40_ram[1854] = 240;
    exp_40_ram[1855] = 32;
    exp_40_ram[1856] = 34;
    exp_40_ram[1857] = 38;
    exp_40_ram[1858] = 0;
    exp_40_ram[1859] = 39;
    exp_40_ram[1860] = 39;
    exp_40_ram[1861] = 86;
    exp_40_ram[1862] = 134;
    exp_40_ram[1863] = 134;
    exp_40_ram[1864] = 6;
    exp_40_ram[1865] = 6;
    exp_40_ram[1866] = 6;
    exp_40_ram[1867] = 86;
    exp_40_ram[1868] = 134;
    exp_40_ram[1869] = 5;
    exp_40_ram[1870] = 57;
    exp_40_ram[1871] = 137;
    exp_40_ram[1872] = 7;
    exp_40_ram[1873] = 137;
    exp_40_ram[1874] = 40;
    exp_40_ram[1875] = 42;
    exp_40_ram[1876] = 39;
    exp_40_ram[1877] = 39;
    exp_40_ram[1878] = 86;
    exp_40_ram[1879] = 134;
    exp_40_ram[1880] = 134;
    exp_40_ram[1881] = 6;
    exp_40_ram[1882] = 6;
    exp_40_ram[1883] = 6;
    exp_40_ram[1884] = 86;
    exp_40_ram[1885] = 134;
    exp_40_ram[1886] = 5;
    exp_40_ram[1887] = 58;
    exp_40_ram[1888] = 138;
    exp_40_ram[1889] = 7;
    exp_40_ram[1890] = 138;
    exp_40_ram[1891] = 40;
    exp_40_ram[1892] = 42;
    exp_40_ram[1893] = 39;
    exp_40_ram[1894] = 39;
    exp_40_ram[1895] = 86;
    exp_40_ram[1896] = 134;
    exp_40_ram[1897] = 134;
    exp_40_ram[1898] = 6;
    exp_40_ram[1899] = 6;
    exp_40_ram[1900] = 6;
    exp_40_ram[1901] = 86;
    exp_40_ram[1902] = 134;
    exp_40_ram[1903] = 5;
    exp_40_ram[1904] = 59;
    exp_40_ram[1905] = 139;
    exp_40_ram[1906] = 7;
    exp_40_ram[1907] = 139;
    exp_40_ram[1908] = 40;
    exp_40_ram[1909] = 42;
    exp_40_ram[1910] = 39;
    exp_40_ram[1911] = 39;
    exp_40_ram[1912] = 86;
    exp_40_ram[1913] = 134;
    exp_40_ram[1914] = 134;
    exp_40_ram[1915] = 6;
    exp_40_ram[1916] = 6;
    exp_40_ram[1917] = 6;
    exp_40_ram[1918] = 86;
    exp_40_ram[1919] = 134;
    exp_40_ram[1920] = 5;
    exp_40_ram[1921] = 60;
    exp_40_ram[1922] = 140;
    exp_40_ram[1923] = 7;
    exp_40_ram[1924] = 140;
    exp_40_ram[1925] = 40;
    exp_40_ram[1926] = 42;
    exp_40_ram[1927] = 39;
    exp_40_ram[1928] = 135;
    exp_40_ram[1929] = 38;
    exp_40_ram[1930] = 240;
    exp_40_ram[1931] = 6;
    exp_40_ram[1932] = 134;
    exp_40_ram[1933] = 37;
    exp_40_ram[1934] = 37;
    exp_40_ram[1935] = 7;
    exp_40_ram[1936] = 8;
    exp_40_ram[1937] = 56;
    exp_40_ram[1938] = 135;
    exp_40_ram[1939] = 134;
    exp_40_ram[1940] = 135;
    exp_40_ram[1941] = 38;
    exp_40_ram[1942] = 166;
    exp_40_ram[1943] = 32;
    exp_40_ram[1944] = 34;
    exp_40_ram[1945] = 37;
    exp_40_ram[1946] = 37;
    exp_40_ram[1947] = 134;
    exp_40_ram[1948] = 134;
    exp_40_ram[1949] = 236;
    exp_40_ram[1950] = 134;
    exp_40_ram[1951] = 134;
    exp_40_ram[1952] = 24;
    exp_40_ram[1953] = 6;
    exp_40_ram[1954] = 7;
    exp_40_ram[1955] = 224;
    exp_40_ram[1956] = 37;
    exp_40_ram[1957] = 5;
    exp_40_ram[1958] = 224;
    exp_40_ram[1959] = 240;
    exp_40_ram[1960] = 32;
    exp_40_ram[1961] = 34;
    exp_40_ram[1962] = 38;
    exp_40_ram[1963] = 0;
    exp_40_ram[1964] = 39;
    exp_40_ram[1965] = 87;
    exp_40_ram[1966] = 135;
    exp_40_ram[1967] = 87;
    exp_40_ram[1968] = 46;
    exp_40_ram[1969] = 39;
    exp_40_ram[1970] = 87;
    exp_40_ram[1971] = 135;
    exp_40_ram[1972] = 87;
    exp_40_ram[1973] = 46;
    exp_40_ram[1974] = 39;
    exp_40_ram[1975] = 87;
    exp_40_ram[1976] = 135;
    exp_40_ram[1977] = 87;
    exp_40_ram[1978] = 46;
    exp_40_ram[1979] = 39;
    exp_40_ram[1980] = 87;
    exp_40_ram[1981] = 135;
    exp_40_ram[1982] = 87;
    exp_40_ram[1983] = 46;
    exp_40_ram[1984] = 39;
    exp_40_ram[1985] = 135;
    exp_40_ram[1986] = 38;
    exp_40_ram[1987] = 240;
    exp_40_ram[1988] = 6;
    exp_40_ram[1989] = 134;
    exp_40_ram[1990] = 37;
    exp_40_ram[1991] = 37;
    exp_40_ram[1992] = 7;
    exp_40_ram[1993] = 8;
    exp_40_ram[1994] = 56;
    exp_40_ram[1995] = 135;
    exp_40_ram[1996] = 134;
    exp_40_ram[1997] = 135;
    exp_40_ram[1998] = 38;
    exp_40_ram[1999] = 166;
    exp_40_ram[2000] = 44;
    exp_40_ram[2001] = 46;
    exp_40_ram[2002] = 37;
    exp_40_ram[2003] = 37;
    exp_40_ram[2004] = 134;
    exp_40_ram[2005] = 134;
    exp_40_ram[2006] = 236;
    exp_40_ram[2007] = 134;
    exp_40_ram[2008] = 134;
    exp_40_ram[2009] = 24;
    exp_40_ram[2010] = 6;
    exp_40_ram[2011] = 7;
    exp_40_ram[2012] = 224;
    exp_40_ram[2013] = 37;
    exp_40_ram[2014] = 5;
    exp_40_ram[2015] = 224;
    exp_40_ram[2016] = 240;
    exp_40_ram[2017] = 32;
    exp_40_ram[2018] = 34;
    exp_40_ram[2019] = 38;
    exp_40_ram[2020] = 0;
    exp_40_ram[2021] = 39;
    exp_40_ram[2022] = 39;
    exp_40_ram[2023] = 86;
    exp_40_ram[2024] = 6;
    exp_40_ram[2025] = 6;
    exp_40_ram[2026] = 5;
    exp_40_ram[2027] = 133;
    exp_40_ram[2028] = 224;
    exp_40_ram[2029] = 7;
    exp_40_ram[2030] = 135;
    exp_40_ram[2031] = 40;
    exp_40_ram[2032] = 42;
    exp_40_ram[2033] = 39;
    exp_40_ram[2034] = 39;
    exp_40_ram[2035] = 86;
    exp_40_ram[2036] = 6;
    exp_40_ram[2037] = 6;
    exp_40_ram[2038] = 5;
    exp_40_ram[2039] = 133;
    exp_40_ram[2040] = 224;
    exp_40_ram[2041] = 7;
    exp_40_ram[2042] = 135;
    exp_40_ram[2043] = 40;
    exp_40_ram[2044] = 42;
    exp_40_ram[2045] = 39;
    exp_40_ram[2046] = 39;
    exp_40_ram[2047] = 86;
    exp_40_ram[2048] = 6;
    exp_40_ram[2049] = 6;
    exp_40_ram[2050] = 5;
    exp_40_ram[2051] = 133;
    exp_40_ram[2052] = 224;
    exp_40_ram[2053] = 7;
    exp_40_ram[2054] = 135;
    exp_40_ram[2055] = 40;
    exp_40_ram[2056] = 42;
    exp_40_ram[2057] = 39;
    exp_40_ram[2058] = 39;
    exp_40_ram[2059] = 86;
    exp_40_ram[2060] = 6;
    exp_40_ram[2061] = 6;
    exp_40_ram[2062] = 5;
    exp_40_ram[2063] = 133;
    exp_40_ram[2064] = 224;
    exp_40_ram[2065] = 7;
    exp_40_ram[2066] = 135;
    exp_40_ram[2067] = 40;
    exp_40_ram[2068] = 42;
    exp_40_ram[2069] = 39;
    exp_40_ram[2070] = 135;
    exp_40_ram[2071] = 38;
    exp_40_ram[2072] = 224;
    exp_40_ram[2073] = 6;
    exp_40_ram[2074] = 134;
    exp_40_ram[2075] = 37;
    exp_40_ram[2076] = 37;
    exp_40_ram[2077] = 7;
    exp_40_ram[2078] = 8;
    exp_40_ram[2079] = 56;
    exp_40_ram[2080] = 135;
    exp_40_ram[2081] = 134;
    exp_40_ram[2082] = 135;
    exp_40_ram[2083] = 38;
    exp_40_ram[2084] = 166;
    exp_40_ram[2085] = 141;
    exp_40_ram[2086] = 13;
    exp_40_ram[2087] = 134;
    exp_40_ram[2088] = 134;
    exp_40_ram[2089] = 232;
    exp_40_ram[2090] = 134;
    exp_40_ram[2091] = 134;
    exp_40_ram[2092] = 24;
    exp_40_ram[2093] = 6;
    exp_40_ram[2094] = 7;
    exp_40_ram[2095] = 236;
    exp_40_ram[2096] = 37;
    exp_40_ram[2097] = 5;
    exp_40_ram[2098] = 224;
    exp_40_ram[2099] = 0;
    exp_40_ram[2100] = 32;
    exp_40_ram[2101] = 36;
    exp_40_ram[2102] = 41;
    exp_40_ram[2103] = 41;
    exp_40_ram[2104] = 42;
    exp_40_ram[2105] = 42;
    exp_40_ram[2106] = 43;
    exp_40_ram[2107] = 43;
    exp_40_ram[2108] = 44;
    exp_40_ram[2109] = 44;
    exp_40_ram[2110] = 45;
    exp_40_ram[2111] = 45;
    exp_40_ram[2112] = 1;
    exp_40_ram[2113] = 128;
    exp_40_ram[2114] = 1;
    exp_40_ram[2115] = 46;
    exp_40_ram[2116] = 44;
    exp_40_ram[2117] = 4;
    exp_40_ram[2118] = 38;
    exp_40_ram[2119] = 0;
    exp_40_ram[2120] = 39;
    exp_40_ram[2121] = 247;
    exp_40_ram[2122] = 39;
    exp_40_ram[2123] = 6;
    exp_40_ram[2124] = 135;
    exp_40_ram[2125] = 128;
    exp_40_ram[2126] = 39;
    exp_40_ram[2127] = 135;
    exp_40_ram[2128] = 38;
    exp_40_ram[2129] = 39;
    exp_40_ram[2130] = 7;
    exp_40_ram[2131] = 218;
    exp_40_ram[2132] = 36;
    exp_40_ram[2133] = 0;
    exp_40_ram[2134] = 37;
    exp_40_ram[2135] = 5;
    exp_40_ram[2136] = 224;
    exp_40_ram[2137] = 39;
    exp_40_ram[2138] = 7;
    exp_40_ram[2139] = 6;
    exp_40_ram[2140] = 7;
    exp_40_ram[2141] = 39;
    exp_40_ram[2142] = 7;
    exp_40_ram[2143] = 135;
    exp_40_ram[2144] = 7;
    exp_40_ram[2145] = 6;
    exp_40_ram[2146] = 133;
    exp_40_ram[2147] = 133;
    exp_40_ram[2148] = 224;
    exp_40_ram[2149] = 39;
    exp_40_ram[2150] = 34;
    exp_40_ram[2151] = 0;
    exp_40_ram[2152] = 39;
    exp_40_ram[2153] = 7;
    exp_40_ram[2154] = 7;
    exp_40_ram[2155] = 199;
    exp_40_ram[2156] = 135;
    exp_40_ram[2157] = 39;
    exp_40_ram[2158] = 6;
    exp_40_ram[2159] = 135;
    exp_40_ram[2160] = 199;
    exp_40_ram[2161] = 134;
    exp_40_ram[2162] = 39;
    exp_40_ram[2163] = 135;
    exp_40_ram[2164] = 8;
    exp_40_ram[2165] = 5;
    exp_40_ram[2166] = 224;
    exp_40_ram[2167] = 0;
    exp_40_ram[2168] = 39;
    exp_40_ram[2169] = 135;
    exp_40_ram[2170] = 34;
    exp_40_ram[2171] = 39;
    exp_40_ram[2172] = 7;
    exp_40_ram[2173] = 214;
    exp_40_ram[2174] = 5;
    exp_40_ram[2175] = 224;
    exp_40_ram[2176] = 39;
    exp_40_ram[2177] = 135;
    exp_40_ram[2178] = 36;
    exp_40_ram[2179] = 39;
    exp_40_ram[2180] = 7;
    exp_40_ram[2181] = 210;
    exp_40_ram[2182] = 5;
    exp_40_ram[2183] = 224;
    exp_40_ram[2184] = 7;
    exp_40_ram[2185] = 32;
    exp_40_ram[2186] = 5;
    exp_40_ram[2187] = 224;
    exp_40_ram[2188] = 7;
    exp_40_ram[2189] = 46;
    exp_40_ram[2190] = 5;
    exp_40_ram[2191] = 224;
    exp_40_ram[2192] = 7;
    exp_40_ram[2193] = 44;
    exp_40_ram[2194] = 42;
    exp_40_ram[2195] = 0;
    exp_40_ram[2196] = 37;
    exp_40_ram[2197] = 224;
    exp_40_ram[2198] = 5;
    exp_40_ram[2199] = 224;
    exp_40_ram[2200] = 7;
    exp_40_ram[2201] = 32;
    exp_40_ram[2202] = 37;
    exp_40_ram[2203] = 224;
    exp_40_ram[2204] = 5;
    exp_40_ram[2205] = 224;
    exp_40_ram[2206] = 7;
    exp_40_ram[2207] = 46;
    exp_40_ram[2208] = 37;
    exp_40_ram[2209] = 224;
    exp_40_ram[2210] = 5;
    exp_40_ram[2211] = 224;
    exp_40_ram[2212] = 7;
    exp_40_ram[2213] = 44;
    exp_40_ram[2214] = 39;
    exp_40_ram[2215] = 39;
    exp_40_ram[2216] = 38;
    exp_40_ram[2217] = 6;
    exp_40_ram[2218] = 133;
    exp_40_ram[2219] = 5;
    exp_40_ram[2220] = 224;
    exp_40_ram[2221] = 39;
    exp_40_ram[2222] = 135;
    exp_40_ram[2223] = 42;
    exp_40_ram[2224] = 39;
    exp_40_ram[2225] = 7;
    exp_40_ram[2226] = 212;
    exp_40_ram[2227] = 37;
    exp_40_ram[2228] = 224;
    exp_40_ram[2229] = 37;
    exp_40_ram[2230] = 224;
    exp_40_ram[2231] = 37;
    exp_40_ram[2232] = 224;
    exp_40_ram[2233] = 32;
    exp_40_ram[2234] = 36;
    exp_40_ram[2235] = 1;
    exp_40_ram[2236] = 128;
    exp_40_ram[2237] = 1;
    exp_40_ram[2238] = 46;
    exp_40_ram[2239] = 44;
    exp_40_ram[2240] = 4;
    exp_40_ram[2241] = 5;
    exp_40_ram[2242] = 224;
    exp_40_ram[2243] = 5;
    exp_40_ram[2244] = 224;
    exp_40_ram[2245] = 5;
    exp_40_ram[2246] = 224;
    exp_40_ram[2247] = 5;
    exp_40_ram[2248] = 224;
    exp_40_ram[2249] = 5;
    exp_40_ram[2250] = 224;
    exp_40_ram[2251] = 5;
    exp_40_ram[2252] = 224;
    exp_40_ram[2253] = 224;
    exp_40_ram[2254] = 7;
    exp_40_ram[2255] = 7;
    exp_40_ram[2256] = 71;
    exp_40_ram[2257] = 135;
    exp_40_ram[2258] = 7;
    exp_40_ram[2259] = 108;
    exp_40_ram[2260] = 151;
    exp_40_ram[2261] = 39;
    exp_40_ram[2262] = 135;
    exp_40_ram[2263] = 7;
    exp_40_ram[2264] = 167;
    exp_40_ram[2265] = 128;
    exp_40_ram[2266] = 240;
    exp_40_ram[2267] = 0;
    exp_40_ram[2268] = 240;
    exp_40_ram[2269] = 0;
    exp_40_ram[2270] = 240;
    exp_40_ram[2271] = 0;
    exp_40_ram[2272] = 240;
    exp_40_ram[2273] = 0;
    exp_40_ram[2274] = 240;
    exp_40_ram[2275] = 0;
    exp_40_ram[2276] = 240;
    exp_40_ram[2277] = 7;
    exp_40_ram[2278] = 135;
    exp_40_ram[2279] = 69;
    exp_40_ram[2280] = 1;
    exp_40_ram[2281] = 101;
    exp_40_ram[2282] = 76;
    exp_40_ram[2283] = 214;
    exp_40_ram[2284] = 5;
    exp_40_ram[2285] = 133;
    exp_40_ram[2286] = 1;
    exp_40_ram[2287] = 128;
    exp_40_ram[2288] = 92;
    exp_40_ram[2289] = 5;
    exp_40_ram[2290] = 133;
    exp_40_ram[2291] = 240;
    exp_40_ram[2292] = 240;
    exp_40_ram[2293] = 1;
    exp_40_ram[2294] = 0;
    exp_40_ram[2295] = 0;
    exp_40_ram[2296] = 0;
    exp_40_ram[2297] = 117;
    exp_40_ram[2298] = 110;
    exp_40_ram[2299] = 87;
    exp_40_ram[2300] = 104;
    exp_40_ram[2301] = 105;
    exp_40_ram[2302] = 0;
    exp_40_ram[2303] = 97;
    exp_40_ram[2304] = 98;
    exp_40_ram[2305] = 65;
    exp_40_ram[2306] = 97;
    exp_40_ram[2307] = 110;
    exp_40_ram[2308] = 65;
    exp_40_ram[2309] = 101;
    exp_40_ram[2310] = 116;
    exp_40_ram[2311] = 68;
    exp_40_ram[2312] = 0;
    exp_40_ram[2313] = 35;
    exp_40_ram[2314] = 35;
    exp_40_ram[2315] = 35;
    exp_40_ram[2316] = 35;
    exp_40_ram[2317] = 35;
    exp_40_ram[2318] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 55;
    exp_33_ram[32] = 19;
    exp_33_ram[33] = 239;
    exp_33_ram[34] = 111;
    exp_33_ram[35] = 147;
    exp_33_ram[36] = 147;
    exp_33_ram[37] = 19;
    exp_33_ram[38] = 19;
    exp_33_ram[39] = 19;
    exp_33_ram[40] = 99;
    exp_33_ram[41] = 147;
    exp_33_ram[42] = 99;
    exp_33_ram[43] = 55;
    exp_33_ram[44] = 99;
    exp_33_ram[45] = 19;
    exp_33_ram[46] = 51;
    exp_33_ram[47] = 19;
    exp_33_ram[48] = 51;
    exp_33_ram[49] = 179;
    exp_33_ram[50] = 131;
    exp_33_ram[51] = 19;
    exp_33_ram[52] = 51;
    exp_33_ram[53] = 179;
    exp_33_ram[54] = 99;
    exp_33_ram[55] = 179;
    exp_33_ram[56] = 51;
    exp_33_ram[57] = 51;
    exp_33_ram[58] = 179;
    exp_33_ram[59] = 51;
    exp_33_ram[60] = 147;
    exp_33_ram[61] = 179;
    exp_33_ram[62] = 19;
    exp_33_ram[63] = 19;
    exp_33_ram[64] = 147;
    exp_33_ram[65] = 51;
    exp_33_ram[66] = 19;
    exp_33_ram[67] = 179;
    exp_33_ram[68] = 19;
    exp_33_ram[69] = 179;
    exp_33_ram[70] = 99;
    exp_33_ram[71] = 179;
    exp_33_ram[72] = 19;
    exp_33_ram[73] = 99;
    exp_33_ram[74] = 99;
    exp_33_ram[75] = 19;
    exp_33_ram[76] = 179;
    exp_33_ram[77] = 179;
    exp_33_ram[78] = 51;
    exp_33_ram[79] = 19;
    exp_33_ram[80] = 19;
    exp_33_ram[81] = 179;
    exp_33_ram[82] = 19;
    exp_33_ram[83] = 51;
    exp_33_ram[84] = 179;
    exp_33_ram[85] = 19;
    exp_33_ram[86] = 99;
    exp_33_ram[87] = 51;
    exp_33_ram[88] = 19;
    exp_33_ram[89] = 99;
    exp_33_ram[90] = 99;
    exp_33_ram[91] = 19;
    exp_33_ram[92] = 19;
    exp_33_ram[93] = 51;
    exp_33_ram[94] = 147;
    exp_33_ram[95] = 111;
    exp_33_ram[96] = 55;
    exp_33_ram[97] = 19;
    exp_33_ram[98] = 227;
    exp_33_ram[99] = 19;
    exp_33_ram[100] = 111;
    exp_33_ram[101] = 99;
    exp_33_ram[102] = 19;
    exp_33_ram[103] = 51;
    exp_33_ram[104] = 55;
    exp_33_ram[105] = 99;
    exp_33_ram[106] = 19;
    exp_33_ram[107] = 99;
    exp_33_ram[108] = 19;
    exp_33_ram[109] = 51;
    exp_33_ram[110] = 179;
    exp_33_ram[111] = 3;
    exp_33_ram[112] = 19;
    exp_33_ram[113] = 51;
    exp_33_ram[114] = 179;
    exp_33_ram[115] = 99;
    exp_33_ram[116] = 179;
    exp_33_ram[117] = 147;
    exp_33_ram[118] = 147;
    exp_33_ram[119] = 19;
    exp_33_ram[120] = 19;
    exp_33_ram[121] = 19;
    exp_33_ram[122] = 179;
    exp_33_ram[123] = 179;
    exp_33_ram[124] = 147;
    exp_33_ram[125] = 51;
    exp_33_ram[126] = 51;
    exp_33_ram[127] = 19;
    exp_33_ram[128] = 99;
    exp_33_ram[129] = 51;
    exp_33_ram[130] = 19;
    exp_33_ram[131] = 99;
    exp_33_ram[132] = 99;
    exp_33_ram[133] = 19;
    exp_33_ram[134] = 51;
    exp_33_ram[135] = 51;
    exp_33_ram[136] = 179;
    exp_33_ram[137] = 19;
    exp_33_ram[138] = 19;
    exp_33_ram[139] = 51;
    exp_33_ram[140] = 147;
    exp_33_ram[141] = 51;
    exp_33_ram[142] = 179;
    exp_33_ram[143] = 19;
    exp_33_ram[144] = 99;
    exp_33_ram[145] = 51;
    exp_33_ram[146] = 19;
    exp_33_ram[147] = 99;
    exp_33_ram[148] = 99;
    exp_33_ram[149] = 19;
    exp_33_ram[150] = 19;
    exp_33_ram[151] = 51;
    exp_33_ram[152] = 103;
    exp_33_ram[153] = 55;
    exp_33_ram[154] = 19;
    exp_33_ram[155] = 227;
    exp_33_ram[156] = 19;
    exp_33_ram[157] = 111;
    exp_33_ram[158] = 51;
    exp_33_ram[159] = 51;
    exp_33_ram[160] = 51;
    exp_33_ram[161] = 179;
    exp_33_ram[162] = 51;
    exp_33_ram[163] = 147;
    exp_33_ram[164] = 51;
    exp_33_ram[165] = 51;
    exp_33_ram[166] = 147;
    exp_33_ram[167] = 147;
    exp_33_ram[168] = 147;
    exp_33_ram[169] = 51;
    exp_33_ram[170] = 19;
    exp_33_ram[171] = 51;
    exp_33_ram[172] = 179;
    exp_33_ram[173] = 147;
    exp_33_ram[174] = 99;
    exp_33_ram[175] = 51;
    exp_33_ram[176] = 147;
    exp_33_ram[177] = 99;
    exp_33_ram[178] = 99;
    exp_33_ram[179] = 147;
    exp_33_ram[180] = 51;
    exp_33_ram[181] = 179;
    exp_33_ram[182] = 51;
    exp_33_ram[183] = 19;
    exp_33_ram[184] = 19;
    exp_33_ram[185] = 179;
    exp_33_ram[186] = 19;
    exp_33_ram[187] = 51;
    exp_33_ram[188] = 179;
    exp_33_ram[189] = 19;
    exp_33_ram[190] = 99;
    exp_33_ram[191] = 179;
    exp_33_ram[192] = 19;
    exp_33_ram[193] = 99;
    exp_33_ram[194] = 99;
    exp_33_ram[195] = 19;
    exp_33_ram[196] = 179;
    exp_33_ram[197] = 147;
    exp_33_ram[198] = 179;
    exp_33_ram[199] = 179;
    exp_33_ram[200] = 111;
    exp_33_ram[201] = 99;
    exp_33_ram[202] = 55;
    exp_33_ram[203] = 99;
    exp_33_ram[204] = 19;
    exp_33_ram[205] = 179;
    exp_33_ram[206] = 147;
    exp_33_ram[207] = 51;
    exp_33_ram[208] = 19;
    exp_33_ram[209] = 51;
    exp_33_ram[210] = 3;
    exp_33_ram[211] = 19;
    exp_33_ram[212] = 51;
    exp_33_ram[213] = 179;
    exp_33_ram[214] = 99;
    exp_33_ram[215] = 19;
    exp_33_ram[216] = 227;
    exp_33_ram[217] = 51;
    exp_33_ram[218] = 19;
    exp_33_ram[219] = 111;
    exp_33_ram[220] = 55;
    exp_33_ram[221] = 147;
    exp_33_ram[222] = 227;
    exp_33_ram[223] = 147;
    exp_33_ram[224] = 111;
    exp_33_ram[225] = 51;
    exp_33_ram[226] = 179;
    exp_33_ram[227] = 51;
    exp_33_ram[228] = 51;
    exp_33_ram[229] = 147;
    exp_33_ram[230] = 179;
    exp_33_ram[231] = 179;
    exp_33_ram[232] = 51;
    exp_33_ram[233] = 51;
    exp_33_ram[234] = 51;
    exp_33_ram[235] = 147;
    exp_33_ram[236] = 147;
    exp_33_ram[237] = 19;
    exp_33_ram[238] = 51;
    exp_33_ram[239] = 147;
    exp_33_ram[240] = 51;
    exp_33_ram[241] = 51;
    exp_33_ram[242] = 19;
    exp_33_ram[243] = 99;
    exp_33_ram[244] = 51;
    exp_33_ram[245] = 19;
    exp_33_ram[246] = 99;
    exp_33_ram[247] = 99;
    exp_33_ram[248] = 19;
    exp_33_ram[249] = 51;
    exp_33_ram[250] = 51;
    exp_33_ram[251] = 179;
    exp_33_ram[252] = 51;
    exp_33_ram[253] = 147;
    exp_33_ram[254] = 51;
    exp_33_ram[255] = 147;
    exp_33_ram[256] = 147;
    exp_33_ram[257] = 179;
    exp_33_ram[258] = 19;
    exp_33_ram[259] = 99;
    exp_33_ram[260] = 179;
    exp_33_ram[261] = 19;
    exp_33_ram[262] = 99;
    exp_33_ram[263] = 99;
    exp_33_ram[264] = 19;
    exp_33_ram[265] = 179;
    exp_33_ram[266] = 19;
    exp_33_ram[267] = 183;
    exp_33_ram[268] = 51;
    exp_33_ram[269] = 147;
    exp_33_ram[270] = 51;
    exp_33_ram[271] = 19;
    exp_33_ram[272] = 179;
    exp_33_ram[273] = 19;
    exp_33_ram[274] = 179;
    exp_33_ram[275] = 51;
    exp_33_ram[276] = 179;
    exp_33_ram[277] = 19;
    exp_33_ram[278] = 51;
    exp_33_ram[279] = 51;
    exp_33_ram[280] = 51;
    exp_33_ram[281] = 51;
    exp_33_ram[282] = 99;
    exp_33_ram[283] = 51;
    exp_33_ram[284] = 147;
    exp_33_ram[285] = 51;
    exp_33_ram[286] = 99;
    exp_33_ram[287] = 227;
    exp_33_ram[288] = 183;
    exp_33_ram[289] = 147;
    exp_33_ram[290] = 51;
    exp_33_ram[291] = 19;
    exp_33_ram[292] = 51;
    exp_33_ram[293] = 179;
    exp_33_ram[294] = 51;
    exp_33_ram[295] = 147;
    exp_33_ram[296] = 227;
    exp_33_ram[297] = 19;
    exp_33_ram[298] = 111;
    exp_33_ram[299] = 147;
    exp_33_ram[300] = 19;
    exp_33_ram[301] = 111;
    exp_33_ram[302] = 19;
    exp_33_ram[303] = 19;
    exp_33_ram[304] = 147;
    exp_33_ram[305] = 99;
    exp_33_ram[306] = 51;
    exp_33_ram[307] = 147;
    exp_33_ram[308] = 19;
    exp_33_ram[309] = 227;
    exp_33_ram[310] = 103;
    exp_33_ram[311] = 99;
    exp_33_ram[312] = 99;
    exp_33_ram[313] = 19;
    exp_33_ram[314] = 147;
    exp_33_ram[315] = 19;
    exp_33_ram[316] = 99;
    exp_33_ram[317] = 147;
    exp_33_ram[318] = 99;
    exp_33_ram[319] = 99;
    exp_33_ram[320] = 19;
    exp_33_ram[321] = 147;
    exp_33_ram[322] = 227;
    exp_33_ram[323] = 19;
    exp_33_ram[324] = 99;
    exp_33_ram[325] = 179;
    exp_33_ram[326] = 51;
    exp_33_ram[327] = 147;
    exp_33_ram[328] = 19;
    exp_33_ram[329] = 227;
    exp_33_ram[330] = 103;
    exp_33_ram[331] = 147;
    exp_33_ram[332] = 239;
    exp_33_ram[333] = 19;
    exp_33_ram[334] = 103;
    exp_33_ram[335] = 51;
    exp_33_ram[336] = 99;
    exp_33_ram[337] = 179;
    exp_33_ram[338] = 111;
    exp_33_ram[339] = 179;
    exp_33_ram[340] = 147;
    exp_33_ram[341] = 239;
    exp_33_ram[342] = 51;
    exp_33_ram[343] = 103;
    exp_33_ram[344] = 147;
    exp_33_ram[345] = 99;
    exp_33_ram[346] = 99;
    exp_33_ram[347] = 239;
    exp_33_ram[348] = 19;
    exp_33_ram[349] = 103;
    exp_33_ram[350] = 179;
    exp_33_ram[351] = 227;
    exp_33_ram[352] = 51;
    exp_33_ram[353] = 239;
    exp_33_ram[354] = 51;
    exp_33_ram[355] = 103;
    exp_33_ram[356] = 72;
    exp_33_ram[357] = 111;
    exp_33_ram[358] = 114;
    exp_33_ram[359] = 0;
    exp_33_ram[360] = 114;
    exp_33_ram[361] = 105;
    exp_33_ram[362] = 107;
    exp_33_ram[363] = 104;
    exp_33_ram[364] = 105;
    exp_33_ram[365] = 32;
    exp_33_ram[366] = 111;
    exp_33_ram[367] = 0;
    exp_33_ram[368] = 37;
    exp_33_ram[369] = 37;
    exp_33_ram[370] = 50;
    exp_33_ram[371] = 116;
    exp_33_ram[372] = 116;
    exp_33_ram[373] = 114;
    exp_33_ram[374] = 108;
    exp_33_ram[375] = 108;
    exp_33_ram[376] = 32;
    exp_33_ram[377] = 49;
    exp_33_ram[378] = 99;
    exp_33_ram[379] = 10;
    exp_33_ram[380] = 37;
    exp_33_ram[381] = 52;
    exp_33_ram[382] = 116;
    exp_33_ram[383] = 116;
    exp_33_ram[384] = 114;
    exp_33_ram[385] = 108;
    exp_33_ram[386] = 108;
    exp_33_ram[387] = 32;
    exp_33_ram[388] = 49;
    exp_33_ram[389] = 99;
    exp_33_ram[390] = 10;
    exp_33_ram[391] = 37;
    exp_33_ram[392] = 50;
    exp_33_ram[393] = 116;
    exp_33_ram[394] = 116;
    exp_33_ram[395] = 114;
    exp_33_ram[396] = 118;
    exp_33_ram[397] = 115;
    exp_33_ram[398] = 32;
    exp_33_ram[399] = 101;
    exp_33_ram[400] = 100;
    exp_33_ram[401] = 37;
    exp_33_ram[402] = 52;
    exp_33_ram[403] = 116;
    exp_33_ram[404] = 116;
    exp_33_ram[405] = 114;
    exp_33_ram[406] = 118;
    exp_33_ram[407] = 115;
    exp_33_ram[408] = 32;
    exp_33_ram[409] = 101;
    exp_33_ram[410] = 100;
    exp_33_ram[411] = 97;
    exp_33_ram[412] = 110;
    exp_33_ram[413] = 116;
    exp_33_ram[414] = 46;
    exp_33_ram[415] = 102;
    exp_33_ram[416] = 0;
    exp_33_ram[417] = 112;
    exp_33_ram[418] = 0;
    exp_33_ram[419] = 65;
    exp_33_ram[420] = 99;
    exp_33_ram[421] = 100;
    exp_33_ram[422] = 56;
    exp_33_ram[423] = 48;
    exp_33_ram[424] = 37;
    exp_33_ram[425] = 10;
    exp_33_ram[426] = 10;
    exp_33_ram[427] = 112;
    exp_33_ram[428] = 32;
    exp_33_ram[429] = 111;
    exp_33_ram[430] = 10;
    exp_33_ram[431] = 72;
    exp_33_ram[432] = 111;
    exp_33_ram[433] = 114;
    exp_33_ram[434] = 98;
    exp_33_ram[435] = 110;
    exp_33_ram[436] = 116;
    exp_33_ram[437] = 100;
    exp_33_ram[438] = 99;
    exp_33_ram[439] = 116;
    exp_33_ram[440] = 87;
    exp_33_ram[441] = 104;
    exp_33_ram[442] = 100;
    exp_33_ram[443] = 101;
    exp_33_ram[444] = 77;
    exp_33_ram[445] = 105;
    exp_33_ram[446] = 99;
    exp_33_ram[447] = 111;
    exp_33_ram[448] = 101;
    exp_33_ram[449] = 101;
    exp_33_ram[450] = 77;
    exp_33_ram[451] = 114;
    exp_33_ram[452] = 0;
    exp_33_ram[453] = 3;
    exp_33_ram[454] = 4;
    exp_33_ram[455] = 4;
    exp_33_ram[456] = 5;
    exp_33_ram[457] = 5;
    exp_33_ram[458] = 5;
    exp_33_ram[459] = 5;
    exp_33_ram[460] = 6;
    exp_33_ram[461] = 6;
    exp_33_ram[462] = 6;
    exp_33_ram[463] = 6;
    exp_33_ram[464] = 6;
    exp_33_ram[465] = 6;
    exp_33_ram[466] = 6;
    exp_33_ram[467] = 6;
    exp_33_ram[468] = 7;
    exp_33_ram[469] = 7;
    exp_33_ram[470] = 7;
    exp_33_ram[471] = 7;
    exp_33_ram[472] = 7;
    exp_33_ram[473] = 7;
    exp_33_ram[474] = 7;
    exp_33_ram[475] = 7;
    exp_33_ram[476] = 7;
    exp_33_ram[477] = 7;
    exp_33_ram[478] = 7;
    exp_33_ram[479] = 7;
    exp_33_ram[480] = 7;
    exp_33_ram[481] = 7;
    exp_33_ram[482] = 7;
    exp_33_ram[483] = 7;
    exp_33_ram[484] = 8;
    exp_33_ram[485] = 8;
    exp_33_ram[486] = 8;
    exp_33_ram[487] = 8;
    exp_33_ram[488] = 8;
    exp_33_ram[489] = 8;
    exp_33_ram[490] = 8;
    exp_33_ram[491] = 8;
    exp_33_ram[492] = 8;
    exp_33_ram[493] = 8;
    exp_33_ram[494] = 8;
    exp_33_ram[495] = 8;
    exp_33_ram[496] = 8;
    exp_33_ram[497] = 8;
    exp_33_ram[498] = 8;
    exp_33_ram[499] = 8;
    exp_33_ram[500] = 8;
    exp_33_ram[501] = 8;
    exp_33_ram[502] = 8;
    exp_33_ram[503] = 8;
    exp_33_ram[504] = 8;
    exp_33_ram[505] = 8;
    exp_33_ram[506] = 8;
    exp_33_ram[507] = 8;
    exp_33_ram[508] = 8;
    exp_33_ram[509] = 8;
    exp_33_ram[510] = 8;
    exp_33_ram[511] = 8;
    exp_33_ram[512] = 8;
    exp_33_ram[513] = 8;
    exp_33_ram[514] = 8;
    exp_33_ram[515] = 8;
    exp_33_ram[516] = 35;
    exp_33_ram[517] = 103;
    exp_33_ram[518] = 183;
    exp_33_ram[519] = 131;
    exp_33_ram[520] = 3;
    exp_33_ram[521] = 103;
    exp_33_ram[522] = 147;
    exp_33_ram[523] = 19;
    exp_33_ram[524] = 51;
    exp_33_ram[525] = 3;
    exp_33_ram[526] = 99;
    exp_33_ram[527] = 103;
    exp_33_ram[528] = 19;
    exp_33_ram[529] = 35;
    exp_33_ram[530] = 111;
    exp_33_ram[531] = 19;
    exp_33_ram[532] = 183;
    exp_33_ram[533] = 35;
    exp_33_ram[534] = 3;
    exp_33_ram[535] = 35;
    exp_33_ram[536] = 147;
    exp_33_ram[537] = 239;
    exp_33_ram[538] = 147;
    exp_33_ram[539] = 131;
    exp_33_ram[540] = 35;
    exp_33_ram[541] = 3;
    exp_33_ram[542] = 19;
    exp_33_ram[543] = 19;
    exp_33_ram[544] = 103;
    exp_33_ram[545] = 19;
    exp_33_ram[546] = 35;
    exp_33_ram[547] = 35;
    exp_33_ram[548] = 19;
    exp_33_ram[549] = 99;
    exp_33_ram[550] = 239;
    exp_33_ram[551] = 131;
    exp_33_ram[552] = 19;
    exp_33_ram[553] = 3;
    exp_33_ram[554] = 19;
    exp_33_ram[555] = 103;
    exp_33_ram[556] = 179;
    exp_33_ram[557] = 35;
    exp_33_ram[558] = 51;
    exp_33_ram[559] = 35;
    exp_33_ram[560] = 111;
    exp_33_ram[561] = 19;
    exp_33_ram[562] = 35;
    exp_33_ram[563] = 35;
    exp_33_ram[564] = 35;
    exp_33_ram[565] = 35;
    exp_33_ram[566] = 35;
    exp_33_ram[567] = 35;
    exp_33_ram[568] = 35;
    exp_33_ram[569] = 147;
    exp_33_ram[570] = 35;
    exp_33_ram[571] = 35;
    exp_33_ram[572] = 35;
    exp_33_ram[573] = 35;
    exp_33_ram[574] = 35;
    exp_33_ram[575] = 35;
    exp_33_ram[576] = 147;
    exp_33_ram[577] = 19;
    exp_33_ram[578] = 147;
    exp_33_ram[579] = 19;
    exp_33_ram[580] = 147;
    exp_33_ram[581] = 19;
    exp_33_ram[582] = 19;
    exp_33_ram[583] = 19;
    exp_33_ram[584] = 99;
    exp_33_ram[585] = 147;
    exp_33_ram[586] = 99;
    exp_33_ram[587] = 19;
    exp_33_ram[588] = 183;
    exp_33_ram[589] = 147;
    exp_33_ram[590] = 19;
    exp_33_ram[591] = 147;
    exp_33_ram[592] = 111;
    exp_33_ram[593] = 147;
    exp_33_ram[594] = 179;
    exp_33_ram[595] = 19;
    exp_33_ram[596] = 99;
    exp_33_ram[597] = 99;
    exp_33_ram[598] = 99;
    exp_33_ram[599] = 147;
    exp_33_ram[600] = 99;
    exp_33_ram[601] = 19;
    exp_33_ram[602] = 19;
    exp_33_ram[603] = 147;
    exp_33_ram[604] = 19;
    exp_33_ram[605] = 147;
    exp_33_ram[606] = 19;
    exp_33_ram[607] = 239;
    exp_33_ram[608] = 147;
    exp_33_ram[609] = 179;
    exp_33_ram[610] = 19;
    exp_33_ram[611] = 179;
    exp_33_ram[612] = 227;
    exp_33_ram[613] = 131;
    exp_33_ram[614] = 3;
    exp_33_ram[615] = 131;
    exp_33_ram[616] = 3;
    exp_33_ram[617] = 131;
    exp_33_ram[618] = 3;
    exp_33_ram[619] = 131;
    exp_33_ram[620] = 3;
    exp_33_ram[621] = 131;
    exp_33_ram[622] = 3;
    exp_33_ram[623] = 131;
    exp_33_ram[624] = 3;
    exp_33_ram[625] = 131;
    exp_33_ram[626] = 19;
    exp_33_ram[627] = 103;
    exp_33_ram[628] = 99;
    exp_33_ram[629] = 19;
    exp_33_ram[630] = 111;
    exp_33_ram[631] = 19;
    exp_33_ram[632] = 111;
    exp_33_ram[633] = 227;
    exp_33_ram[634] = 147;
    exp_33_ram[635] = 19;
    exp_33_ram[636] = 147;
    exp_33_ram[637] = 19;
    exp_33_ram[638] = 239;
    exp_33_ram[639] = 111;
    exp_33_ram[640] = 19;
    exp_33_ram[641] = 183;
    exp_33_ram[642] = 111;
    exp_33_ram[643] = 183;
    exp_33_ram[644] = 19;
    exp_33_ram[645] = 147;
    exp_33_ram[646] = 19;
    exp_33_ram[647] = 111;
    exp_33_ram[648] = 131;
    exp_33_ram[649] = 99;
    exp_33_ram[650] = 19;
    exp_33_ram[651] = 35;
    exp_33_ram[652] = 35;
    exp_33_ram[653] = 35;
    exp_33_ram[654] = 35;
    exp_33_ram[655] = 35;
    exp_33_ram[656] = 35;
    exp_33_ram[657] = 35;
    exp_33_ram[658] = 35;
    exp_33_ram[659] = 35;
    exp_33_ram[660] = 147;
    exp_33_ram[661] = 35;
    exp_33_ram[662] = 35;
    exp_33_ram[663] = 35;
    exp_33_ram[664] = 35;
    exp_33_ram[665] = 19;
    exp_33_ram[666] = 147;
    exp_33_ram[667] = 147;
    exp_33_ram[668] = 19;
    exp_33_ram[669] = 19;
    exp_33_ram[670] = 147;
    exp_33_ram[671] = 19;
    exp_33_ram[672] = 147;
    exp_33_ram[673] = 19;
    exp_33_ram[674] = 147;
    exp_33_ram[675] = 179;
    exp_33_ram[676] = 3;
    exp_33_ram[677] = 19;
    exp_33_ram[678] = 51;
    exp_33_ram[679] = 99;
    exp_33_ram[680] = 131;
    exp_33_ram[681] = 99;
    exp_33_ram[682] = 147;
    exp_33_ram[683] = 99;
    exp_33_ram[684] = 19;
    exp_33_ram[685] = 51;
    exp_33_ram[686] = 3;
    exp_33_ram[687] = 99;
    exp_33_ram[688] = 131;
    exp_33_ram[689] = 3;
    exp_33_ram[690] = 131;
    exp_33_ram[691] = 3;
    exp_33_ram[692] = 131;
    exp_33_ram[693] = 3;
    exp_33_ram[694] = 131;
    exp_33_ram[695] = 3;
    exp_33_ram[696] = 131;
    exp_33_ram[697] = 3;
    exp_33_ram[698] = 131;
    exp_33_ram[699] = 3;
    exp_33_ram[700] = 131;
    exp_33_ram[701] = 19;
    exp_33_ram[702] = 19;
    exp_33_ram[703] = 103;
    exp_33_ram[704] = 147;
    exp_33_ram[705] = 147;
    exp_33_ram[706] = 19;
    exp_33_ram[707] = 239;
    exp_33_ram[708] = 19;
    exp_33_ram[709] = 131;
    exp_33_ram[710] = 227;
    exp_33_ram[711] = 19;
    exp_33_ram[712] = 111;
    exp_33_ram[713] = 147;
    exp_33_ram[714] = 19;
    exp_33_ram[715] = 179;
    exp_33_ram[716] = 131;
    exp_33_ram[717] = 19;
    exp_33_ram[718] = 51;
    exp_33_ram[719] = 147;
    exp_33_ram[720] = 99;
    exp_33_ram[721] = 99;
    exp_33_ram[722] = 99;
    exp_33_ram[723] = 147;
    exp_33_ram[724] = 99;
    exp_33_ram[725] = 99;
    exp_33_ram[726] = 99;
    exp_33_ram[727] = 147;
    exp_33_ram[728] = 227;
    exp_33_ram[729] = 19;
    exp_33_ram[730] = 147;
    exp_33_ram[731] = 111;
    exp_33_ram[732] = 51;
    exp_33_ram[733] = 131;
    exp_33_ram[734] = 51;
    exp_33_ram[735] = 227;
    exp_33_ram[736] = 111;
    exp_33_ram[737] = 147;
    exp_33_ram[738] = 227;
    exp_33_ram[739] = 19;
    exp_33_ram[740] = 131;
    exp_33_ram[741] = 99;
    exp_33_ram[742] = 147;
    exp_33_ram[743] = 147;
    exp_33_ram[744] = 19;
    exp_33_ram[745] = 19;
    exp_33_ram[746] = 35;
    exp_33_ram[747] = 35;
    exp_33_ram[748] = 239;
    exp_33_ram[749] = 3;
    exp_33_ram[750] = 131;
    exp_33_ram[751] = 19;
    exp_33_ram[752] = 147;
    exp_33_ram[753] = 19;
    exp_33_ram[754] = 19;
    exp_33_ram[755] = 179;
    exp_33_ram[756] = 147;
    exp_33_ram[757] = 19;
    exp_33_ram[758] = 239;
    exp_33_ram[759] = 111;
    exp_33_ram[760] = 99;
    exp_33_ram[761] = 99;
    exp_33_ram[762] = 147;
    exp_33_ram[763] = 99;
    exp_33_ram[764] = 147;
    exp_33_ram[765] = 227;
    exp_33_ram[766] = 3;
    exp_33_ram[767] = 147;
    exp_33_ram[768] = 3;
    exp_33_ram[769] = 99;
    exp_33_ram[770] = 147;
    exp_33_ram[771] = 111;
    exp_33_ram[772] = 147;
    exp_33_ram[773] = 227;
    exp_33_ram[774] = 19;
    exp_33_ram[775] = 147;
    exp_33_ram[776] = 19;
    exp_33_ram[777] = 111;
    exp_33_ram[778] = 147;
    exp_33_ram[779] = 147;
    exp_33_ram[780] = 19;
    exp_33_ram[781] = 19;
    exp_33_ram[782] = 111;
    exp_33_ram[783] = 3;
    exp_33_ram[784] = 147;
    exp_33_ram[785] = 147;
    exp_33_ram[786] = 19;
    exp_33_ram[787] = 19;
    exp_33_ram[788] = 239;
    exp_33_ram[789] = 19;
    exp_33_ram[790] = 147;
    exp_33_ram[791] = 111;
    exp_33_ram[792] = 147;
    exp_33_ram[793] = 147;
    exp_33_ram[794] = 19;
    exp_33_ram[795] = 35;
    exp_33_ram[796] = 239;
    exp_33_ram[797] = 131;
    exp_33_ram[798] = 19;
    exp_33_ram[799] = 19;
    exp_33_ram[800] = 111;
    exp_33_ram[801] = 147;
    exp_33_ram[802] = 19;
    exp_33_ram[803] = 147;
    exp_33_ram[804] = 111;
    exp_33_ram[805] = 19;
    exp_33_ram[806] = 147;
    exp_33_ram[807] = 19;
    exp_33_ram[808] = 131;
    exp_33_ram[809] = 111;
    exp_33_ram[810] = 19;
    exp_33_ram[811] = 147;
    exp_33_ram[812] = 19;
    exp_33_ram[813] = 111;
    exp_33_ram[814] = 19;
    exp_33_ram[815] = 19;
    exp_33_ram[816] = 103;
    exp_33_ram[817] = 19;
    exp_33_ram[818] = 35;
    exp_33_ram[819] = 183;
    exp_33_ram[820] = 35;
    exp_33_ram[821] = 19;
    exp_33_ram[822] = 3;
    exp_33_ram[823] = 35;
    exp_33_ram[824] = 35;
    exp_33_ram[825] = 147;
    exp_33_ram[826] = 147;
    exp_33_ram[827] = 35;
    exp_33_ram[828] = 35;
    exp_33_ram[829] = 35;
    exp_33_ram[830] = 35;
    exp_33_ram[831] = 35;
    exp_33_ram[832] = 239;
    exp_33_ram[833] = 131;
    exp_33_ram[834] = 19;
    exp_33_ram[835] = 103;
    exp_33_ram[836] = 147;
    exp_33_ram[837] = 147;
    exp_33_ram[838] = 55;
    exp_33_ram[839] = 19;
    exp_33_ram[840] = 99;
    exp_33_ram[841] = 19;
    exp_33_ram[842] = 19;
    exp_33_ram[843] = 51;
    exp_33_ram[844] = 103;
    exp_33_ram[845] = 55;
    exp_33_ram[846] = 3;
    exp_33_ram[847] = 3;
    exp_33_ram[848] = 99;
    exp_33_ram[849] = 19;
    exp_33_ram[850] = 35;
    exp_33_ram[851] = 183;
    exp_33_ram[852] = 19;
    exp_33_ram[853] = 147;
    exp_33_ram[854] = 183;
    exp_33_ram[855] = 227;
    exp_33_ram[856] = 147;
    exp_33_ram[857] = 179;
    exp_33_ram[858] = 3;
    exp_33_ram[859] = 51;
    exp_33_ram[860] = 99;
    exp_33_ram[861] = 51;
    exp_33_ram[862] = 99;
    exp_33_ram[863] = 51;
    exp_33_ram[864] = 19;
    exp_33_ram[865] = 111;
    exp_33_ram[866] = 179;
    exp_33_ram[867] = 35;
    exp_33_ram[868] = 99;
    exp_33_ram[869] = 179;
    exp_33_ram[870] = 147;
    exp_33_ram[871] = 147;
    exp_33_ram[872] = 147;
    exp_33_ram[873] = 179;
    exp_33_ram[874] = 179;
    exp_33_ram[875] = 35;
    exp_33_ram[876] = 19;
    exp_33_ram[877] = 111;
    exp_33_ram[878] = 55;
    exp_33_ram[879] = 147;
    exp_33_ram[880] = 51;
    exp_33_ram[881] = 19;
    exp_33_ram[882] = 19;
    exp_33_ram[883] = 51;
    exp_33_ram[884] = 131;
    exp_33_ram[885] = 183;
    exp_33_ram[886] = 147;
    exp_33_ram[887] = 179;
    exp_33_ram[888] = 35;
    exp_33_ram[889] = 183;
    exp_33_ram[890] = 131;
    exp_33_ram[891] = 19;
    exp_33_ram[892] = 147;
    exp_33_ram[893] = 55;
    exp_33_ram[894] = 19;
    exp_33_ram[895] = 99;
    exp_33_ram[896] = 147;
    exp_33_ram[897] = 179;
    exp_33_ram[898] = 3;
    exp_33_ram[899] = 179;
    exp_33_ram[900] = 179;
    exp_33_ram[901] = 51;
    exp_33_ram[902] = 147;
    exp_33_ram[903] = 227;
    exp_33_ram[904] = 19;
    exp_33_ram[905] = 51;
    exp_33_ram[906] = 99;
    exp_33_ram[907] = 19;
    exp_33_ram[908] = 51;
    exp_33_ram[909] = 3;
    exp_33_ram[910] = 51;
    exp_33_ram[911] = 51;
    exp_33_ram[912] = 227;
    exp_33_ram[913] = 179;
    exp_33_ram[914] = 147;
    exp_33_ram[915] = 19;
    exp_33_ram[916] = 35;
    exp_33_ram[917] = 179;
    exp_33_ram[918] = 111;
    exp_33_ram[919] = 103;
    exp_33_ram[920] = 179;
    exp_33_ram[921] = 147;
    exp_33_ram[922] = 147;
    exp_33_ram[923] = 99;
    exp_33_ram[924] = 19;
    exp_33_ram[925] = 51;
    exp_33_ram[926] = 19;
    exp_33_ram[927] = 111;
    exp_33_ram[928] = 131;
    exp_33_ram[929] = 19;
    exp_33_ram[930] = 147;
    exp_33_ram[931] = 35;
    exp_33_ram[932] = 131;
    exp_33_ram[933] = 35;
    exp_33_ram[934] = 131;
    exp_33_ram[935] = 35;
    exp_33_ram[936] = 131;
    exp_33_ram[937] = 35;
    exp_33_ram[938] = 179;
    exp_33_ram[939] = 227;
    exp_33_ram[940] = 19;
    exp_33_ram[941] = 19;
    exp_33_ram[942] = 179;
    exp_33_ram[943] = 179;
    exp_33_ram[944] = 19;
    exp_33_ram[945] = 51;
    exp_33_ram[946] = 99;
    exp_33_ram[947] = 19;
    exp_33_ram[948] = 19;
    exp_33_ram[949] = 179;
    exp_33_ram[950] = 179;
    exp_33_ram[951] = 147;
    exp_33_ram[952] = 99;
    exp_33_ram[953] = 103;
    exp_33_ram[954] = 51;
    exp_33_ram[955] = 131;
    exp_33_ram[956] = 51;
    exp_33_ram[957] = 147;
    exp_33_ram[958] = 35;
    exp_33_ram[959] = 111;
    exp_33_ram[960] = 51;
    exp_33_ram[961] = 3;
    exp_33_ram[962] = 51;
    exp_33_ram[963] = 147;
    exp_33_ram[964] = 35;
    exp_33_ram[965] = 111;
    exp_33_ram[966] = 147;
    exp_33_ram[967] = 99;
    exp_33_ram[968] = 19;
    exp_33_ram[969] = 147;
    exp_33_ram[970] = 35;
    exp_33_ram[971] = 35;
    exp_33_ram[972] = 19;
    exp_33_ram[973] = 239;
    exp_33_ram[974] = 147;
    exp_33_ram[975] = 99;
    exp_33_ram[976] = 147;
    exp_33_ram[977] = 19;
    exp_33_ram[978] = 239;
    exp_33_ram[979] = 147;
    exp_33_ram[980] = 131;
    exp_33_ram[981] = 3;
    exp_33_ram[982] = 19;
    exp_33_ram[983] = 19;
    exp_33_ram[984] = 103;
    exp_33_ram[985] = 147;
    exp_33_ram[986] = 19;
    exp_33_ram[987] = 103;
    exp_33_ram[988] = 147;
    exp_33_ram[989] = 147;
    exp_33_ram[990] = 99;
    exp_33_ram[991] = 19;
    exp_33_ram[992] = 147;
    exp_33_ram[993] = 147;
    exp_33_ram[994] = 99;
    exp_33_ram[995] = 19;
    exp_33_ram[996] = 147;
    exp_33_ram[997] = 99;
    exp_33_ram[998] = 19;
    exp_33_ram[999] = 35;
    exp_33_ram[1000] = 239;
    exp_33_ram[1001] = 131;
    exp_33_ram[1002] = 179;
    exp_33_ram[1003] = 147;
    exp_33_ram[1004] = 19;
    exp_33_ram[1005] = 19;
    exp_33_ram[1006] = 103;
    exp_33_ram[1007] = 147;
    exp_33_ram[1008] = 19;
    exp_33_ram[1009] = 103;
    exp_33_ram[1010] = 183;
    exp_33_ram[1011] = 3;
    exp_33_ram[1012] = 131;
    exp_33_ram[1013] = 131;
    exp_33_ram[1014] = 19;
    exp_33_ram[1015] = 131;
    exp_33_ram[1016] = 179;
    exp_33_ram[1017] = 103;
    exp_33_ram[1018] = 19;
    exp_33_ram[1019] = 35;
    exp_33_ram[1020] = 131;
    exp_33_ram[1021] = 35;
    exp_33_ram[1022] = 183;
    exp_33_ram[1023] = 35;
    exp_33_ram[1024] = 35;
    exp_33_ram[1025] = 35;
    exp_33_ram[1026] = 35;
    exp_33_ram[1027] = 35;
    exp_33_ram[1028] = 35;
    exp_33_ram[1029] = 19;
    exp_33_ram[1030] = 19;
    exp_33_ram[1031] = 19;
    exp_33_ram[1032] = 147;
    exp_33_ram[1033] = 147;
    exp_33_ram[1034] = 147;
    exp_33_ram[1035] = 99;
    exp_33_ram[1036] = 3;
    exp_33_ram[1037] = 183;
    exp_33_ram[1038] = 147;
    exp_33_ram[1039] = 147;
    exp_33_ram[1040] = 99;
    exp_33_ram[1041] = 147;
    exp_33_ram[1042] = 19;
    exp_33_ram[1043] = 239;
    exp_33_ram[1044] = 147;
    exp_33_ram[1045] = 239;
    exp_33_ram[1046] = 51;
    exp_33_ram[1047] = 179;
    exp_33_ram[1048] = 179;
    exp_33_ram[1049] = 19;
    exp_33_ram[1050] = 147;
    exp_33_ram[1051] = 111;
    exp_33_ram[1052] = 19;
    exp_33_ram[1053] = 239;
    exp_33_ram[1054] = 51;
    exp_33_ram[1055] = 147;
    exp_33_ram[1056] = 19;
    exp_33_ram[1057] = 239;
    exp_33_ram[1058] = 51;
    exp_33_ram[1059] = 179;
    exp_33_ram[1060] = 179;
    exp_33_ram[1061] = 19;
    exp_33_ram[1062] = 19;
    exp_33_ram[1063] = 111;
    exp_33_ram[1064] = 3;
    exp_33_ram[1065] = 3;
    exp_33_ram[1066] = 131;
    exp_33_ram[1067] = 147;
    exp_33_ram[1068] = 179;
    exp_33_ram[1069] = 147;
    exp_33_ram[1070] = 179;
    exp_33_ram[1071] = 19;
    exp_33_ram[1072] = 51;
    exp_33_ram[1073] = 147;
    exp_33_ram[1074] = 19;
    exp_33_ram[1075] = 3;
    exp_33_ram[1076] = 19;
    exp_33_ram[1077] = 147;
    exp_33_ram[1078] = 51;
    exp_33_ram[1079] = 179;
    exp_33_ram[1080] = 179;
    exp_33_ram[1081] = 179;
    exp_33_ram[1082] = 183;
    exp_33_ram[1083] = 147;
    exp_33_ram[1084] = 179;
    exp_33_ram[1085] = 51;
    exp_33_ram[1086] = 179;
    exp_33_ram[1087] = 147;
    exp_33_ram[1088] = 19;
    exp_33_ram[1089] = 51;
    exp_33_ram[1090] = 239;
    exp_33_ram[1091] = 179;
    exp_33_ram[1092] = 147;
    exp_33_ram[1093] = 179;
    exp_33_ram[1094] = 179;
    exp_33_ram[1095] = 51;
    exp_33_ram[1096] = 51;
    exp_33_ram[1097] = 51;
    exp_33_ram[1098] = 179;
    exp_33_ram[1099] = 131;
    exp_33_ram[1100] = 179;
    exp_33_ram[1101] = 3;
    exp_33_ram[1102] = 131;
    exp_33_ram[1103] = 3;
    exp_33_ram[1104] = 131;
    exp_33_ram[1105] = 3;
    exp_33_ram[1106] = 131;
    exp_33_ram[1107] = 3;
    exp_33_ram[1108] = 19;
    exp_33_ram[1109] = 103;
    exp_33_ram[1110] = 19;
    exp_33_ram[1111] = 35;
    exp_33_ram[1112] = 35;
    exp_33_ram[1113] = 19;
    exp_33_ram[1114] = 239;
    exp_33_ram[1115] = 183;
    exp_33_ram[1116] = 3;
    exp_33_ram[1117] = 147;
    exp_33_ram[1118] = 239;
    exp_33_ram[1119] = 183;
    exp_33_ram[1120] = 131;
    exp_33_ram[1121] = 51;
    exp_33_ram[1122] = 99;
    exp_33_ram[1123] = 35;
    exp_33_ram[1124] = 35;
    exp_33_ram[1125] = 131;
    exp_33_ram[1126] = 3;
    exp_33_ram[1127] = 147;
    exp_33_ram[1128] = 19;
    exp_33_ram[1129] = 103;
    exp_33_ram[1130] = 19;
    exp_33_ram[1131] = 35;
    exp_33_ram[1132] = 147;
    exp_33_ram[1133] = 19;
    exp_33_ram[1134] = 35;
    exp_33_ram[1135] = 35;
    exp_33_ram[1136] = 19;
    exp_33_ram[1137] = 239;
    exp_33_ram[1138] = 51;
    exp_33_ram[1139] = 179;
    exp_33_ram[1140] = 183;
    exp_33_ram[1141] = 51;
    exp_33_ram[1142] = 51;
    exp_33_ram[1143] = 147;
    exp_33_ram[1144] = 131;
    exp_33_ram[1145] = 35;
    exp_33_ram[1146] = 3;
    exp_33_ram[1147] = 35;
    exp_33_ram[1148] = 131;
    exp_33_ram[1149] = 19;
    exp_33_ram[1150] = 103;
    exp_33_ram[1151] = 19;
    exp_33_ram[1152] = 183;
    exp_33_ram[1153] = 35;
    exp_33_ram[1154] = 19;
    exp_33_ram[1155] = 147;
    exp_33_ram[1156] = 147;
    exp_33_ram[1157] = 19;
    exp_33_ram[1158] = 35;
    exp_33_ram[1159] = 35;
    exp_33_ram[1160] = 35;
    exp_33_ram[1161] = 35;
    exp_33_ram[1162] = 35;
    exp_33_ram[1163] = 239;
    exp_33_ram[1164] = 183;
    exp_33_ram[1165] = 19;
    exp_33_ram[1166] = 147;
    exp_33_ram[1167] = 19;
    exp_33_ram[1168] = 239;
    exp_33_ram[1169] = 131;
    exp_33_ram[1170] = 183;
    exp_33_ram[1171] = 19;
    exp_33_ram[1172] = 147;
    exp_33_ram[1173] = 179;
    exp_33_ram[1174] = 147;
    exp_33_ram[1175] = 19;
    exp_33_ram[1176] = 179;
    exp_33_ram[1177] = 19;
    exp_33_ram[1178] = 19;
    exp_33_ram[1179] = 239;
    exp_33_ram[1180] = 163;
    exp_33_ram[1181] = 131;
    exp_33_ram[1182] = 19;
    exp_33_ram[1183] = 19;
    exp_33_ram[1184] = 147;
    exp_33_ram[1185] = 179;
    exp_33_ram[1186] = 147;
    exp_33_ram[1187] = 179;
    exp_33_ram[1188] = 239;
    exp_33_ram[1189] = 163;
    exp_33_ram[1190] = 3;
    exp_33_ram[1191] = 147;
    exp_33_ram[1192] = 19;
    exp_33_ram[1193] = 239;
    exp_33_ram[1194] = 35;
    exp_33_ram[1195] = 131;
    exp_33_ram[1196] = 35;
    exp_33_ram[1197] = 35;
    exp_33_ram[1198] = 147;
    exp_33_ram[1199] = 35;
    exp_33_ram[1200] = 131;
    exp_33_ram[1201] = 147;
    exp_33_ram[1202] = 147;
    exp_33_ram[1203] = 163;
    exp_33_ram[1204] = 3;
    exp_33_ram[1205] = 239;
    exp_33_ram[1206] = 35;
    exp_33_ram[1207] = 131;
    exp_33_ram[1208] = 35;
    exp_33_ram[1209] = 163;
    exp_33_ram[1210] = 147;
    exp_33_ram[1211] = 163;
    exp_33_ram[1212] = 131;
    exp_33_ram[1213] = 147;
    exp_33_ram[1214] = 147;
    exp_33_ram[1215] = 35;
    exp_33_ram[1216] = 3;
    exp_33_ram[1217] = 239;
    exp_33_ram[1218] = 35;
    exp_33_ram[1219] = 131;
    exp_33_ram[1220] = 35;
    exp_33_ram[1221] = 35;
    exp_33_ram[1222] = 147;
    exp_33_ram[1223] = 35;
    exp_33_ram[1224] = 131;
    exp_33_ram[1225] = 147;
    exp_33_ram[1226] = 147;
    exp_33_ram[1227] = 163;
    exp_33_ram[1228] = 3;
    exp_33_ram[1229] = 239;
    exp_33_ram[1230] = 35;
    exp_33_ram[1231] = 131;
    exp_33_ram[1232] = 35;
    exp_33_ram[1233] = 163;
    exp_33_ram[1234] = 147;
    exp_33_ram[1235] = 163;
    exp_33_ram[1236] = 131;
    exp_33_ram[1237] = 147;
    exp_33_ram[1238] = 147;
    exp_33_ram[1239] = 35;
    exp_33_ram[1240] = 3;
    exp_33_ram[1241] = 19;
    exp_33_ram[1242] = 239;
    exp_33_ram[1243] = 35;
    exp_33_ram[1244] = 35;
    exp_33_ram[1245] = 131;
    exp_33_ram[1246] = 3;
    exp_33_ram[1247] = 147;
    exp_33_ram[1248] = 147;
    exp_33_ram[1249] = 35;
    exp_33_ram[1250] = 239;
    exp_33_ram[1251] = 35;
    exp_33_ram[1252] = 35;
    exp_33_ram[1253] = 131;
    exp_33_ram[1254] = 3;
    exp_33_ram[1255] = 147;
    exp_33_ram[1256] = 147;
    exp_33_ram[1257] = 163;
    exp_33_ram[1258] = 239;
    exp_33_ram[1259] = 35;
    exp_33_ram[1260] = 131;
    exp_33_ram[1261] = 35;
    exp_33_ram[1262] = 131;
    exp_33_ram[1263] = 147;
    exp_33_ram[1264] = 35;
    exp_33_ram[1265] = 131;
    exp_33_ram[1266] = 131;
    exp_33_ram[1267] = 3;
    exp_33_ram[1268] = 147;
    exp_33_ram[1269] = 163;
    exp_33_ram[1270] = 147;
    exp_33_ram[1271] = 35;
    exp_33_ram[1272] = 3;
    exp_33_ram[1273] = 3;
    exp_33_ram[1274] = 19;
    exp_33_ram[1275] = 131;
    exp_33_ram[1276] = 19;
    exp_33_ram[1277] = 103;
    exp_33_ram[1278] = 19;
    exp_33_ram[1279] = 35;
    exp_33_ram[1280] = 55;
    exp_33_ram[1281] = 35;
    exp_33_ram[1282] = 35;
    exp_33_ram[1283] = 35;
    exp_33_ram[1284] = 35;
    exp_33_ram[1285] = 35;
    exp_33_ram[1286] = 35;
    exp_33_ram[1287] = 35;
    exp_33_ram[1288] = 35;
    exp_33_ram[1289] = 35;
    exp_33_ram[1290] = 35;
    exp_33_ram[1291] = 19;
    exp_33_ram[1292] = 147;
    exp_33_ram[1293] = 19;
    exp_33_ram[1294] = 147;
    exp_33_ram[1295] = 147;
    exp_33_ram[1296] = 19;
    exp_33_ram[1297] = 19;
    exp_33_ram[1298] = 239;
    exp_33_ram[1299] = 51;
    exp_33_ram[1300] = 147;
    exp_33_ram[1301] = 19;
    exp_33_ram[1302] = 239;
    exp_33_ram[1303] = 147;
    exp_33_ram[1304] = 99;
    exp_33_ram[1305] = 99;
    exp_33_ram[1306] = 179;
    exp_33_ram[1307] = 51;
    exp_33_ram[1308] = 51;
    exp_33_ram[1309] = 51;
    exp_33_ram[1310] = 147;
    exp_33_ram[1311] = 147;
    exp_33_ram[1312] = 111;
    exp_33_ram[1313] = 55;
    exp_33_ram[1314] = 147;
    exp_33_ram[1315] = 19;
    exp_33_ram[1316] = 19;
    exp_33_ram[1317] = 147;
    exp_33_ram[1318] = 19;
    exp_33_ram[1319] = 239;
    exp_33_ram[1320] = 147;
    exp_33_ram[1321] = 19;
    exp_33_ram[1322] = 147;
    exp_33_ram[1323] = 147;
    exp_33_ram[1324] = 239;
    exp_33_ram[1325] = 99;
    exp_33_ram[1326] = 99;
    exp_33_ram[1327] = 51;
    exp_33_ram[1328] = 179;
    exp_33_ram[1329] = 179;
    exp_33_ram[1330] = 51;
    exp_33_ram[1331] = 147;
    exp_33_ram[1332] = 51;
    exp_33_ram[1333] = 111;
    exp_33_ram[1334] = 183;
    exp_33_ram[1335] = 19;
    exp_33_ram[1336] = 147;
    exp_33_ram[1337] = 239;
    exp_33_ram[1338] = 35;
    exp_33_ram[1339] = 147;
    exp_33_ram[1340] = 35;
    exp_33_ram[1341] = 51;
    exp_33_ram[1342] = 3;
    exp_33_ram[1343] = 183;
    exp_33_ram[1344] = 147;
    exp_33_ram[1345] = 239;
    exp_33_ram[1346] = 35;
    exp_33_ram[1347] = 19;
    exp_33_ram[1348] = 35;
    exp_33_ram[1349] = 3;
    exp_33_ram[1350] = 147;
    exp_33_ram[1351] = 147;
    exp_33_ram[1352] = 239;
    exp_33_ram[1353] = 147;
    exp_33_ram[1354] = 35;
    exp_33_ram[1355] = 35;
    exp_33_ram[1356] = 35;
    exp_33_ram[1357] = 35;
    exp_33_ram[1358] = 35;
    exp_33_ram[1359] = 35;
    exp_33_ram[1360] = 35;
    exp_33_ram[1361] = 51;
    exp_33_ram[1362] = 35;
    exp_33_ram[1363] = 147;
    exp_33_ram[1364] = 239;
    exp_33_ram[1365] = 35;
    exp_33_ram[1366] = 35;
    exp_33_ram[1367] = 131;
    exp_33_ram[1368] = 19;
    exp_33_ram[1369] = 3;
    exp_33_ram[1370] = 131;
    exp_33_ram[1371] = 3;
    exp_33_ram[1372] = 131;
    exp_33_ram[1373] = 3;
    exp_33_ram[1374] = 131;
    exp_33_ram[1375] = 3;
    exp_33_ram[1376] = 131;
    exp_33_ram[1377] = 3;
    exp_33_ram[1378] = 131;
    exp_33_ram[1379] = 19;
    exp_33_ram[1380] = 103;
    exp_33_ram[1381] = 19;
    exp_33_ram[1382] = 35;
    exp_33_ram[1383] = 3;
    exp_33_ram[1384] = 19;
    exp_33_ram[1385] = 35;
    exp_33_ram[1386] = 35;
    exp_33_ram[1387] = 147;
    exp_33_ram[1388] = 35;
    exp_33_ram[1389] = 35;
    exp_33_ram[1390] = 19;
    exp_33_ram[1391] = 19;
    exp_33_ram[1392] = 147;
    exp_33_ram[1393] = 147;
    exp_33_ram[1394] = 19;
    exp_33_ram[1395] = 35;
    exp_33_ram[1396] = 35;
    exp_33_ram[1397] = 35;
    exp_33_ram[1398] = 35;
    exp_33_ram[1399] = 35;
    exp_33_ram[1400] = 35;
    exp_33_ram[1401] = 35;
    exp_33_ram[1402] = 35;
    exp_33_ram[1403] = 35;
    exp_33_ram[1404] = 35;
    exp_33_ram[1405] = 239;
    exp_33_ram[1406] = 19;
    exp_33_ram[1407] = 239;
    exp_33_ram[1408] = 19;
    exp_33_ram[1409] = 147;
    exp_33_ram[1410] = 19;
    exp_33_ram[1411] = 239;
    exp_33_ram[1412] = 3;
    exp_33_ram[1413] = 131;
    exp_33_ram[1414] = 19;
    exp_33_ram[1415] = 147;
    exp_33_ram[1416] = 179;
    exp_33_ram[1417] = 19;
    exp_33_ram[1418] = 35;
    exp_33_ram[1419] = 239;
    exp_33_ram[1420] = 19;
    exp_33_ram[1421] = 239;
    exp_33_ram[1422] = 19;
    exp_33_ram[1423] = 147;
    exp_33_ram[1424] = 19;
    exp_33_ram[1425] = 19;
    exp_33_ram[1426] = 147;
    exp_33_ram[1427] = 35;
    exp_33_ram[1428] = 35;
    exp_33_ram[1429] = 35;
    exp_33_ram[1430] = 35;
    exp_33_ram[1431] = 35;
    exp_33_ram[1432] = 35;
    exp_33_ram[1433] = 239;
    exp_33_ram[1434] = 19;
    exp_33_ram[1435] = 239;
    exp_33_ram[1436] = 19;
    exp_33_ram[1437] = 147;
    exp_33_ram[1438] = 19;
    exp_33_ram[1439] = 239;
    exp_33_ram[1440] = 19;
    exp_33_ram[1441] = 147;
    exp_33_ram[1442] = 19;
    exp_33_ram[1443] = 35;
    exp_33_ram[1444] = 239;
    exp_33_ram[1445] = 19;
    exp_33_ram[1446] = 239;
    exp_33_ram[1447] = 19;
    exp_33_ram[1448] = 19;
    exp_33_ram[1449] = 147;
    exp_33_ram[1450] = 19;
    exp_33_ram[1451] = 147;
    exp_33_ram[1452] = 239;
    exp_33_ram[1453] = 19;
    exp_33_ram[1454] = 239;
    exp_33_ram[1455] = 19;
    exp_33_ram[1456] = 147;
    exp_33_ram[1457] = 99;
    exp_33_ram[1458] = 99;
    exp_33_ram[1459] = 99;
    exp_33_ram[1460] = 19;
    exp_33_ram[1461] = 99;
    exp_33_ram[1462] = 99;
    exp_33_ram[1463] = 99;
    exp_33_ram[1464] = 19;
    exp_33_ram[1465] = 131;
    exp_33_ram[1466] = 3;
    exp_33_ram[1467] = 131;
    exp_33_ram[1468] = 3;
    exp_33_ram[1469] = 131;
    exp_33_ram[1470] = 3;
    exp_33_ram[1471] = 131;
    exp_33_ram[1472] = 3;
    exp_33_ram[1473] = 19;
    exp_33_ram[1474] = 103;
    exp_33_ram[1475] = 19;
    exp_33_ram[1476] = 147;
    exp_33_ram[1477] = 35;
    exp_33_ram[1478] = 19;
    exp_33_ram[1479] = 19;
    exp_33_ram[1480] = 19;
    exp_33_ram[1481] = 35;
    exp_33_ram[1482] = 35;
    exp_33_ram[1483] = 35;
    exp_33_ram[1484] = 35;
    exp_33_ram[1485] = 239;
    exp_33_ram[1486] = 19;
    exp_33_ram[1487] = 147;
    exp_33_ram[1488] = 19;
    exp_33_ram[1489] = 131;
    exp_33_ram[1490] = 239;
    exp_33_ram[1491] = 19;
    exp_33_ram[1492] = 239;
    exp_33_ram[1493] = 19;
    exp_33_ram[1494] = 147;
    exp_33_ram[1495] = 99;
    exp_33_ram[1496] = 183;
    exp_33_ram[1497] = 147;
    exp_33_ram[1498] = 179;
    exp_33_ram[1499] = 51;
    exp_33_ram[1500] = 19;
    exp_33_ram[1501] = 179;
    exp_33_ram[1502] = 147;
    exp_33_ram[1503] = 19;
    exp_33_ram[1504] = 19;
    exp_33_ram[1505] = 239;
    exp_33_ram[1506] = 19;
    exp_33_ram[1507] = 147;
    exp_33_ram[1508] = 19;
    exp_33_ram[1509] = 239;
    exp_33_ram[1510] = 99;
    exp_33_ram[1511] = 147;
    exp_33_ram[1512] = 35;
    exp_33_ram[1513] = 131;
    exp_33_ram[1514] = 19;
    exp_33_ram[1515] = 3;
    exp_33_ram[1516] = 3;
    exp_33_ram[1517] = 131;
    exp_33_ram[1518] = 147;
    exp_33_ram[1519] = 131;
    exp_33_ram[1520] = 19;
    exp_33_ram[1521] = 103;
    exp_33_ram[1522] = 227;
    exp_33_ram[1523] = 147;
    exp_33_ram[1524] = 19;
    exp_33_ram[1525] = 19;
    exp_33_ram[1526] = 239;
    exp_33_ram[1527] = 19;
    exp_33_ram[1528] = 239;
    exp_33_ram[1529] = 147;
    exp_33_ram[1530] = 51;
    exp_33_ram[1531] = 179;
    exp_33_ram[1532] = 179;
    exp_33_ram[1533] = 179;
    exp_33_ram[1534] = 179;
    exp_33_ram[1535] = 19;
    exp_33_ram[1536] = 227;
    exp_33_ram[1537] = 55;
    exp_33_ram[1538] = 19;
    exp_33_ram[1539] = 147;
    exp_33_ram[1540] = 111;
    exp_33_ram[1541] = 99;
    exp_33_ram[1542] = 19;
    exp_33_ram[1543] = 147;
    exp_33_ram[1544] = 19;
    exp_33_ram[1545] = 239;
    exp_33_ram[1546] = 19;
    exp_33_ram[1547] = 239;
    exp_33_ram[1548] = 99;
    exp_33_ram[1549] = 55;
    exp_33_ram[1550] = 19;
    exp_33_ram[1551] = 35;
    exp_33_ram[1552] = 111;
    exp_33_ram[1553] = 35;
    exp_33_ram[1554] = 111;
    exp_33_ram[1555] = 19;
    exp_33_ram[1556] = 19;
    exp_33_ram[1557] = 147;
    exp_33_ram[1558] = 19;
    exp_33_ram[1559] = 35;
    exp_33_ram[1560] = 239;
    exp_33_ram[1561] = 147;
    exp_33_ram[1562] = 19;
    exp_33_ram[1563] = 19;
    exp_33_ram[1564] = 239;
    exp_33_ram[1565] = 19;
    exp_33_ram[1566] = 239;
    exp_33_ram[1567] = 131;
    exp_33_ram[1568] = 19;
    exp_33_ram[1569] = 103;
    exp_33_ram[1570] = 19;
    exp_33_ram[1571] = 35;
    exp_33_ram[1572] = 35;
    exp_33_ram[1573] = 131;
    exp_33_ram[1574] = 3;
    exp_33_ram[1575] = 35;
    exp_33_ram[1576] = 147;
    exp_33_ram[1577] = 19;
    exp_33_ram[1578] = 35;
    exp_33_ram[1579] = 35;
    exp_33_ram[1580] = 239;
    exp_33_ram[1581] = 19;
    exp_33_ram[1582] = 99;
    exp_33_ram[1583] = 55;
    exp_33_ram[1584] = 19;
    exp_33_ram[1585] = 179;
    exp_33_ram[1586] = 51;
    exp_33_ram[1587] = 51;
    exp_33_ram[1588] = 19;
    exp_33_ram[1589] = 239;
    exp_33_ram[1590] = 55;
    exp_33_ram[1591] = 147;
    exp_33_ram[1592] = 19;
    exp_33_ram[1593] = 19;
    exp_33_ram[1594] = 239;
    exp_33_ram[1595] = 19;
    exp_33_ram[1596] = 147;
    exp_33_ram[1597] = 239;
    exp_33_ram[1598] = 147;
    exp_33_ram[1599] = 35;
    exp_33_ram[1600] = 131;
    exp_33_ram[1601] = 19;
    exp_33_ram[1602] = 3;
    exp_33_ram[1603] = 131;
    exp_33_ram[1604] = 3;
    exp_33_ram[1605] = 131;
    exp_33_ram[1606] = 19;
    exp_33_ram[1607] = 103;
    exp_33_ram[1608] = 19;
    exp_33_ram[1609] = 35;
    exp_33_ram[1610] = 35;
    exp_33_ram[1611] = 35;
    exp_33_ram[1612] = 35;
    exp_33_ram[1613] = 19;
    exp_33_ram[1614] = 35;
    exp_33_ram[1615] = 239;
    exp_33_ram[1616] = 35;
    exp_33_ram[1617] = 35;
    exp_33_ram[1618] = 19;
    exp_33_ram[1619] = 239;
    exp_33_ram[1620] = 19;
    exp_33_ram[1621] = 147;
    exp_33_ram[1622] = 3;
    exp_33_ram[1623] = 131;
    exp_33_ram[1624] = 51;
    exp_33_ram[1625] = 19;
    exp_33_ram[1626] = 51;
    exp_33_ram[1627] = 179;
    exp_33_ram[1628] = 179;
    exp_33_ram[1629] = 147;
    exp_33_ram[1630] = 131;
    exp_33_ram[1631] = 19;
    exp_33_ram[1632] = 147;
    exp_33_ram[1633] = 19;
    exp_33_ram[1634] = 147;
    exp_33_ram[1635] = 227;
    exp_33_ram[1636] = 19;
    exp_33_ram[1637] = 147;
    exp_33_ram[1638] = 99;
    exp_33_ram[1639] = 147;
    exp_33_ram[1640] = 147;
    exp_33_ram[1641] = 227;
    exp_33_ram[1642] = 19;
    exp_33_ram[1643] = 19;
    exp_33_ram[1644] = 131;
    exp_33_ram[1645] = 3;
    exp_33_ram[1646] = 3;
    exp_33_ram[1647] = 131;
    exp_33_ram[1648] = 19;
    exp_33_ram[1649] = 103;
    exp_33_ram[1650] = 19;
    exp_33_ram[1651] = 35;
    exp_33_ram[1652] = 35;
    exp_33_ram[1653] = 19;
    exp_33_ram[1654] = 19;
    exp_33_ram[1655] = 239;
    exp_33_ram[1656] = 19;
    exp_33_ram[1657] = 131;
    exp_33_ram[1658] = 3;
    exp_33_ram[1659] = 19;
    exp_33_ram[1660] = 103;
    exp_33_ram[1661] = 19;
    exp_33_ram[1662] = 35;
    exp_33_ram[1663] = 35;
    exp_33_ram[1664] = 19;
    exp_33_ram[1665] = 19;
    exp_33_ram[1666] = 239;
    exp_33_ram[1667] = 147;
    exp_33_ram[1668] = 35;
    exp_33_ram[1669] = 35;
    exp_33_ram[1670] = 111;
    exp_33_ram[1671] = 131;
    exp_33_ram[1672] = 19;
    exp_33_ram[1673] = 239;
    exp_33_ram[1674] = 111;
    exp_33_ram[1675] = 131;
    exp_33_ram[1676] = 147;
    exp_33_ram[1677] = 35;
    exp_33_ram[1678] = 183;
    exp_33_ram[1679] = 131;
    exp_33_ram[1680] = 147;
    exp_33_ram[1681] = 3;
    exp_33_ram[1682] = 239;
    exp_33_ram[1683] = 183;
    exp_33_ram[1684] = 3;
    exp_33_ram[1685] = 147;
    exp_33_ram[1686] = 179;
    exp_33_ram[1687] = 19;
    exp_33_ram[1688] = 239;
    exp_33_ram[1689] = 3;
    exp_33_ram[1690] = 147;
    exp_33_ram[1691] = 227;
    exp_33_ram[1692] = 111;
    exp_33_ram[1693] = 131;
    exp_33_ram[1694] = 147;
    exp_33_ram[1695] = 35;
    exp_33_ram[1696] = 183;
    exp_33_ram[1697] = 131;
    exp_33_ram[1698] = 147;
    exp_33_ram[1699] = 3;
    exp_33_ram[1700] = 239;
    exp_33_ram[1701] = 183;
    exp_33_ram[1702] = 3;
    exp_33_ram[1703] = 147;
    exp_33_ram[1704] = 179;
    exp_33_ram[1705] = 19;
    exp_33_ram[1706] = 239;
    exp_33_ram[1707] = 3;
    exp_33_ram[1708] = 147;
    exp_33_ram[1709] = 227;
    exp_33_ram[1710] = 131;
    exp_33_ram[1711] = 147;
    exp_33_ram[1712] = 35;
    exp_33_ram[1713] = 3;
    exp_33_ram[1714] = 147;
    exp_33_ram[1715] = 227;
    exp_33_ram[1716] = 183;
    exp_33_ram[1717] = 131;
    exp_33_ram[1718] = 147;
    exp_33_ram[1719] = 19;
    exp_33_ram[1720] = 239;
    exp_33_ram[1721] = 19;
    exp_33_ram[1722] = 131;
    exp_33_ram[1723] = 3;
    exp_33_ram[1724] = 19;
    exp_33_ram[1725] = 103;
    exp_33_ram[1726] = 19;
    exp_33_ram[1727] = 35;
    exp_33_ram[1728] = 35;
    exp_33_ram[1729] = 19;
    exp_33_ram[1730] = 131;
    exp_33_ram[1731] = 19;
    exp_33_ram[1732] = 35;
    exp_33_ram[1733] = 131;
    exp_33_ram[1734] = 19;
    exp_33_ram[1735] = 35;
    exp_33_ram[1736] = 131;
    exp_33_ram[1737] = 19;
    exp_33_ram[1738] = 35;
    exp_33_ram[1739] = 131;
    exp_33_ram[1740] = 19;
    exp_33_ram[1741] = 35;
    exp_33_ram[1742] = 131;
    exp_33_ram[1743] = 19;
    exp_33_ram[1744] = 35;
    exp_33_ram[1745] = 131;
    exp_33_ram[1746] = 35;
    exp_33_ram[1747] = 131;
    exp_33_ram[1748] = 19;
    exp_33_ram[1749] = 35;
    exp_33_ram[1750] = 3;
    exp_33_ram[1751] = 239;
    exp_33_ram[1752] = 19;
    exp_33_ram[1753] = 147;
    exp_33_ram[1754] = 19;
    exp_33_ram[1755] = 147;
    exp_33_ram[1756] = 239;
    exp_33_ram[1757] = 19;
    exp_33_ram[1758] = 239;
    exp_33_ram[1759] = 19;
    exp_33_ram[1760] = 147;
    exp_33_ram[1761] = 35;
    exp_33_ram[1762] = 35;
    exp_33_ram[1763] = 147;
    exp_33_ram[1764] = 19;
    exp_33_ram[1765] = 239;
    exp_33_ram[1766] = 35;
    exp_33_ram[1767] = 3;
    exp_33_ram[1768] = 239;
    exp_33_ram[1769] = 147;
    exp_33_ram[1770] = 19;
    exp_33_ram[1771] = 239;
    exp_33_ram[1772] = 183;
    exp_33_ram[1773] = 131;
    exp_33_ram[1774] = 19;
    exp_33_ram[1775] = 239;
    exp_33_ram[1776] = 111;
    exp_33_ram[1777] = 19;
    exp_33_ram[1778] = 35;
    exp_33_ram[1779] = 35;
    exp_33_ram[1780] = 35;
    exp_33_ram[1781] = 35;
    exp_33_ram[1782] = 35;
    exp_33_ram[1783] = 35;
    exp_33_ram[1784] = 35;
    exp_33_ram[1785] = 35;
    exp_33_ram[1786] = 35;
    exp_33_ram[1787] = 35;
    exp_33_ram[1788] = 35;
    exp_33_ram[1789] = 35;
    exp_33_ram[1790] = 19;
    exp_33_ram[1791] = 147;
    exp_33_ram[1792] = 35;
    exp_33_ram[1793] = 19;
    exp_33_ram[1794] = 147;
    exp_33_ram[1795] = 35;
    exp_33_ram[1796] = 35;
    exp_33_ram[1797] = 239;
    exp_33_ram[1798] = 35;
    exp_33_ram[1799] = 35;
    exp_33_ram[1800] = 35;
    exp_33_ram[1801] = 111;
    exp_33_ram[1802] = 3;
    exp_33_ram[1803] = 183;
    exp_33_ram[1804] = 147;
    exp_33_ram[1805] = 179;
    exp_33_ram[1806] = 35;
    exp_33_ram[1807] = 3;
    exp_33_ram[1808] = 183;
    exp_33_ram[1809] = 147;
    exp_33_ram[1810] = 179;
    exp_33_ram[1811] = 35;
    exp_33_ram[1812] = 3;
    exp_33_ram[1813] = 183;
    exp_33_ram[1814] = 147;
    exp_33_ram[1815] = 179;
    exp_33_ram[1816] = 35;
    exp_33_ram[1817] = 3;
    exp_33_ram[1818] = 183;
    exp_33_ram[1819] = 147;
    exp_33_ram[1820] = 179;
    exp_33_ram[1821] = 35;
    exp_33_ram[1822] = 131;
    exp_33_ram[1823] = 147;
    exp_33_ram[1824] = 35;
    exp_33_ram[1825] = 239;
    exp_33_ram[1826] = 19;
    exp_33_ram[1827] = 147;
    exp_33_ram[1828] = 3;
    exp_33_ram[1829] = 131;
    exp_33_ram[1830] = 51;
    exp_33_ram[1831] = 19;
    exp_33_ram[1832] = 51;
    exp_33_ram[1833] = 179;
    exp_33_ram[1834] = 179;
    exp_33_ram[1835] = 147;
    exp_33_ram[1836] = 183;
    exp_33_ram[1837] = 131;
    exp_33_ram[1838] = 35;
    exp_33_ram[1839] = 35;
    exp_33_ram[1840] = 3;
    exp_33_ram[1841] = 131;
    exp_33_ram[1842] = 19;
    exp_33_ram[1843] = 147;
    exp_33_ram[1844] = 227;
    exp_33_ram[1845] = 19;
    exp_33_ram[1846] = 147;
    exp_33_ram[1847] = 99;
    exp_33_ram[1848] = 147;
    exp_33_ram[1849] = 147;
    exp_33_ram[1850] = 227;
    exp_33_ram[1851] = 131;
    exp_33_ram[1852] = 19;
    exp_33_ram[1853] = 239;
    exp_33_ram[1854] = 239;
    exp_33_ram[1855] = 35;
    exp_33_ram[1856] = 35;
    exp_33_ram[1857] = 35;
    exp_33_ram[1858] = 111;
    exp_33_ram[1859] = 3;
    exp_33_ram[1860] = 131;
    exp_33_ram[1861] = 183;
    exp_33_ram[1862] = 147;
    exp_33_ram[1863] = 51;
    exp_33_ram[1864] = 147;
    exp_33_ram[1865] = 179;
    exp_33_ram[1866] = 51;
    exp_33_ram[1867] = 183;
    exp_33_ram[1868] = 147;
    exp_33_ram[1869] = 179;
    exp_33_ram[1870] = 179;
    exp_33_ram[1871] = 19;
    exp_33_ram[1872] = 179;
    exp_33_ram[1873] = 147;
    exp_33_ram[1874] = 35;
    exp_33_ram[1875] = 35;
    exp_33_ram[1876] = 3;
    exp_33_ram[1877] = 131;
    exp_33_ram[1878] = 183;
    exp_33_ram[1879] = 147;
    exp_33_ram[1880] = 51;
    exp_33_ram[1881] = 147;
    exp_33_ram[1882] = 179;
    exp_33_ram[1883] = 51;
    exp_33_ram[1884] = 183;
    exp_33_ram[1885] = 147;
    exp_33_ram[1886] = 179;
    exp_33_ram[1887] = 179;
    exp_33_ram[1888] = 19;
    exp_33_ram[1889] = 179;
    exp_33_ram[1890] = 147;
    exp_33_ram[1891] = 35;
    exp_33_ram[1892] = 35;
    exp_33_ram[1893] = 3;
    exp_33_ram[1894] = 131;
    exp_33_ram[1895] = 183;
    exp_33_ram[1896] = 147;
    exp_33_ram[1897] = 51;
    exp_33_ram[1898] = 147;
    exp_33_ram[1899] = 179;
    exp_33_ram[1900] = 51;
    exp_33_ram[1901] = 183;
    exp_33_ram[1902] = 147;
    exp_33_ram[1903] = 179;
    exp_33_ram[1904] = 179;
    exp_33_ram[1905] = 19;
    exp_33_ram[1906] = 179;
    exp_33_ram[1907] = 147;
    exp_33_ram[1908] = 35;
    exp_33_ram[1909] = 35;
    exp_33_ram[1910] = 3;
    exp_33_ram[1911] = 131;
    exp_33_ram[1912] = 183;
    exp_33_ram[1913] = 147;
    exp_33_ram[1914] = 51;
    exp_33_ram[1915] = 147;
    exp_33_ram[1916] = 179;
    exp_33_ram[1917] = 51;
    exp_33_ram[1918] = 183;
    exp_33_ram[1919] = 147;
    exp_33_ram[1920] = 179;
    exp_33_ram[1921] = 179;
    exp_33_ram[1922] = 19;
    exp_33_ram[1923] = 179;
    exp_33_ram[1924] = 147;
    exp_33_ram[1925] = 35;
    exp_33_ram[1926] = 35;
    exp_33_ram[1927] = 131;
    exp_33_ram[1928] = 147;
    exp_33_ram[1929] = 35;
    exp_33_ram[1930] = 239;
    exp_33_ram[1931] = 19;
    exp_33_ram[1932] = 147;
    exp_33_ram[1933] = 3;
    exp_33_ram[1934] = 131;
    exp_33_ram[1935] = 51;
    exp_33_ram[1936] = 19;
    exp_33_ram[1937] = 51;
    exp_33_ram[1938] = 179;
    exp_33_ram[1939] = 179;
    exp_33_ram[1940] = 147;
    exp_33_ram[1941] = 183;
    exp_33_ram[1942] = 131;
    exp_33_ram[1943] = 35;
    exp_33_ram[1944] = 35;
    exp_33_ram[1945] = 3;
    exp_33_ram[1946] = 131;
    exp_33_ram[1947] = 19;
    exp_33_ram[1948] = 147;
    exp_33_ram[1949] = 227;
    exp_33_ram[1950] = 19;
    exp_33_ram[1951] = 147;
    exp_33_ram[1952] = 99;
    exp_33_ram[1953] = 147;
    exp_33_ram[1954] = 147;
    exp_33_ram[1955] = 227;
    exp_33_ram[1956] = 131;
    exp_33_ram[1957] = 19;
    exp_33_ram[1958] = 239;
    exp_33_ram[1959] = 239;
    exp_33_ram[1960] = 35;
    exp_33_ram[1961] = 35;
    exp_33_ram[1962] = 35;
    exp_33_ram[1963] = 111;
    exp_33_ram[1964] = 3;
    exp_33_ram[1965] = 183;
    exp_33_ram[1966] = 147;
    exp_33_ram[1967] = 179;
    exp_33_ram[1968] = 35;
    exp_33_ram[1969] = 3;
    exp_33_ram[1970] = 183;
    exp_33_ram[1971] = 147;
    exp_33_ram[1972] = 179;
    exp_33_ram[1973] = 35;
    exp_33_ram[1974] = 3;
    exp_33_ram[1975] = 183;
    exp_33_ram[1976] = 147;
    exp_33_ram[1977] = 179;
    exp_33_ram[1978] = 35;
    exp_33_ram[1979] = 3;
    exp_33_ram[1980] = 183;
    exp_33_ram[1981] = 147;
    exp_33_ram[1982] = 179;
    exp_33_ram[1983] = 35;
    exp_33_ram[1984] = 131;
    exp_33_ram[1985] = 147;
    exp_33_ram[1986] = 35;
    exp_33_ram[1987] = 239;
    exp_33_ram[1988] = 19;
    exp_33_ram[1989] = 147;
    exp_33_ram[1990] = 3;
    exp_33_ram[1991] = 131;
    exp_33_ram[1992] = 51;
    exp_33_ram[1993] = 19;
    exp_33_ram[1994] = 51;
    exp_33_ram[1995] = 179;
    exp_33_ram[1996] = 179;
    exp_33_ram[1997] = 147;
    exp_33_ram[1998] = 183;
    exp_33_ram[1999] = 131;
    exp_33_ram[2000] = 35;
    exp_33_ram[2001] = 35;
    exp_33_ram[2002] = 3;
    exp_33_ram[2003] = 131;
    exp_33_ram[2004] = 19;
    exp_33_ram[2005] = 147;
    exp_33_ram[2006] = 227;
    exp_33_ram[2007] = 19;
    exp_33_ram[2008] = 147;
    exp_33_ram[2009] = 99;
    exp_33_ram[2010] = 147;
    exp_33_ram[2011] = 147;
    exp_33_ram[2012] = 227;
    exp_33_ram[2013] = 131;
    exp_33_ram[2014] = 19;
    exp_33_ram[2015] = 239;
    exp_33_ram[2016] = 239;
    exp_33_ram[2017] = 35;
    exp_33_ram[2018] = 35;
    exp_33_ram[2019] = 35;
    exp_33_ram[2020] = 111;
    exp_33_ram[2021] = 3;
    exp_33_ram[2022] = 131;
    exp_33_ram[2023] = 55;
    exp_33_ram[2024] = 19;
    exp_33_ram[2025] = 147;
    exp_33_ram[2026] = 19;
    exp_33_ram[2027] = 147;
    exp_33_ram[2028] = 239;
    exp_33_ram[2029] = 19;
    exp_33_ram[2030] = 147;
    exp_33_ram[2031] = 35;
    exp_33_ram[2032] = 35;
    exp_33_ram[2033] = 3;
    exp_33_ram[2034] = 131;
    exp_33_ram[2035] = 55;
    exp_33_ram[2036] = 19;
    exp_33_ram[2037] = 147;
    exp_33_ram[2038] = 19;
    exp_33_ram[2039] = 147;
    exp_33_ram[2040] = 239;
    exp_33_ram[2041] = 19;
    exp_33_ram[2042] = 147;
    exp_33_ram[2043] = 35;
    exp_33_ram[2044] = 35;
    exp_33_ram[2045] = 3;
    exp_33_ram[2046] = 131;
    exp_33_ram[2047] = 55;
    exp_33_ram[2048] = 19;
    exp_33_ram[2049] = 147;
    exp_33_ram[2050] = 19;
    exp_33_ram[2051] = 147;
    exp_33_ram[2052] = 239;
    exp_33_ram[2053] = 19;
    exp_33_ram[2054] = 147;
    exp_33_ram[2055] = 35;
    exp_33_ram[2056] = 35;
    exp_33_ram[2057] = 3;
    exp_33_ram[2058] = 131;
    exp_33_ram[2059] = 55;
    exp_33_ram[2060] = 19;
    exp_33_ram[2061] = 147;
    exp_33_ram[2062] = 19;
    exp_33_ram[2063] = 147;
    exp_33_ram[2064] = 239;
    exp_33_ram[2065] = 19;
    exp_33_ram[2066] = 147;
    exp_33_ram[2067] = 35;
    exp_33_ram[2068] = 35;
    exp_33_ram[2069] = 131;
    exp_33_ram[2070] = 147;
    exp_33_ram[2071] = 35;
    exp_33_ram[2072] = 239;
    exp_33_ram[2073] = 19;
    exp_33_ram[2074] = 147;
    exp_33_ram[2075] = 3;
    exp_33_ram[2076] = 131;
    exp_33_ram[2077] = 51;
    exp_33_ram[2078] = 19;
    exp_33_ram[2079] = 51;
    exp_33_ram[2080] = 179;
    exp_33_ram[2081] = 179;
    exp_33_ram[2082] = 147;
    exp_33_ram[2083] = 183;
    exp_33_ram[2084] = 131;
    exp_33_ram[2085] = 19;
    exp_33_ram[2086] = 147;
    exp_33_ram[2087] = 19;
    exp_33_ram[2088] = 147;
    exp_33_ram[2089] = 227;
    exp_33_ram[2090] = 19;
    exp_33_ram[2091] = 147;
    exp_33_ram[2092] = 99;
    exp_33_ram[2093] = 147;
    exp_33_ram[2094] = 147;
    exp_33_ram[2095] = 227;
    exp_33_ram[2096] = 131;
    exp_33_ram[2097] = 19;
    exp_33_ram[2098] = 239;
    exp_33_ram[2099] = 19;
    exp_33_ram[2100] = 131;
    exp_33_ram[2101] = 3;
    exp_33_ram[2102] = 3;
    exp_33_ram[2103] = 131;
    exp_33_ram[2104] = 3;
    exp_33_ram[2105] = 131;
    exp_33_ram[2106] = 3;
    exp_33_ram[2107] = 131;
    exp_33_ram[2108] = 3;
    exp_33_ram[2109] = 131;
    exp_33_ram[2110] = 3;
    exp_33_ram[2111] = 131;
    exp_33_ram[2112] = 19;
    exp_33_ram[2113] = 103;
    exp_33_ram[2114] = 19;
    exp_33_ram[2115] = 35;
    exp_33_ram[2116] = 35;
    exp_33_ram[2117] = 19;
    exp_33_ram[2118] = 35;
    exp_33_ram[2119] = 111;
    exp_33_ram[2120] = 131;
    exp_33_ram[2121] = 19;
    exp_33_ram[2122] = 131;
    exp_33_ram[2123] = 147;
    exp_33_ram[2124] = 179;
    exp_33_ram[2125] = 35;
    exp_33_ram[2126] = 131;
    exp_33_ram[2127] = 147;
    exp_33_ram[2128] = 35;
    exp_33_ram[2129] = 3;
    exp_33_ram[2130] = 147;
    exp_33_ram[2131] = 227;
    exp_33_ram[2132] = 35;
    exp_33_ram[2133] = 111;
    exp_33_ram[2134] = 131;
    exp_33_ram[2135] = 19;
    exp_33_ram[2136] = 239;
    exp_33_ram[2137] = 131;
    exp_33_ram[2138] = 19;
    exp_33_ram[2139] = 179;
    exp_33_ram[2140] = 19;
    exp_33_ram[2141] = 131;
    exp_33_ram[2142] = 179;
    exp_33_ram[2143] = 19;
    exp_33_ram[2144] = 147;
    exp_33_ram[2145] = 19;
    exp_33_ram[2146] = 147;
    exp_33_ram[2147] = 19;
    exp_33_ram[2148] = 239;
    exp_33_ram[2149] = 131;
    exp_33_ram[2150] = 35;
    exp_33_ram[2151] = 111;
    exp_33_ram[2152] = 131;
    exp_33_ram[2153] = 19;
    exp_33_ram[2154] = 179;
    exp_33_ram[2155] = 131;
    exp_33_ram[2156] = 19;
    exp_33_ram[2157] = 131;
    exp_33_ram[2158] = 147;
    exp_33_ram[2159] = 179;
    exp_33_ram[2160] = 131;
    exp_33_ram[2161] = 147;
    exp_33_ram[2162] = 131;
    exp_33_ram[2163] = 179;
    exp_33_ram[2164] = 99;
    exp_33_ram[2165] = 19;
    exp_33_ram[2166] = 239;
    exp_33_ram[2167] = 111;
    exp_33_ram[2168] = 131;
    exp_33_ram[2169] = 147;
    exp_33_ram[2170] = 35;
    exp_33_ram[2171] = 3;
    exp_33_ram[2172] = 147;
    exp_33_ram[2173] = 227;
    exp_33_ram[2174] = 19;
    exp_33_ram[2175] = 239;
    exp_33_ram[2176] = 131;
    exp_33_ram[2177] = 147;
    exp_33_ram[2178] = 35;
    exp_33_ram[2179] = 3;
    exp_33_ram[2180] = 147;
    exp_33_ram[2181] = 227;
    exp_33_ram[2182] = 19;
    exp_33_ram[2183] = 239;
    exp_33_ram[2184] = 147;
    exp_33_ram[2185] = 35;
    exp_33_ram[2186] = 19;
    exp_33_ram[2187] = 239;
    exp_33_ram[2188] = 147;
    exp_33_ram[2189] = 35;
    exp_33_ram[2190] = 19;
    exp_33_ram[2191] = 239;
    exp_33_ram[2192] = 147;
    exp_33_ram[2193] = 35;
    exp_33_ram[2194] = 35;
    exp_33_ram[2195] = 111;
    exp_33_ram[2196] = 3;
    exp_33_ram[2197] = 239;
    exp_33_ram[2198] = 19;
    exp_33_ram[2199] = 239;
    exp_33_ram[2200] = 147;
    exp_33_ram[2201] = 35;
    exp_33_ram[2202] = 3;
    exp_33_ram[2203] = 239;
    exp_33_ram[2204] = 19;
    exp_33_ram[2205] = 239;
    exp_33_ram[2206] = 147;
    exp_33_ram[2207] = 35;
    exp_33_ram[2208] = 3;
    exp_33_ram[2209] = 239;
    exp_33_ram[2210] = 19;
    exp_33_ram[2211] = 239;
    exp_33_ram[2212] = 147;
    exp_33_ram[2213] = 35;
    exp_33_ram[2214] = 131;
    exp_33_ram[2215] = 3;
    exp_33_ram[2216] = 131;
    exp_33_ram[2217] = 19;
    exp_33_ram[2218] = 147;
    exp_33_ram[2219] = 19;
    exp_33_ram[2220] = 239;
    exp_33_ram[2221] = 131;
    exp_33_ram[2222] = 147;
    exp_33_ram[2223] = 35;
    exp_33_ram[2224] = 3;
    exp_33_ram[2225] = 147;
    exp_33_ram[2226] = 227;
    exp_33_ram[2227] = 3;
    exp_33_ram[2228] = 239;
    exp_33_ram[2229] = 3;
    exp_33_ram[2230] = 239;
    exp_33_ram[2231] = 3;
    exp_33_ram[2232] = 239;
    exp_33_ram[2233] = 131;
    exp_33_ram[2234] = 3;
    exp_33_ram[2235] = 19;
    exp_33_ram[2236] = 103;
    exp_33_ram[2237] = 19;
    exp_33_ram[2238] = 35;
    exp_33_ram[2239] = 35;
    exp_33_ram[2240] = 19;
    exp_33_ram[2241] = 19;
    exp_33_ram[2242] = 239;
    exp_33_ram[2243] = 19;
    exp_33_ram[2244] = 239;
    exp_33_ram[2245] = 19;
    exp_33_ram[2246] = 239;
    exp_33_ram[2247] = 19;
    exp_33_ram[2248] = 239;
    exp_33_ram[2249] = 19;
    exp_33_ram[2250] = 239;
    exp_33_ram[2251] = 19;
    exp_33_ram[2252] = 239;
    exp_33_ram[2253] = 239;
    exp_33_ram[2254] = 147;
    exp_33_ram[2255] = 163;
    exp_33_ram[2256] = 131;
    exp_33_ram[2257] = 147;
    exp_33_ram[2258] = 19;
    exp_33_ram[2259] = 227;
    exp_33_ram[2260] = 19;
    exp_33_ram[2261] = 183;
    exp_33_ram[2262] = 147;
    exp_33_ram[2263] = 179;
    exp_33_ram[2264] = 131;
    exp_33_ram[2265] = 103;
    exp_33_ram[2266] = 239;
    exp_33_ram[2267] = 111;
    exp_33_ram[2268] = 239;
    exp_33_ram[2269] = 111;
    exp_33_ram[2270] = 239;
    exp_33_ram[2271] = 111;
    exp_33_ram[2272] = 239;
    exp_33_ram[2273] = 111;
    exp_33_ram[2274] = 239;
    exp_33_ram[2275] = 19;
    exp_33_ram[2276] = 111;
    exp_33_ram[2277] = 19;
    exp_33_ram[2278] = 147;
    exp_33_ram[2279] = 51;
    exp_33_ram[2280] = 19;
    exp_33_ram[2281] = 179;
    exp_33_ram[2282] = 99;
    exp_33_ram[2283] = 99;
    exp_33_ram[2284] = 19;
    exp_33_ram[2285] = 179;
    exp_33_ram[2286] = 19;
    exp_33_ram[2287] = 103;
    exp_33_ram[2288] = 227;
    exp_33_ram[2289] = 19;
    exp_33_ram[2290] = 179;
    exp_33_ram[2291] = 111;
    exp_33_ram[2292] = 128;
    exp_33_ram[2293] = 0;
    exp_33_ram[2294] = 8;
    exp_33_ram[2295] = 12;
    exp_33_ram[2296] = 16;
    exp_33_ram[2297] = 83;
    exp_33_ram[2298] = 111;
    exp_33_ram[2299] = 101;
    exp_33_ram[2300] = 84;
    exp_33_ram[2301] = 114;
    exp_33_ram[2302] = 116;
    exp_33_ram[2303] = 74;
    exp_33_ram[2304] = 101;
    exp_33_ram[2305] = 114;
    exp_33_ram[2306] = 77;
    exp_33_ram[2307] = 117;
    exp_33_ram[2308] = 108;
    exp_33_ram[2309] = 83;
    exp_33_ram[2310] = 99;
    exp_33_ram[2311] = 118;
    exp_33_ram[2312] = 0;
    exp_33_ram[2313] = 104;
    exp_33_ram[2314] = 112;
    exp_33_ram[2315] = 120;
    exp_33_ram[2316] = 128;
    exp_33_ram[2317] = 136;
    exp_33_ram[2318] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_179;

  reg [31:0] exp_179_reg;
  always@(*) begin
    case (exp_177)
      0:exp_179_reg <= exp_157;
      1:exp_179_reg <= exp_167;
      default:exp_179_reg <= exp_178;
    endcase
  end
  assign exp_179 = exp_179_reg;
  assign exp_177 = exp_139[2:2];
  assign exp_139 = exp_1;
  assign exp_178 = 0;

      reg [31:0] exp_157_reg = 0;
      always@(posedge clk) begin
        if (exp_156) begin
          exp_157_reg <= exp_164;
        end
      end
      assign exp_157 = exp_157_reg;
    
  reg [31:0] exp_164_reg;
  always@(*) begin
    case (exp_159)
      0:exp_164_reg <= exp_161;
      1:exp_164_reg <= exp_162;
      default:exp_164_reg <= exp_163;
    endcase
  end
  assign exp_164 = exp_164_reg;
  assign exp_159 = exp_157 == exp_158;
  assign exp_158 = 4294967295;
  assign exp_163 = 0;
  assign exp_161 = exp_157 + exp_160;
  assign exp_160 = 1;
  assign exp_162 = 0;
  assign exp_156 = 1;

      reg [31:0] exp_167_reg = 0;
      always@(posedge clk) begin
        if (exp_166) begin
          exp_167_reg <= exp_174;
        end
      end
      assign exp_167 = exp_167_reg;
    
  reg [31:0] exp_174_reg;
  always@(*) begin
    case (exp_169)
      0:exp_174_reg <= exp_171;
      1:exp_174_reg <= exp_172;
      default:exp_174_reg <= exp_173;
    endcase
  end
  assign exp_174 = exp_174_reg;
  assign exp_169 = exp_167 == exp_168;
  assign exp_168 = 4294967295;
  assign exp_173 = 0;
  assign exp_171 = exp_167 + exp_170;
  assign exp_170 = 1;
  assign exp_172 = 0;
  assign exp_166 = exp_159 & exp_165;
  assign exp_165 = 1;
  assign exp_182 = exp_201;
  assign exp_201 = 0;
  assign exp_204 = exp_222;
  assign exp_222 = 0;
  assign exp_226 = exp_241;
  assign exp_241 = stdin_in;
  assign exp_461 = exp_248[15:8];
  assign exp_462 = exp_248[23:16];
  assign exp_463 = exp_248[31:24];
  assign exp_475 = $signed(exp_474);
  assign exp_474 = exp_473 + exp_469;
  assign exp_473 = 0;

  reg [15:0] exp_469_reg;
  always@(*) begin
    case (exp_459)
      0:exp_469_reg <= exp_466;
      1:exp_469_reg <= exp_467;
      default:exp_469_reg <= exp_468;
    endcase
  end
  assign exp_469 = exp_469_reg;
  assign exp_468 = 0;
  assign exp_466 = exp_248[15:0];
  assign exp_467 = exp_248[31:16];
  assign exp_476 = 0;
  assign exp_477 = exp_465;
  assign exp_478 = exp_469;
  assign exp_479 = 0;
  assign exp_480 = 0;

  reg [31:0] exp_839_reg;
  always@(*) begin
    case (exp_629)
      0:exp_839_reg <= exp_835;
      1:exp_839_reg <= exp_837;
      default:exp_839_reg <= exp_838;
    endcase
  end
  assign exp_839 = exp_839_reg;
  assign exp_838 = 0;

  reg [31:0] exp_835_reg;
  always@(*) begin
    case (exp_606)
      0:exp_835_reg <= exp_830;
      1:exp_835_reg <= exp_831;
      default:exp_835_reg <= exp_834;
    endcase
  end
  assign exp_835 = exp_835_reg;
  assign exp_606 = exp_605 & exp_603;
  assign exp_605 = exp_598 == exp_604;
  assign exp_604 = 0;
  assign exp_834 = 0;
  assign exp_830 = exp_829[63:32];

  reg [63:0] exp_829_reg;
  always@(*) begin
    case (exp_826)
      0:exp_829_reg <= exp_825;
      1:exp_829_reg <= exp_827;
      default:exp_829_reg <= exp_828;
    endcase
  end
  assign exp_829 = exp_829_reg;

      reg [0:0] exp_826_reg = 0;
      always@(posedge clk) begin
        if (exp_811) begin
          exp_826_reg <= exp_809;
        end
      end
      assign exp_826 = exp_826_reg;
    
      reg [0:0] exp_809_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_809_reg <= exp_786;
        end
      end
      assign exp_809 = exp_809_reg;
    
      reg [0:0] exp_786_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_786_reg <= exp_783;
        end
      end
      assign exp_786 = exp_786_reg;
      assign exp_783 = exp_781 ^ exp_782;
  assign exp_781 = exp_763 & exp_746;
  assign exp_763 = exp_762 + exp_761;
  assign exp_762 = 0;
  assign exp_761 = exp_759[31:31];

      reg [31:0] exp_759_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_759_reg <= exp_376;
        end
      end
      assign exp_759 = exp_759_reg;
      assign exp_758 = exp_748 == exp_757;
  assign exp_757 = 0;
  assign exp_746 = exp_745 | exp_612;
  assign exp_745 = exp_606 | exp_609;
  assign exp_609 = exp_608 & exp_603;
  assign exp_608 = exp_598 == exp_607;
  assign exp_607 = 1;
  assign exp_612 = exp_611 & exp_603;
  assign exp_611 = exp_598 == exp_610;
  assign exp_610 = 2;
  assign exp_782 = exp_766 & exp_747;
  assign exp_766 = exp_765 + exp_764;
  assign exp_765 = 0;
  assign exp_764 = exp_760[31:31];

      reg [31:0] exp_760_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_760_reg <= exp_377;
        end
      end
      assign exp_760 = exp_760_reg;
      assign exp_747 = exp_606 | exp_609;
  assign exp_768 = exp_748 == exp_767;
  assign exp_767 = 1;
  assign exp_788 = exp_748 == exp_787;
  assign exp_787 = 2;
  assign exp_811 = exp_748 == exp_810;
  assign exp_810 = 3;
  assign exp_828 = 0;

      reg [63:0] exp_825_reg = 0;
      always@(posedge clk) begin
        if (exp_811) begin
          exp_825_reg <= exp_824;
        end
      end
      assign exp_825 = exp_825_reg;
      assign exp_824 = exp_820 + exp_823;
  assign exp_820 = exp_816 + exp_819;
  assign exp_816 = exp_812 + exp_815;
  assign exp_812 = exp_805;

      reg [31:0] exp_805_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_805_reg <= exp_792;
        end
      end
      assign exp_805 = exp_805_reg;
      assign exp_792 = exp_790 * exp_791;
  assign exp_790 = exp_789;
  assign exp_789 = exp_784[15:0];

      reg [31:0] exp_784_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_784_reg <= exp_774;
        end
      end
      assign exp_784 = exp_784_reg;
      assign exp_774 = exp_773 + exp_772;
  assign exp_773 = 0;

  reg [31:0] exp_772_reg;
  always@(*) begin
    case (exp_769)
      0:exp_772_reg <= exp_759;
      1:exp_772_reg <= exp_770;
      default:exp_772_reg <= exp_771;
    endcase
  end
  assign exp_772 = exp_772_reg;
  assign exp_769 = exp_763 & exp_746;
  assign exp_771 = 0;
  assign exp_770 = -exp_759;
  assign exp_791 = exp_785[15:0];

      reg [31:0] exp_785_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_785_reg <= exp_780;
        end
      end
      assign exp_785 = exp_785_reg;
      assign exp_780 = exp_779 + exp_778;
  assign exp_779 = 0;

  reg [31:0] exp_778_reg;
  always@(*) begin
    case (exp_775)
      0:exp_778_reg <= exp_760;
      1:exp_778_reg <= exp_776;
      default:exp_778_reg <= exp_777;
    endcase
  end
  assign exp_778 = exp_778_reg;
  assign exp_775 = exp_766 & exp_747;
  assign exp_777 = 0;
  assign exp_776 = -exp_760;
  assign exp_815 = exp_813 << exp_814;
  assign exp_813 = exp_806;

      reg [31:0] exp_806_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_806_reg <= exp_796;
        end
      end
      assign exp_806 = exp_806_reg;
      assign exp_796 = exp_794 * exp_795;
  assign exp_794 = exp_793;
  assign exp_793 = exp_784[15:0];
  assign exp_795 = exp_785[31:16];
  assign exp_814 = 16;
  assign exp_819 = exp_817 << exp_818;
  assign exp_817 = exp_807;

      reg [31:0] exp_807_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_807_reg <= exp_800;
        end
      end
      assign exp_807 = exp_807_reg;
      assign exp_800 = exp_798 * exp_799;
  assign exp_798 = exp_797;
  assign exp_797 = exp_784[31:16];
  assign exp_799 = exp_785[15:0];
  assign exp_818 = 16;
  assign exp_823 = exp_821 << exp_822;
  assign exp_821 = exp_808;

      reg [31:0] exp_808_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_808_reg <= exp_804;
        end
      end
      assign exp_808 = exp_808_reg;
      assign exp_804 = exp_802 * exp_803;
  assign exp_802 = exp_801;
  assign exp_801 = exp_784[31:16];
  assign exp_803 = exp_785[31:16];
  assign exp_822 = 32;
  assign exp_827 = -exp_825;
  assign exp_831 = exp_829[31:0];

  reg [31:0] exp_837_reg;
  always@(*) begin
    case (exp_630)
      0:exp_837_reg <= exp_740;
      1:exp_837_reg <= exp_741;
      default:exp_837_reg <= exp_836;
    endcase
  end
  assign exp_837 = exp_837_reg;
  assign exp_630 = exp_598[1:1];
  assign exp_836 = 0;

      reg [31:0] exp_740_reg = 0;
      always@(posedge clk) begin
        if (exp_649) begin
          exp_740_reg <= exp_734;
        end
      end
      assign exp_740 = exp_740_reg;
    
  reg [31:0] exp_734_reg;
  always@(*) begin
    case (exp_730)
      0:exp_734_reg <= exp_721;
      1:exp_734_reg <= exp_732;
      default:exp_734_reg <= exp_733;
    endcase
  end
  assign exp_734 = exp_734_reg;
  assign exp_730 = exp_729 & exp_632;
  assign exp_729 = exp_678 == exp_728;

      reg [31:0] exp_678_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_678_reg <= exp_675;
        end
      end
      assign exp_678 = exp_678_reg;
      assign exp_675 = exp_674 + exp_673;
  assign exp_674 = 0;

  reg [31:0] exp_673_reg;
  always@(*) begin
    case (exp_670)
      0:exp_673_reg <= exp_655;
      1:exp_673_reg <= exp_671;
      default:exp_673_reg <= exp_672;
    endcase
  end
  assign exp_673 = exp_673_reg;
  assign exp_670 = exp_661 & exp_632;
  assign exp_661 = exp_660 + exp_659;
  assign exp_660 = 0;
  assign exp_659 = exp_655[31:31];

      reg [31:0] exp_655_reg = 0;
      always@(posedge clk) begin
        if (exp_653) begin
          exp_655_reg <= exp_377;
        end
      end
      assign exp_655 = exp_655_reg;
      assign exp_653 = exp_635 == exp_652;
  assign exp_652 = 0;
  assign exp_632 = ~exp_631;
  assign exp_631 = exp_598[0:0];
  assign exp_672 = 0;
  assign exp_671 = -exp_655;
  assign exp_663 = exp_635 == exp_662;
  assign exp_662 = 1;
  assign exp_728 = 0;
  assign exp_733 = 0;
  assign exp_721 = exp_720 + exp_719;
  assign exp_720 = 0;

  reg [31:0] exp_719_reg;
  always@(*) begin
    case (exp_716)
      0:exp_719_reg <= exp_714;
      1:exp_719_reg <= exp_717;
      default:exp_719_reg <= exp_718;
    endcase
  end
  assign exp_719 = exp_719_reg;
  assign exp_716 = exp_680 & exp_632;

      reg [0:0] exp_680_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_680_reg <= exp_676;
        end
      end
      assign exp_680 = exp_680_reg;
      assign exp_676 = exp_658 ^ exp_661;
  assign exp_658 = exp_657 + exp_656;
  assign exp_657 = 0;
  assign exp_656 = exp_654[31:31];

      reg [31:0] exp_654_reg = 0;
      always@(posedge clk) begin
        if (exp_653) begin
          exp_654_reg <= exp_376;
        end
      end
      assign exp_654 = exp_654_reg;
      assign exp_718 = 0;

      reg [31:0] exp_714_reg = 0;
      always@(posedge clk) begin
        if (exp_647) begin
          exp_714_reg <= exp_684;
        end
      end
      assign exp_714 = exp_714_reg;
    
      reg [31:0] exp_684_reg = 0;
      always@(posedge clk) begin
        if (exp_683) begin
          exp_684_reg <= exp_711;
        end
      end
      assign exp_684 = exp_684_reg;
    
  reg [31:0] exp_711_reg;
  always@(*) begin
    case (exp_645)
      0:exp_711_reg <= exp_703;
      1:exp_711_reg <= exp_709;
      default:exp_711_reg <= exp_710;
    endcase
  end
  assign exp_711 = exp_711_reg;
  assign exp_645 = exp_635 == exp_644;
  assign exp_644 = 2;
  assign exp_710 = 0;

  reg [31:0] exp_703_reg;
  always@(*) begin
    case (exp_693)
      0:exp_703_reg <= exp_697;
      1:exp_703_reg <= exp_701;
      default:exp_703_reg <= exp_702;
    endcase
  end
  assign exp_703 = exp_703_reg;
  assign exp_693 = ~exp_692;
  assign exp_692 = exp_691[32:32];
  assign exp_691 = exp_690 - exp_678;
  assign exp_690 = exp_689;
  assign exp_689 = {exp_687, exp_688};  assign exp_687 = exp_682[31:0];

      reg [31:0] exp_682_reg = 0;
      always@(posedge clk) begin
        if (exp_681) begin
          exp_682_reg <= exp_708;
        end
      end
      assign exp_682 = exp_682_reg;
    
  reg [32:0] exp_708_reg;
  always@(*) begin
    case (exp_645)
      0:exp_708_reg <= exp_695;
      1:exp_708_reg <= exp_706;
      default:exp_708_reg <= exp_707;
    endcase
  end
  assign exp_708 = exp_708_reg;
  assign exp_707 = 0;

  reg [32:0] exp_695_reg;
  always@(*) begin
    case (exp_693)
      0:exp_695_reg <= exp_689;
      1:exp_695_reg <= exp_691;
      default:exp_695_reg <= exp_694;
    endcase
  end
  assign exp_695 = exp_695_reg;
  assign exp_694 = 0;
  assign exp_706 = 0;
  assign exp_681 = 1;
  assign exp_688 = exp_686[31:31];

      reg [31:0] exp_686_reg = 0;
      always@(posedge clk) begin
        if (exp_685) begin
          exp_686_reg <= exp_713;
        end
      end
      assign exp_686 = exp_686_reg;
    
  reg [31:0] exp_713_reg;
  always@(*) begin
    case (exp_645)
      0:exp_713_reg <= exp_705;
      1:exp_713_reg <= exp_677;
      default:exp_713_reg <= exp_712;
    endcase
  end
  assign exp_713 = exp_713_reg;
  assign exp_712 = 0;
  assign exp_705 = exp_686 << exp_704;
  assign exp_704 = 1;

      reg [31:0] exp_677_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_677_reg <= exp_669;
        end
      end
      assign exp_677 = exp_677_reg;
      assign exp_669 = exp_668 + exp_667;
  assign exp_668 = 0;

  reg [31:0] exp_667_reg;
  always@(*) begin
    case (exp_664)
      0:exp_667_reg <= exp_654;
      1:exp_667_reg <= exp_665;
      default:exp_667_reg <= exp_666;
    endcase
  end
  assign exp_667 = exp_667_reg;
  assign exp_664 = exp_658 & exp_632;
  assign exp_666 = 0;
  assign exp_665 = -exp_654;
  assign exp_685 = 1;
  assign exp_702 = 0;
  assign exp_697 = exp_684 << exp_696;
  assign exp_696 = 1;
  assign exp_701 = exp_699 | exp_700;
  assign exp_699 = exp_684 << exp_698;
  assign exp_698 = 1;
  assign exp_700 = 1;
  assign exp_709 = 0;
  assign exp_683 = 1;
  assign exp_647 = exp_635 == exp_646;
  assign exp_646 = 35;
  assign exp_717 = -exp_714;
  assign exp_732 = $signed(exp_731);
  assign exp_731 = -1;
  assign exp_649 = exp_635 == exp_648;
  assign exp_648 = 36;

      reg [31:0] exp_741_reg = 0;
      always@(posedge clk) begin
        if (exp_649) begin
          exp_741_reg <= exp_739;
        end
      end
      assign exp_741 = exp_741_reg;
    
  reg [31:0] exp_739_reg;
  always@(*) begin
    case (exp_737)
      0:exp_739_reg <= exp_727;
      1:exp_739_reg <= exp_654;
      default:exp_739_reg <= exp_738;
    endcase
  end
  assign exp_739 = exp_739_reg;
  assign exp_737 = exp_736 & exp_632;
  assign exp_736 = exp_678 == exp_735;
  assign exp_735 = 0;
  assign exp_738 = 0;
  assign exp_727 = exp_726 + exp_725;
  assign exp_726 = 0;

  reg [31:0] exp_725_reg;
  always@(*) begin
    case (exp_722)
      0:exp_725_reg <= exp_715;
      1:exp_725_reg <= exp_723;
      default:exp_725_reg <= exp_724;
    endcase
  end
  assign exp_725 = exp_725_reg;
  assign exp_722 = exp_679 & exp_632;

      reg [0:0] exp_679_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_679_reg <= exp_658;
        end
      end
      assign exp_679 = exp_679_reg;
      assign exp_724 = 0;

      reg [31:0] exp_715_reg = 0;
      always@(posedge clk) begin
        if (exp_647) begin
          exp_715_reg <= exp_682;
        end
      end
      assign exp_715 = exp_715_reg;
      assign exp_723 = -exp_715;
  assign exp_310 = $signed(exp_309);
  assign exp_309 = 0;
  assign exp_539 = exp_374 != exp_375;
  assign exp_552 = 0;
  assign exp_553 = 0;
  assign exp_540 = $signed(exp_374) < $signed(exp_375);
  assign exp_541 = $signed(exp_374) >= $signed(exp_375);
  assign exp_546 = exp_543 < exp_545;
  assign exp_543 = exp_542 + exp_374;
  assign exp_542 = 0;
  assign exp_545 = exp_544 + exp_375;
  assign exp_544 = 0;
  assign exp_551 = exp_548 >= exp_550;
  assign exp_548 = exp_547 + exp_374;
  assign exp_547 = 0;
  assign exp_550 = exp_549 + exp_375;
  assign exp_549 = 0;
  assign exp_866 = 0;
  assign exp_865 = exp_264 + exp_864;
  assign exp_864 = 4;

  reg [32:0] exp_596_reg;
  always@(*) begin
    case (exp_397)
      0:exp_596_reg <= exp_586;
      1:exp_596_reg <= exp_594;
      default:exp_596_reg <= exp_595;
    endcase
  end
  assign exp_596 = exp_596_reg;
  assign exp_595 = 0;
  assign exp_586 = exp_585 + exp_383;

  reg [31:0] exp_585_reg;
  always@(*) begin
    case (exp_395)
      0:exp_585_reg <= exp_571;
      1:exp_585_reg <= exp_583;
      default:exp_585_reg <= exp_584;
    endcase
  end
  assign exp_585 = exp_585_reg;
  assign exp_584 = 0;
  assign exp_571 = $signed(exp_570);
  assign exp_570 = exp_569 + exp_568;
  assign exp_569 = 0;
  assign exp_568 = {exp_567, exp_564};  assign exp_567 = {exp_566, exp_563};  assign exp_566 = {exp_565, exp_562};  assign exp_565 = {exp_560, exp_561};  assign exp_560 = exp_382[31:31];
  assign exp_561 = exp_382[7:7];
  assign exp_562 = exp_382[30:25];
  assign exp_563 = exp_382[11:8];
  assign exp_564 = 0;
  assign exp_583 = $signed(exp_582);
  assign exp_582 = exp_581 + exp_580;
  assign exp_581 = 0;
  assign exp_580 = {exp_579, exp_576};  assign exp_579 = {exp_578, exp_575};  assign exp_578 = {exp_577, exp_574};  assign exp_577 = {exp_572, exp_573};  assign exp_572 = exp_382[31:31];
  assign exp_573 = exp_382[19:12];
  assign exp_574 = exp_382[20:20];
  assign exp_575 = exp_382[30:21];
  assign exp_576 = 0;

      reg [31:0] exp_383_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_383_reg <= exp_266;
        end
      end
      assign exp_383 = exp_383_reg;
      assign exp_594 = exp_593 & exp_592;
  assign exp_593 = $signed(exp_591);
  assign exp_591 = exp_374 + exp_590;
  assign exp_590 = $signed(exp_589);
  assign exp_589 = exp_588 + exp_587;
  assign exp_588 = 0;
  assign exp_587 = exp_382[31:20];
  assign exp_592 = 4294967294;
  assign exp_263 = exp_256 & exp_254;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_265;
  assign exp_398 = 3;
  assign exp_244 = ~exp_229;
  assign exp_229 = exp_6;
  assign exp_200 = exp_184 & exp_185;
  assign exp_184 = exp_192;
  assign exp_192 = exp_5 & exp_191;
  assign exp_185 = exp_6;
  assign exp_181 = exp_2;

      reg [31:0] exp_221_reg = 0;
      always@(posedge clk) begin
        if (exp_220) begin
          exp_221_reg <= exp_203;
        end
      end
      assign exp_221 = exp_221_reg;
      assign exp_203 = exp_2;
  assign exp_220 = exp_206 & exp_207;
  assign exp_206 = exp_214;
  assign exp_214 = exp_5 & exp_213;
  assign exp_207 = exp_6;
  assign stdin_ready_out = exp_245;
  assign stdout_valid_out = exp_200;
  assign stdout_out = exp_181;
  assign leds_out = exp_221;

endmodule