
module soc(clk, stdin_valid_in, stdin_in, stdout_ready_in, stdin_ready_out, stdout_valid_out, stdout_out, leds_out);
  input [0:0] stdin_valid_in;
  input [31:0] stdin_in;
  input [0:0] stdout_ready_in;
  input [0:0] clk;
  output [0:0] stdin_ready_out;
  output [0:0] stdout_valid_out;
  output [31:0] stdout_out;
  output [31:0] leds_out;
  wire [0:0] exp_245;
  wire [0:0] exp_228;
  wire [0:0] exp_236;
  wire [0:0] exp_5;
  wire [0:0] exp_250;
  wire [0:0] exp_597;
  wire [0:0] exp_534;
  wire [0:0] exp_399;
  wire [6:0] exp_384;
  wire [31:0] exp_382;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [12:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_264;
  wire [32:0] exp_867;
  wire [0:0] exp_863;
  wire [0:0] exp_559;
  wire [0:0] exp_537;
  wire [0:0] exp_395;
  wire [6:0] exp_394;
  wire [0:0] exp_397;
  wire [6:0] exp_396;
  wire [0:0] exp_558;
  wire [0:0] exp_403;
  wire [6:0] exp_402;
  wire [0:0] exp_557;
  wire [0:0] exp_556;
  wire [0:0] exp_555;
  wire [2:0] exp_385;
  wire [0:0] exp_554;
  wire [0:0] exp_538;
  wire [31:0] exp_374;
  wire [31:0] exp_312;
  wire [0:0] exp_308;
  wire [4:0] exp_288;
  wire [0:0] exp_307;
  wire [0:0] exp_311;
  wire [31:0] exp_304;
  wire [0:0] exp_285;
  wire [0:0] exp_858;
  wire [0:0] exp_857;
  wire [0:0] exp_856;
  wire [0:0] exp_855;
  wire [4:0] exp_267;
  wire [4:0] exp_850;
  wire [0:0] exp_849;
  wire [0:0] exp_441;
  wire [0:0] exp_440;
  wire [0:0] exp_439;
  wire [0:0] exp_438;
  wire [0:0] exp_437;
  wire [0:0] exp_436;
  wire [0:0] exp_387;
  wire [4:0] exp_386;
  wire [0:0] exp_389;
  wire [5:0] exp_388;
  wire [0:0] exp_391;
  wire [5:0] exp_390;
  wire [0:0] exp_393;
  wire [4:0] exp_392;
  wire [0:0] exp_844;
  wire [0:0] exp_843;
  wire [0:0] exp_629;
  wire [0:0] exp_603;
  wire [0:0] exp_601;
  wire [6:0] exp_599;
  wire [5:0] exp_600;
  wire [0:0] exp_602;
  wire [0:0] exp_628;
  wire [2:0] exp_598;
  wire [0:0] exp_842;
  wire [0:0] exp_840;
  wire [0:0] exp_833;
  wire [2:0] exp_748;
  wire [2:0] exp_755;
  wire [0:0] exp_750;
  wire [2:0] exp_749;
  wire [0:0] exp_754;
  wire [2:0] exp_752;
  wire [0:0] exp_751;
  wire [0:0] exp_753;
  wire [0:0] exp_744;
  wire [0:0] exp_743;
  wire [0:0] exp_742;
  wire [2:0] exp_832;
  wire [0:0] exp_841;
  wire [0:0] exp_651;
  wire [5:0] exp_635;
  wire [5:0] exp_642;
  wire [0:0] exp_637;
  wire [5:0] exp_636;
  wire [0:0] exp_641;
  wire [5:0] exp_639;
  wire [0:0] exp_638;
  wire [0:0] exp_640;
  wire [5:0] exp_650;
  wire [0:0] exp_262;
  wire [0:0] exp_261;
  wire [0:0] exp_259;
  wire [0:0] exp_258;
  wire [0:0] exp_256;
  wire [0:0] exp_257;
  wire [0:0] exp_255;
  wire [0:0] exp_868;
  wire [0:0] exp_254;
  wire [0:0] exp_253;
  wire [0:0] exp_872;
  wire [0:0] exp_871;
  wire [0:0] exp_870;
  wire [0:0] exp_869;
  wire [0:0] exp_249;
  wire [0:0] exp_240;
  wire [0:0] exp_235;
  wire [0:0] exp_232;
  wire [31:0] exp_1;
  wire [31:0] exp_246;
  wire [31:0] exp_453;
  wire [31:0] exp_452;
  wire [31:0] exp_451;
  wire [31:0] exp_450;
  wire [11:0] exp_449;
  wire [11:0] exp_448;
  wire [11:0] exp_447;
  wire [0:0] exp_401;
  wire [5:0] exp_400;
  wire [0:0] exp_446;
  wire [11:0] exp_442;
  wire [11:0] exp_445;
  wire [6:0] exp_443;
  wire [4:0] exp_444;
  wire [31:0] exp_231;
  wire [0:0] exp_234;
  wire [31:0] exp_233;
  wire [0:0] exp_239;
  wire [0:0] exp_218;
  wire [0:0] exp_213;
  wire [0:0] exp_210;
  wire [31:0] exp_209;
  wire [0:0] exp_212;
  wire [31:0] exp_211;
  wire [0:0] exp_217;
  wire [0:0] exp_196;
  wire [0:0] exp_191;
  wire [0:0] exp_188;
  wire [31:0] exp_187;
  wire [0:0] exp_190;
  wire [31:0] exp_189;
  wire [0:0] exp_195;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [31:0] exp_146;
  wire [0:0] exp_149;
  wire [31:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [14:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_251;
  wire [0:0] exp_536;
  wire [0:0] exp_535;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_176;
  wire [0:0] exp_183;
  wire [0:0] exp_198;
  wire [0:0] exp_205;
  wire [0:0] exp_223;
  wire [0:0] exp_227;
  wire [0:0] exp_243;
  wire [0:0] exp_846;
  wire [0:0] exp_845;
  wire [0:0] exp_260;
  wire [0:0] exp_303;
  wire [31:0] exp_275;
  wire [0:0] exp_274;
  wire [1:0] exp_283;
  wire [4:0] exp_270;
  wire [0:0] exp_273;
  wire [0:0] exp_852;
  wire [0:0] exp_851;
  wire [4:0] exp_269;
  wire [31:0] exp_271;
  wire [31:0] exp_848;
  wire [0:0] exp_847;
  wire [31:0] exp_484;
  wire [0:0] exp_483;
  wire [31:0] exp_435;
  wire [2:0] exp_378;
  wire [2:0] exp_369;
  wire [0:0] exp_366;
  wire [0:0] exp_300;
  wire [6:0] exp_290;
  wire [6:0] exp_299;
  wire [0:0] exp_302;
  wire [6:0] exp_301;
  wire [0:0] exp_368;
  wire [2:0] exp_356;
  wire [0:0] exp_298;
  wire [4:0] exp_297;
  wire [0:0] exp_355;
  wire [2:0] exp_343;
  wire [0:0] exp_296;
  wire [5:0] exp_295;
  wire [0:0] exp_342;
  wire [2:0] exp_292;
  wire [0:0] exp_341;
  wire [0:0] exp_354;
  wire [0:0] exp_367;
  wire [0:0] exp_373;
  wire [0:0] exp_434;
  wire [31:0] exp_414;
  wire [0:0] exp_380;
  wire [0:0] exp_372;
  wire [0:0] exp_358;
  wire [0:0] exp_345;
  wire [0:0] exp_331;
  wire [0:0] exp_329;
  wire [0:0] exp_330;
  wire [0:0] exp_294;
  wire [4:0] exp_293;
  wire [0:0] exp_344;
  wire [0:0] exp_357;
  wire [0:0] exp_371;
  wire [0:0] exp_370;
  wire [0:0] exp_413;
  wire [31:0] exp_411;
  wire [31:0] exp_376;
  wire [31:0] exp_362;
  wire [0:0] exp_359;
  wire [0:0] exp_361;
  wire [31:0] exp_351;
  wire [0:0] exp_350;
  wire [31:0] exp_337;
  wire [0:0] exp_336;
  wire [31:0] exp_335;
  wire [31:0] exp_333;
  wire [19:0] exp_332;
  wire [3:0] exp_334;
  wire [31:0] exp_349;
  wire [31:0] exp_347;
  wire [19:0] exp_346;
  wire [3:0] exp_348;
  wire [31:0] exp_360;
  wire [31:0] exp_377;
  wire [31:0] exp_365;
  wire [0:0] exp_363;
  wire [0:0] exp_364;
  wire [31:0] exp_353;
  wire [0:0] exp_352;
  wire [31:0] exp_340;
  wire [0:0] exp_339;
  wire [31:0] exp_324;
  wire [0:0] exp_323;
  wire [31:0] exp_318;
  wire [0:0] exp_314;
  wire [4:0] exp_289;
  wire [0:0] exp_313;
  wire [0:0] exp_317;
  wire [31:0] exp_306;
  wire [0:0] exp_286;
  wire [0:0] exp_862;
  wire [0:0] exp_861;
  wire [0:0] exp_860;
  wire [0:0] exp_859;
  wire [4:0] exp_268;
  wire [0:0] exp_305;
  wire [31:0] exp_282;
  wire [0:0] exp_281;
  wire [1:0] exp_284;
  wire [4:0] exp_277;
  wire [0:0] exp_280;
  wire [0:0] exp_854;
  wire [0:0] exp_853;
  wire [4:0] exp_276;
  wire [31:0] exp_278;
  wire [31:0] exp_287;
  wire [31:0] exp_316;
  wire [0:0] exp_315;
  wire [31:0] exp_322;
  wire [31:0] exp_319;
  wire [31:0] exp_321;
  wire [11:0] exp_320;
  wire [31:0] exp_338;
  wire [31:0] exp_266;
  wire [0:0] exp_265;
  wire [31:0] exp_412;
  wire [31:0] exp_416;
  wire [31:0] exp_415;
  wire [5:0] exp_410;
  wire [5:0] exp_409;
  wire [5:0] exp_408;
  wire [4:0] exp_379;
  wire [4:0] exp_328;
  wire [0:0] exp_327;
  wire [4:0] exp_326;
  wire [4:0] exp_291;
  wire [31:0] exp_432;
  wire [1:0] exp_418;
  wire [0:0] exp_417;
  wire [31:0] exp_433;
  wire [1:0] exp_424;
  wire [0:0] exp_423;
  wire [31:0] exp_420;
  wire [31:0] exp_419;
  wire [31:0] exp_422;
  wire [31:0] exp_421;
  wire [31:0] exp_425;
  wire [31:0] exp_429;
  wire [32:0] exp_428;
  wire [32:0] exp_426;
  wire [0:0] exp_407;
  wire [0:0] exp_381;
  wire [0:0] exp_325;
  wire [0:0] exp_406;
  wire [0:0] exp_405;
  wire [0:0] exp_404;
  wire [32:0] exp_427;
  wire [31:0] exp_430;
  wire [31:0] exp_431;
  wire [31:0] exp_482;
  wire [0:0] exp_481;
  wire [31:0] exp_472;
  wire [7:0] exp_471;
  wire [7:0] exp_470;
  wire [7:0] exp_465;
  wire [1:0] exp_456;
  wire [1:0] exp_455;
  wire [1:0] exp_454;
  wire [0:0] exp_464;
  wire [7:0] exp_460;
  wire [31:0] exp_248;
  wire [31:0] exp_238;
  wire [0:0] exp_237;
  wire [31:0] exp_216;
  wire [0:0] exp_215;
  wire [31:0] exp_194;
  wire [0:0] exp_193;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [12:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_252;
  wire [3:0] exp_533;
  wire [0:0] exp_532;
  wire [3:0] exp_520;
  wire [3:0] exp_516;
  wire [1:0] exp_519;
  wire [1:0] exp_518;
  wire [1:0] exp_517;
  wire [3:0] exp_525;
  wire [3:0] exp_521;
  wire [0:0] exp_524;
  wire [0:0] exp_523;
  wire [0:0] exp_522;
  wire [3:0] exp_526;
  wire [3:0] exp_527;
  wire [3:0] exp_528;
  wire [3:0] exp_529;
  wire [3:0] exp_530;
  wire [3:0] exp_531;
  wire [12:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_247;
  wire [31:0] exp_515;
  wire [0:0] exp_514;
  wire [31:0] exp_502;
  wire [0:0] exp_501;
  wire [31:0] exp_488;
  wire [7:0] exp_487;
  wire [7:0] exp_486;
  wire [7:0] exp_485;
  wire [31:0] exp_375;
  wire [31:0] exp_496;
  wire [3:0] exp_495;
  wire [31:0] exp_498;
  wire [4:0] exp_497;
  wire [31:0] exp_500;
  wire [4:0] exp_499;
  wire [31:0] exp_506;
  wire [0:0] exp_459;
  wire [0:0] exp_458;
  wire [0:0] exp_457;
  wire [0:0] exp_505;
  wire [31:0] exp_492;
  wire [15:0] exp_491;
  wire [15:0] exp_490;
  wire [15:0] exp_489;
  wire [31:0] exp_504;
  wire [4:0] exp_503;
  wire [31:0] exp_508;
  wire [31:0] exp_507;
  wire [31:0] exp_494;
  wire [31:0] exp_493;
  wire [31:0] exp_509;
  wire [31:0] exp_510;
  wire [31:0] exp_511;
  wire [31:0] exp_512;
  wire [31:0] exp_513;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [12:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [12:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [12:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [12:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [12:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [12:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [12:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [12:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [12:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [12:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [12:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [12:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_179;
  wire [0:0] exp_177;
  wire [31:0] exp_139;
  wire [0:0] exp_178;
  wire [31:0] exp_157;
  wire [31:0] exp_164;
  wire [0:0] exp_159;
  wire [31:0] exp_158;
  wire [0:0] exp_163;
  wire [31:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [31:0] exp_167;
  wire [31:0] exp_174;
  wire [0:0] exp_169;
  wire [31:0] exp_168;
  wire [0:0] exp_173;
  wire [31:0] exp_171;
  wire [0:0] exp_170;
  wire [0:0] exp_172;
  wire [0:0] exp_166;
  wire [0:0] exp_165;
  wire [31:0] exp_182;
  wire [31:0] exp_201;
  wire [31:0] exp_204;
  wire [31:0] exp_222;
  wire [31:0] exp_226;
  wire [31:0] exp_241;
  wire [7:0] exp_461;
  wire [7:0] exp_462;
  wire [7:0] exp_463;
  wire [31:0] exp_475;
  wire [15:0] exp_474;
  wire [15:0] exp_473;
  wire [15:0] exp_469;
  wire [0:0] exp_468;
  wire [15:0] exp_466;
  wire [15:0] exp_467;
  wire [31:0] exp_476;
  wire [31:0] exp_477;
  wire [31:0] exp_478;
  wire [31:0] exp_479;
  wire [31:0] exp_480;
  wire [31:0] exp_839;
  wire [0:0] exp_838;
  wire [31:0] exp_835;
  wire [0:0] exp_606;
  wire [0:0] exp_605;
  wire [0:0] exp_604;
  wire [0:0] exp_834;
  wire [31:0] exp_830;
  wire [63:0] exp_829;
  wire [0:0] exp_826;
  wire [0:0] exp_809;
  wire [0:0] exp_786;
  wire [0:0] exp_783;
  wire [0:0] exp_781;
  wire [0:0] exp_763;
  wire [0:0] exp_762;
  wire [0:0] exp_761;
  wire [31:0] exp_759;
  wire [0:0] exp_758;
  wire [0:0] exp_757;
  wire [0:0] exp_746;
  wire [0:0] exp_745;
  wire [0:0] exp_609;
  wire [0:0] exp_608;
  wire [0:0] exp_607;
  wire [0:0] exp_612;
  wire [0:0] exp_611;
  wire [1:0] exp_610;
  wire [0:0] exp_782;
  wire [0:0] exp_766;
  wire [0:0] exp_765;
  wire [0:0] exp_764;
  wire [31:0] exp_760;
  wire [0:0] exp_747;
  wire [0:0] exp_768;
  wire [0:0] exp_767;
  wire [0:0] exp_788;
  wire [1:0] exp_787;
  wire [0:0] exp_811;
  wire [1:0] exp_810;
  wire [0:0] exp_828;
  wire [63:0] exp_825;
  wire [63:0] exp_824;
  wire [63:0] exp_820;
  wire [63:0] exp_816;
  wire [63:0] exp_812;
  wire [31:0] exp_805;
  wire [31:0] exp_792;
  wire [31:0] exp_790;
  wire [15:0] exp_789;
  wire [31:0] exp_784;
  wire [31:0] exp_774;
  wire [31:0] exp_773;
  wire [31:0] exp_772;
  wire [0:0] exp_769;
  wire [0:0] exp_771;
  wire [31:0] exp_770;
  wire [15:0] exp_791;
  wire [31:0] exp_785;
  wire [31:0] exp_780;
  wire [31:0] exp_779;
  wire [31:0] exp_778;
  wire [0:0] exp_775;
  wire [0:0] exp_777;
  wire [31:0] exp_776;
  wire [63:0] exp_815;
  wire [63:0] exp_813;
  wire [31:0] exp_806;
  wire [31:0] exp_796;
  wire [31:0] exp_794;
  wire [15:0] exp_793;
  wire [15:0] exp_795;
  wire [4:0] exp_814;
  wire [63:0] exp_819;
  wire [63:0] exp_817;
  wire [31:0] exp_807;
  wire [31:0] exp_800;
  wire [31:0] exp_798;
  wire [15:0] exp_797;
  wire [15:0] exp_799;
  wire [4:0] exp_818;
  wire [63:0] exp_823;
  wire [63:0] exp_821;
  wire [31:0] exp_808;
  wire [31:0] exp_804;
  wire [31:0] exp_802;
  wire [15:0] exp_801;
  wire [15:0] exp_803;
  wire [5:0] exp_822;
  wire [63:0] exp_827;
  wire [31:0] exp_831;
  wire [31:0] exp_837;
  wire [0:0] exp_630;
  wire [0:0] exp_836;
  wire [31:0] exp_740;
  wire [31:0] exp_734;
  wire [0:0] exp_730;
  wire [0:0] exp_729;
  wire [31:0] exp_678;
  wire [31:0] exp_675;
  wire [31:0] exp_674;
  wire [31:0] exp_673;
  wire [0:0] exp_670;
  wire [0:0] exp_661;
  wire [0:0] exp_660;
  wire [0:0] exp_659;
  wire [31:0] exp_655;
  wire [0:0] exp_653;
  wire [0:0] exp_652;
  wire [0:0] exp_632;
  wire [0:0] exp_631;
  wire [0:0] exp_672;
  wire [31:0] exp_671;
  wire [0:0] exp_663;
  wire [0:0] exp_662;
  wire [0:0] exp_728;
  wire [0:0] exp_733;
  wire [31:0] exp_721;
  wire [31:0] exp_720;
  wire [31:0] exp_719;
  wire [0:0] exp_716;
  wire [0:0] exp_680;
  wire [0:0] exp_676;
  wire [0:0] exp_658;
  wire [0:0] exp_657;
  wire [0:0] exp_656;
  wire [31:0] exp_654;
  wire [0:0] exp_718;
  wire [31:0] exp_714;
  wire [31:0] exp_684;
  wire [31:0] exp_711;
  wire [0:0] exp_645;
  wire [1:0] exp_644;
  wire [0:0] exp_710;
  wire [31:0] exp_703;
  wire [0:0] exp_693;
  wire [0:0] exp_692;
  wire [32:0] exp_691;
  wire [32:0] exp_690;
  wire [32:0] exp_689;
  wire [31:0] exp_687;
  wire [31:0] exp_682;
  wire [32:0] exp_708;
  wire [0:0] exp_707;
  wire [32:0] exp_695;
  wire [0:0] exp_694;
  wire [0:0] exp_706;
  wire [0:0] exp_681;
  wire [0:0] exp_688;
  wire [31:0] exp_686;
  wire [31:0] exp_713;
  wire [0:0] exp_712;
  wire [31:0] exp_705;
  wire [0:0] exp_704;
  wire [31:0] exp_677;
  wire [31:0] exp_669;
  wire [31:0] exp_668;
  wire [31:0] exp_667;
  wire [0:0] exp_664;
  wire [0:0] exp_666;
  wire [31:0] exp_665;
  wire [0:0] exp_685;
  wire [0:0] exp_702;
  wire [31:0] exp_697;
  wire [0:0] exp_696;
  wire [31:0] exp_701;
  wire [31:0] exp_699;
  wire [0:0] exp_698;
  wire [0:0] exp_700;
  wire [0:0] exp_709;
  wire [0:0] exp_683;
  wire [0:0] exp_647;
  wire [5:0] exp_646;
  wire [31:0] exp_717;
  wire [31:0] exp_732;
  wire [0:0] exp_731;
  wire [0:0] exp_649;
  wire [5:0] exp_648;
  wire [31:0] exp_741;
  wire [31:0] exp_739;
  wire [0:0] exp_737;
  wire [0:0] exp_736;
  wire [0:0] exp_735;
  wire [0:0] exp_738;
  wire [31:0] exp_727;
  wire [31:0] exp_726;
  wire [31:0] exp_725;
  wire [0:0] exp_722;
  wire [0:0] exp_679;
  wire [0:0] exp_724;
  wire [31:0] exp_715;
  wire [31:0] exp_723;
  wire [31:0] exp_310;
  wire [0:0] exp_309;
  wire [0:0] exp_539;
  wire [0:0] exp_552;
  wire [0:0] exp_553;
  wire [0:0] exp_540;
  wire [0:0] exp_541;
  wire [0:0] exp_546;
  wire [31:0] exp_543;
  wire [31:0] exp_542;
  wire [31:0] exp_545;
  wire [31:0] exp_544;
  wire [0:0] exp_551;
  wire [31:0] exp_548;
  wire [31:0] exp_547;
  wire [31:0] exp_550;
  wire [31:0] exp_549;
  wire [0:0] exp_866;
  wire [31:0] exp_865;
  wire [2:0] exp_864;
  wire [32:0] exp_596;
  wire [0:0] exp_595;
  wire [31:0] exp_586;
  wire [31:0] exp_585;
  wire [0:0] exp_584;
  wire [31:0] exp_571;
  wire [12:0] exp_570;
  wire [12:0] exp_569;
  wire [12:0] exp_568;
  wire [11:0] exp_567;
  wire [7:0] exp_566;
  wire [1:0] exp_565;
  wire [0:0] exp_560;
  wire [0:0] exp_561;
  wire [5:0] exp_562;
  wire [3:0] exp_563;
  wire [0:0] exp_564;
  wire [31:0] exp_583;
  wire [20:0] exp_582;
  wire [20:0] exp_581;
  wire [20:0] exp_580;
  wire [19:0] exp_579;
  wire [9:0] exp_578;
  wire [8:0] exp_577;
  wire [0:0] exp_572;
  wire [7:0] exp_573;
  wire [0:0] exp_574;
  wire [9:0] exp_575;
  wire [0:0] exp_576;
  wire [31:0] exp_383;
  wire [32:0] exp_594;
  wire [32:0] exp_593;
  wire [31:0] exp_591;
  wire [31:0] exp_590;
  wire [11:0] exp_589;
  wire [11:0] exp_588;
  wire [11:0] exp_587;
  wire [32:0] exp_592;
  wire [0:0] exp_263;
  wire [0:0] exp_80;
  wire [12:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_398;
  wire [0:0] exp_244;
  wire [0:0] exp_229;
  wire [0:0] exp_200;
  wire [0:0] exp_184;
  wire [0:0] exp_192;
  wire [0:0] exp_185;
  wire [31:0] exp_181;
  wire [31:0] exp_221;
  wire [31:0] exp_203;
  wire [0:0] exp_220;
  wire [0:0] exp_206;
  wire [0:0] exp_214;
  wire [0:0] exp_207;

  assign exp_245 = exp_228 & exp_244;
  assign exp_228 = exp_236;
  assign exp_236 = exp_5 & exp_235;
  assign exp_5 = exp_250;
  assign exp_250 = exp_597;
  assign exp_597 = exp_534 & exp_262;
  assign exp_534 = exp_399 | exp_401;
  assign exp_399 = exp_384 == exp_398;
  assign exp_384 = exp_382[6:0];

      reg [31:0] exp_382_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_382_reg <= exp_96;
        end
      end
      assign exp_382 = exp_382_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_264;

      reg [31:0] exp_264_reg = 0;
      always@(posedge clk) begin
        if (exp_263) begin
          exp_264_reg <= exp_867;
        end
      end
      assign exp_264 = exp_264_reg;
    
  reg [32:0] exp_867_reg;
  always@(*) begin
    case (exp_863)
      0:exp_867_reg <= exp_865;
      1:exp_867_reg <= exp_596;
      default:exp_867_reg <= exp_866;
    endcase
  end
  assign exp_867 = exp_867_reg;
  assign exp_863 = exp_559 & exp_262;
  assign exp_559 = exp_537 | exp_558;
  assign exp_537 = exp_395 | exp_397;
  assign exp_395 = exp_384 == exp_394;
  assign exp_394 = 111;
  assign exp_397 = exp_384 == exp_396;
  assign exp_396 = 103;

  reg [0:0] exp_558_reg;
  always@(*) begin
    case (exp_403)
      0:exp_558_reg <= exp_556;
      1:exp_558_reg <= exp_555;
      default:exp_558_reg <= exp_557;
    endcase
  end
  assign exp_558 = exp_558_reg;
  assign exp_403 = exp_384 == exp_402;
  assign exp_402 = 99;
  assign exp_557 = 0;
  assign exp_556 = 0;

  reg [0:0] exp_555_reg;
  always@(*) begin
    case (exp_385)
      0:exp_555_reg <= exp_538;
      1:exp_555_reg <= exp_539;
      2:exp_555_reg <= exp_552;
      3:exp_555_reg <= exp_553;
      4:exp_555_reg <= exp_540;
      5:exp_555_reg <= exp_541;
      6:exp_555_reg <= exp_546;
      7:exp_555_reg <= exp_551;
      default:exp_555_reg <= exp_554;
    endcase
  end
  assign exp_555 = exp_555_reg;
  assign exp_385 = exp_382[14:12];
  assign exp_554 = 0;
  assign exp_538 = exp_374 == exp_375;

      reg [31:0] exp_374_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_374_reg <= exp_312;
        end
      end
      assign exp_374 = exp_374_reg;
    
  reg [31:0] exp_312_reg;
  always@(*) begin
    case (exp_308)
      0:exp_312_reg <= exp_304;
      1:exp_312_reg <= exp_310;
      default:exp_312_reg <= exp_311;
    endcase
  end
  assign exp_312 = exp_312_reg;
  assign exp_308 = exp_288 == exp_307;
  assign exp_288 = exp_96[19:15];
  assign exp_307 = 0;
  assign exp_311 = 0;

  reg [31:0] exp_304_reg;
  always@(*) begin
    case (exp_285)
      0:exp_304_reg <= exp_275;
      1:exp_304_reg <= exp_287;
      default:exp_304_reg <= exp_303;
    endcase
  end
  assign exp_304 = exp_304_reg;
  assign exp_285 = exp_858;
  assign exp_858 = exp_857 & exp_254;
  assign exp_857 = exp_856 & exp_262;
  assign exp_856 = exp_855 & exp_849;
  assign exp_855 = exp_267 == exp_850;
  assign exp_267 = exp_96[19:15];
  assign exp_850 = exp_382[11:7];
  assign exp_849 = exp_441 | exp_844;
  assign exp_441 = exp_440 | exp_399;
  assign exp_440 = exp_439 | exp_393;
  assign exp_439 = exp_438 | exp_391;
  assign exp_438 = exp_437 | exp_397;
  assign exp_437 = exp_436 | exp_395;
  assign exp_436 = exp_387 | exp_389;
  assign exp_387 = exp_384 == exp_386;
  assign exp_386 = 19;
  assign exp_389 = exp_384 == exp_388;
  assign exp_388 = 51;
  assign exp_391 = exp_384 == exp_390;
  assign exp_390 = 55;
  assign exp_393 = exp_384 == exp_392;
  assign exp_392 = 23;
  assign exp_844 = exp_843 & exp_603;

  reg [0:0] exp_843_reg;
  always@(*) begin
    case (exp_629)
      0:exp_843_reg <= exp_840;
      1:exp_843_reg <= exp_841;
      default:exp_843_reg <= exp_842;
    endcase
  end
  assign exp_843 = exp_843_reg;
  assign exp_629 = exp_603 & exp_628;
  assign exp_603 = exp_601 & exp_602;
  assign exp_601 = exp_599 == exp_600;
  assign exp_599 = exp_382[6:0];
  assign exp_600 = 51;
  assign exp_602 = exp_382[25:25];
  assign exp_628 = exp_598[2:2];
  assign exp_598 = exp_382[14:12];
  assign exp_842 = 0;
  assign exp_840 = exp_833 & exp_603;
  assign exp_833 = exp_748 == exp_832;

      reg [2:0] exp_748_reg = 0;
      always@(posedge clk) begin
        if (exp_744) begin
          exp_748_reg <= exp_755;
        end
      end
      assign exp_748 = exp_748_reg;
    
  reg [2:0] exp_755_reg;
  always@(*) begin
    case (exp_750)
      0:exp_755_reg <= exp_752;
      1:exp_755_reg <= exp_753;
      default:exp_755_reg <= exp_754;
    endcase
  end
  assign exp_755 = exp_755_reg;
  assign exp_750 = exp_748 == exp_749;
  assign exp_749 = 4;
  assign exp_754 = 0;
  assign exp_752 = exp_748 + exp_751;
  assign exp_751 = 1;
  assign exp_753 = 0;
  assign exp_744 = exp_603 & exp_743;
  assign exp_743 = ~exp_742;
  assign exp_742 = exp_598[2:2];
  assign exp_832 = 4;
  assign exp_841 = exp_651 & exp_603;
  assign exp_651 = exp_635 == exp_650;

      reg [5:0] exp_635_reg = 0;
      always@(posedge clk) begin
        if (exp_629) begin
          exp_635_reg <= exp_642;
        end
      end
      assign exp_635 = exp_635_reg;
    
  reg [5:0] exp_642_reg;
  always@(*) begin
    case (exp_637)
      0:exp_642_reg <= exp_639;
      1:exp_642_reg <= exp_640;
      default:exp_642_reg <= exp_641;
    endcase
  end
  assign exp_642 = exp_642_reg;
  assign exp_637 = exp_635 == exp_636;
  assign exp_636 = 37;
  assign exp_641 = 0;
  assign exp_639 = exp_635 + exp_638;
  assign exp_638 = 1;
  assign exp_640 = 0;
  assign exp_650 = 37;

      reg [0:0] exp_262_reg = 0;
      always@(posedge clk) begin
        if (exp_254) begin
          exp_262_reg <= exp_261;
        end
      end
      assign exp_262 = exp_262_reg;
      assign exp_261 = exp_259 & exp_260;

      reg [0:0] exp_259_reg = 0;
      always@(posedge clk) begin
        if (exp_254) begin
          exp_259_reg <= exp_258;
        end
      end
      assign exp_259 = exp_259_reg;
      assign exp_258 = exp_256 & exp_257;
  assign exp_256 = 1;
  assign exp_257 = ~exp_255;
  assign exp_255 = exp_868;
  assign exp_868 = exp_262 & exp_559;
  assign exp_254 = ~exp_253;
  assign exp_253 = exp_872;
  assign exp_872 = exp_262 & exp_871;
  assign exp_871 = exp_870 | exp_846;
  assign exp_870 = exp_250 & exp_869;
  assign exp_869 = ~exp_249;
  assign exp_249 = exp_240;

  reg [0:0] exp_240_reg;
  always@(*) begin
    case (exp_235)
      0:exp_240_reg <= exp_218;
      1:exp_240_reg <= exp_227;
      default:exp_240_reg <= exp_239;
    endcase
  end
  assign exp_240 = exp_240_reg;
  assign exp_235 = exp_232 & exp_234;
  assign exp_232 = exp_1 >= exp_231;
  assign exp_1 = exp_246;
  assign exp_246 = exp_453;
  assign exp_453 = exp_452 + exp_451;
  assign exp_452 = 0;
  assign exp_451 = exp_374 + exp_450;
  assign exp_450 = $signed(exp_449);
  assign exp_449 = exp_448 + exp_447;
  assign exp_448 = 0;

  reg [11:0] exp_447_reg;
  always@(*) begin
    case (exp_401)
      0:exp_447_reg <= exp_442;
      1:exp_447_reg <= exp_445;
      default:exp_447_reg <= exp_446;
    endcase
  end
  assign exp_447 = exp_447_reg;
  assign exp_401 = exp_384 == exp_400;
  assign exp_400 = 35;
  assign exp_446 = 0;
  assign exp_442 = exp_382[31:20];
  assign exp_445 = {exp_443, exp_444};  assign exp_443 = exp_382[31:25];
  assign exp_444 = exp_382[11:7];
  assign exp_231 = 2147483664;
  assign exp_234 = exp_1 <= exp_233;
  assign exp_233 = 2147483664;
  assign exp_239 = 0;

  reg [0:0] exp_218_reg;
  always@(*) begin
    case (exp_213)
      0:exp_218_reg <= exp_196;
      1:exp_218_reg <= exp_205;
      default:exp_218_reg <= exp_217;
    endcase
  end
  assign exp_218 = exp_218_reg;
  assign exp_213 = exp_210 & exp_212;
  assign exp_210 = exp_1 >= exp_209;
  assign exp_209 = 2147483660;
  assign exp_212 = exp_1 <= exp_211;
  assign exp_211 = 2147483660;
  assign exp_217 = 0;

  reg [0:0] exp_196_reg;
  always@(*) begin
    case (exp_191)
      0:exp_196_reg <= exp_155;
      1:exp_196_reg <= exp_183;
      default:exp_196_reg <= exp_195;
    endcase
  end
  assign exp_196 = exp_196_reg;
  assign exp_191 = exp_188 & exp_190;
  assign exp_188 = exp_1 >= exp_187;
  assign exp_187 = 2147483656;
  assign exp_190 = exp_1 <= exp_189;
  assign exp_189 = 2147483656;
  assign exp_195 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 2147483648;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 2147483652;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 20476;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_251;
  assign exp_251 = exp_536;
  assign exp_536 = exp_535 + exp_401;
  assign exp_535 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_176;
  assign exp_176 = 1;
  assign exp_183 = exp_198;
  assign exp_198 = stdout_ready_in;
  assign exp_205 = exp_223;
  assign exp_223 = 1;
  assign exp_227 = exp_243;
  assign exp_243 = stdin_valid_in;
  assign exp_846 = exp_603 & exp_845;
  assign exp_845 = ~exp_843;
  assign exp_260 = ~exp_255;
  assign exp_303 = 0;

  //Create RAM
  reg [31:0] exp_275_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_273) begin
      exp_275_ram[exp_269] <= exp_271;
    end
  end
  assign exp_275 = exp_275_ram[exp_270];
  assign exp_274 = exp_283;
  assign exp_283 = 1;
  assign exp_270 = exp_267;
  assign exp_273 = exp_852;
  assign exp_852 = exp_851 & exp_254;
  assign exp_851 = exp_849 & exp_262;
  assign exp_269 = exp_850;
  assign exp_271 = exp_848;

  reg [31:0] exp_848_reg;
  always@(*) begin
    case (exp_844)
      0:exp_848_reg <= exp_484;
      1:exp_848_reg <= exp_839;
      default:exp_848_reg <= exp_847;
    endcase
  end
  assign exp_848 = exp_848_reg;
  assign exp_847 = 0;

  reg [31:0] exp_484_reg;
  always@(*) begin
    case (exp_399)
      0:exp_484_reg <= exp_435;
      1:exp_484_reg <= exp_482;
      default:exp_484_reg <= exp_483;
    endcase
  end
  assign exp_484 = exp_484_reg;
  assign exp_483 = 0;

  reg [31:0] exp_435_reg;
  always@(*) begin
    case (exp_378)
      0:exp_435_reg <= exp_414;
      1:exp_435_reg <= exp_416;
      2:exp_435_reg <= exp_432;
      3:exp_435_reg <= exp_433;
      4:exp_435_reg <= exp_425;
      5:exp_435_reg <= exp_429;
      6:exp_435_reg <= exp_430;
      7:exp_435_reg <= exp_431;
      default:exp_435_reg <= exp_434;
    endcase
  end
  assign exp_435 = exp_435_reg;

      reg [2:0] exp_378_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_378_reg <= exp_369;
        end
      end
      assign exp_378 = exp_378_reg;
    
  reg [2:0] exp_369_reg;
  always@(*) begin
    case (exp_366)
      0:exp_369_reg <= exp_356;
      1:exp_369_reg <= exp_367;
      default:exp_369_reg <= exp_368;
    endcase
  end
  assign exp_369 = exp_369_reg;
  assign exp_366 = exp_300 | exp_302;
  assign exp_300 = exp_290 == exp_299;
  assign exp_290 = exp_96[6:0];
  assign exp_299 = 111;
  assign exp_302 = exp_290 == exp_301;
  assign exp_301 = 103;
  assign exp_368 = 0;

  reg [2:0] exp_356_reg;
  always@(*) begin
    case (exp_298)
      0:exp_356_reg <= exp_343;
      1:exp_356_reg <= exp_354;
      default:exp_356_reg <= exp_355;
    endcase
  end
  assign exp_356 = exp_356_reg;
  assign exp_298 = exp_290 == exp_297;
  assign exp_297 = 23;
  assign exp_355 = 0;

  reg [2:0] exp_343_reg;
  always@(*) begin
    case (exp_296)
      0:exp_343_reg <= exp_292;
      1:exp_343_reg <= exp_341;
      default:exp_343_reg <= exp_342;
    endcase
  end
  assign exp_343 = exp_343_reg;
  assign exp_296 = exp_290 == exp_295;
  assign exp_295 = 55;
  assign exp_342 = 0;
  assign exp_292 = exp_96[14:12];
  assign exp_341 = 0;
  assign exp_354 = 0;
  assign exp_367 = 0;
  assign exp_373 = exp_254 & exp_259;
  assign exp_434 = 0;

  reg [31:0] exp_414_reg;
  always@(*) begin
    case (exp_380)
      0:exp_414_reg <= exp_411;
      1:exp_414_reg <= exp_412;
      default:exp_414_reg <= exp_413;
    endcase
  end
  assign exp_414 = exp_414_reg;

      reg [0:0] exp_380_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_380_reg <= exp_372;
        end
      end
      assign exp_380 = exp_380_reg;
      assign exp_372 = exp_358 & exp_371;
  assign exp_358 = exp_345 & exp_357;
  assign exp_345 = exp_331 & exp_344;
  assign exp_331 = exp_329 & exp_330;
  assign exp_329 = exp_96[30:30];
  assign exp_330 = ~exp_294;
  assign exp_294 = exp_290 == exp_293;
  assign exp_293 = 19;
  assign exp_344 = ~exp_296;
  assign exp_357 = ~exp_298;
  assign exp_371 = ~exp_370;
  assign exp_370 = exp_300 | exp_302;
  assign exp_413 = 0;
  assign exp_411 = exp_376 + exp_377;

      reg [31:0] exp_376_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_376_reg <= exp_362;
        end
      end
      assign exp_376 = exp_376_reg;
    
  reg [31:0] exp_362_reg;
  always@(*) begin
    case (exp_359)
      0:exp_362_reg <= exp_351;
      1:exp_362_reg <= exp_360;
      default:exp_362_reg <= exp_361;
    endcase
  end
  assign exp_362 = exp_362_reg;
  assign exp_359 = exp_300 | exp_302;
  assign exp_361 = 0;

  reg [31:0] exp_351_reg;
  always@(*) begin
    case (exp_298)
      0:exp_351_reg <= exp_337;
      1:exp_351_reg <= exp_349;
      default:exp_351_reg <= exp_350;
    endcase
  end
  assign exp_351 = exp_351_reg;
  assign exp_350 = 0;

  reg [31:0] exp_337_reg;
  always@(*) begin
    case (exp_296)
      0:exp_337_reg <= exp_312;
      1:exp_337_reg <= exp_335;
      default:exp_337_reg <= exp_336;
    endcase
  end
  assign exp_337 = exp_337_reg;
  assign exp_336 = 0;
  assign exp_335 = exp_333 << exp_334;
  assign exp_333 = exp_332;
  assign exp_332 = exp_96[31:12];
  assign exp_334 = 12;
  assign exp_349 = exp_347 << exp_348;
  assign exp_347 = exp_346;
  assign exp_346 = exp_96[31:12];
  assign exp_348 = 12;
  assign exp_360 = 4;

      reg [31:0] exp_377_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_377_reg <= exp_365;
        end
      end
      assign exp_377 = exp_377_reg;
    
  reg [31:0] exp_365_reg;
  always@(*) begin
    case (exp_363)
      0:exp_365_reg <= exp_353;
      1:exp_365_reg <= exp_266;
      default:exp_365_reg <= exp_364;
    endcase
  end
  assign exp_365 = exp_365_reg;
  assign exp_363 = exp_300 | exp_302;
  assign exp_364 = 0;

  reg [31:0] exp_353_reg;
  always@(*) begin
    case (exp_298)
      0:exp_353_reg <= exp_340;
      1:exp_353_reg <= exp_266;
      default:exp_353_reg <= exp_352;
    endcase
  end
  assign exp_353 = exp_353_reg;
  assign exp_352 = 0;

  reg [31:0] exp_340_reg;
  always@(*) begin
    case (exp_296)
      0:exp_340_reg <= exp_324;
      1:exp_340_reg <= exp_338;
      default:exp_340_reg <= exp_339;
    endcase
  end
  assign exp_340 = exp_340_reg;
  assign exp_339 = 0;

  reg [31:0] exp_324_reg;
  always@(*) begin
    case (exp_294)
      0:exp_324_reg <= exp_318;
      1:exp_324_reg <= exp_322;
      default:exp_324_reg <= exp_323;
    endcase
  end
  assign exp_324 = exp_324_reg;
  assign exp_323 = 0;

  reg [31:0] exp_318_reg;
  always@(*) begin
    case (exp_314)
      0:exp_318_reg <= exp_306;
      1:exp_318_reg <= exp_316;
      default:exp_318_reg <= exp_317;
    endcase
  end
  assign exp_318 = exp_318_reg;
  assign exp_314 = exp_289 == exp_313;
  assign exp_289 = exp_96[24:20];
  assign exp_313 = 0;
  assign exp_317 = 0;

  reg [31:0] exp_306_reg;
  always@(*) begin
    case (exp_286)
      0:exp_306_reg <= exp_282;
      1:exp_306_reg <= exp_287;
      default:exp_306_reg <= exp_305;
    endcase
  end
  assign exp_306 = exp_306_reg;
  assign exp_286 = exp_862;
  assign exp_862 = exp_861 & exp_254;
  assign exp_861 = exp_860 & exp_262;
  assign exp_860 = exp_859 & exp_849;
  assign exp_859 = exp_268 == exp_850;
  assign exp_268 = exp_96[24:20];
  assign exp_305 = 0;

  //Create RAM
  reg [31:0] exp_282_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_280) begin
      exp_282_ram[exp_276] <= exp_278;
    end
  end
  assign exp_282 = exp_282_ram[exp_277];
  assign exp_281 = exp_284;
  assign exp_284 = 1;
  assign exp_277 = exp_268;
  assign exp_280 = exp_854;
  assign exp_854 = exp_853 & exp_254;
  assign exp_853 = exp_849 & exp_262;
  assign exp_276 = exp_850;
  assign exp_278 = exp_848;
  assign exp_287 = exp_848;
  assign exp_316 = $signed(exp_315);
  assign exp_315 = 0;
  assign exp_322 = exp_319 + exp_321;
  assign exp_319 = 0;
  assign exp_321 = $signed(exp_320);
  assign exp_320 = exp_96[31:20];
  assign exp_338 = 0;

      reg [31:0] exp_266_reg = 0;
      always@(posedge clk) begin
        if (exp_265) begin
          exp_266_reg <= exp_264;
        end
      end
      assign exp_266 = exp_266_reg;
      assign exp_265 = exp_256 & exp_254;
  assign exp_412 = exp_376 - exp_377;
  assign exp_416 = exp_376 << exp_415;
  assign exp_415 = $signed(exp_410);
  assign exp_410 = exp_409 + exp_408;
  assign exp_409 = 0;
  assign exp_408 = exp_379;

      reg [4:0] exp_379_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_379_reg <= exp_328;
        end
      end
      assign exp_379 = exp_379_reg;
    
  reg [4:0] exp_328_reg;
  always@(*) begin
    case (exp_294)
      0:exp_328_reg <= exp_326;
      1:exp_328_reg <= exp_291;
      default:exp_328_reg <= exp_327;
    endcase
  end
  assign exp_328 = exp_328_reg;
  assign exp_327 = 0;
  assign exp_326 = exp_324[4:0];
  assign exp_291 = exp_96[24:20];
  assign exp_432 = $signed(exp_418);
  assign exp_418 = exp_417;
  assign exp_417 = $signed(exp_376) < $signed(exp_377);
  assign exp_433 = $signed(exp_424);
  assign exp_424 = exp_423;
  assign exp_423 = exp_420 < exp_422;
  assign exp_420 = exp_419 + exp_376;
  assign exp_419 = 0;
  assign exp_422 = exp_421 + exp_377;
  assign exp_421 = 0;
  assign exp_425 = exp_376 ^ exp_377;
  assign exp_429 = exp_428[31:0];
  assign exp_428 = $signed(exp_426) >>> $signed(exp_427);
  assign exp_426 = {exp_407, exp_376};
  reg [0:0] exp_407_reg;
  always@(*) begin
    case (exp_381)
      0:exp_407_reg <= exp_405;
      1:exp_407_reg <= exp_404;
      default:exp_407_reg <= exp_406;
    endcase
  end
  assign exp_407 = exp_407_reg;

      reg [0:0] exp_381_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_381_reg <= exp_325;
        end
      end
      assign exp_381 = exp_381_reg;
      assign exp_325 = exp_96[30:30];
  assign exp_406 = 0;
  assign exp_405 = 0;
  assign exp_404 = exp_376[31:31];
  assign exp_427 = $signed(exp_410);
  assign exp_430 = exp_376 | exp_377;
  assign exp_431 = exp_376 & exp_377;

  reg [31:0] exp_482_reg;
  always@(*) begin
    case (exp_385)
      0:exp_482_reg <= exp_472;
      1:exp_482_reg <= exp_475;
      2:exp_482_reg <= exp_248;
      3:exp_482_reg <= exp_476;
      4:exp_482_reg <= exp_477;
      5:exp_482_reg <= exp_478;
      6:exp_482_reg <= exp_479;
      7:exp_482_reg <= exp_480;
      default:exp_482_reg <= exp_481;
    endcase
  end
  assign exp_482 = exp_482_reg;
  assign exp_481 = 0;
  assign exp_472 = $signed(exp_471);
  assign exp_471 = exp_470 + exp_465;
  assign exp_470 = 0;

  reg [7:0] exp_465_reg;
  always@(*) begin
    case (exp_456)
      0:exp_465_reg <= exp_460;
      1:exp_465_reg <= exp_461;
      2:exp_465_reg <= exp_462;
      3:exp_465_reg <= exp_463;
      default:exp_465_reg <= exp_464;
    endcase
  end
  assign exp_465 = exp_465_reg;
  assign exp_456 = exp_455 + exp_454;
  assign exp_455 = 0;
  assign exp_454 = exp_453[1:0];
  assign exp_464 = 0;
  assign exp_460 = exp_248[7:0];
  assign exp_248 = exp_238;

  reg [31:0] exp_238_reg;
  always@(*) begin
    case (exp_235)
      0:exp_238_reg <= exp_216;
      1:exp_238_reg <= exp_226;
      default:exp_238_reg <= exp_237;
    endcase
  end
  assign exp_238 = exp_238_reg;
  assign exp_237 = 0;

  reg [31:0] exp_216_reg;
  always@(*) begin
    case (exp_213)
      0:exp_216_reg <= exp_194;
      1:exp_216_reg <= exp_204;
      default:exp_216_reg <= exp_215;
    endcase
  end
  assign exp_216 = exp_216_reg;
  assign exp_215 = 0;

  reg [31:0] exp_194_reg;
  always@(*) begin
    case (exp_191)
      0:exp_194_reg <= exp_153;
      1:exp_194_reg <= exp_182;
      default:exp_194_reg <= exp_193;
    endcase
  end
  assign exp_194 = exp_194_reg;
  assign exp_193 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 0;
    exp_54_ram[32] = 252;
    exp_54_ram[33] = 81;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 0;
    exp_54_ram[36] = 99;
    exp_54_ram[37] = 46;
    exp_54_ram[38] = 0;
    exp_54_ram[39] = 0;
    exp_54_ram[40] = 108;
    exp_54_ram[41] = 0;
    exp_54_ram[42] = 97;
    exp_54_ram[43] = 0;
    exp_54_ram[44] = 97;
    exp_54_ram[45] = 0;
    exp_54_ram[46] = 0;
    exp_54_ram[47] = 97;
    exp_54_ram[48] = 0;
    exp_54_ram[49] = 97;
    exp_54_ram[50] = 0;
    exp_54_ram[51] = 115;
    exp_54_ram[52] = 0;
    exp_54_ram[53] = 110;
    exp_54_ram[54] = 46;
    exp_54_ram[55] = 0;
    exp_54_ram[56] = 120;
    exp_54_ram[57] = 0;
    exp_54_ram[58] = 99;
    exp_54_ram[59] = 46;
    exp_54_ram[60] = 0;
    exp_54_ram[61] = 99;
    exp_54_ram[62] = 46;
    exp_54_ram[63] = 0;
    exp_54_ram[64] = 110;
    exp_54_ram[65] = 46;
    exp_54_ram[66] = 0;
    exp_54_ram[67] = 99;
    exp_54_ram[68] = 46;
    exp_54_ram[69] = 0;
    exp_54_ram[70] = 97;
    exp_54_ram[71] = 0;
    exp_54_ram[72] = 99;
    exp_54_ram[73] = 46;
    exp_54_ram[74] = 0;
    exp_54_ram[75] = 97;
    exp_54_ram[76] = 0;
    exp_54_ram[77] = 99;
    exp_54_ram[78] = 46;
    exp_54_ram[79] = 0;
    exp_54_ram[80] = 102;
    exp_54_ram[81] = 0;
    exp_54_ram[82] = 102;
    exp_54_ram[83] = 102;
    exp_54_ram[84] = 0;
    exp_54_ram[85] = 102;
    exp_54_ram[86] = 102;
    exp_54_ram[87] = 0;
    exp_54_ram[88] = 97;
    exp_54_ram[89] = 52;
    exp_54_ram[90] = 0;
    exp_54_ram[91] = 102;
    exp_54_ram[92] = 102;
    exp_54_ram[93] = 0;
    exp_54_ram[94] = 112;
    exp_54_ram[95] = 46;
    exp_54_ram[96] = 0;
    exp_54_ram[97] = 102;
    exp_54_ram[98] = 49;
    exp_54_ram[99] = 0;
    exp_54_ram[100] = 50;
    exp_54_ram[101] = 0;
    exp_54_ram[102] = 51;
    exp_54_ram[103] = 0;
    exp_54_ram[104] = 100;
    exp_54_ram[105] = 0;
    exp_54_ram[106] = 102;
    exp_54_ram[107] = 102;
    exp_54_ram[108] = 0;
    exp_54_ram[109] = 114;
    exp_54_ram[110] = 46;
    exp_54_ram[111] = 0;
    exp_54_ram[112] = 115;
    exp_54_ram[113] = 46;
    exp_54_ram[114] = 0;
    exp_54_ram[115] = 100;
    exp_54_ram[116] = 0;
    exp_54_ram[117] = 100;
    exp_54_ram[118] = 115;
    exp_54_ram[119] = 0;
    exp_54_ram[120] = 102;
    exp_54_ram[121] = 50;
    exp_54_ram[122] = 0;
    exp_54_ram[123] = 100;
    exp_54_ram[124] = 52;
    exp_54_ram[125] = 102;
    exp_54_ram[126] = 0;
    exp_54_ram[127] = 115;
    exp_54_ram[128] = 46;
    exp_54_ram[129] = 0;
    exp_54_ram[130] = 52;
    exp_54_ram[131] = 0;
    exp_54_ram[132] = 0;
    exp_54_ram[133] = 0;
    exp_54_ram[134] = 115;
    exp_54_ram[135] = 46;
    exp_54_ram[136] = 0;
    exp_54_ram[137] = 52;
    exp_54_ram[138] = 0;
    exp_54_ram[139] = 52;
    exp_54_ram[140] = 0;
    exp_54_ram[141] = 52;
    exp_54_ram[142] = 0;
    exp_54_ram[143] = 100;
    exp_54_ram[144] = 0;
    exp_54_ram[145] = 108;
    exp_54_ram[146] = 46;
    exp_54_ram[147] = 0;
    exp_54_ram[148] = 101;
    exp_54_ram[149] = 0;
    exp_54_ram[150] = 32;
    exp_54_ram[151] = 32;
    exp_54_ram[152] = 48;
    exp_54_ram[153] = 49;
    exp_54_ram[154] = 32;
    exp_54_ram[155] = 48;
    exp_54_ram[156] = 0;
    exp_54_ram[157] = 32;
    exp_54_ram[158] = 32;
    exp_54_ram[159] = 48;
    exp_54_ram[160] = 49;
    exp_54_ram[161] = 32;
    exp_54_ram[162] = 48;
    exp_54_ram[163] = 0;
    exp_54_ram[164] = 97;
    exp_54_ram[165] = 0;
    exp_54_ram[166] = 97;
    exp_54_ram[167] = 0;
    exp_54_ram[168] = 97;
    exp_54_ram[169] = 0;
    exp_54_ram[170] = 32;
    exp_54_ram[171] = 32;
    exp_54_ram[172] = 48;
    exp_54_ram[173] = 49;
    exp_54_ram[174] = 32;
    exp_54_ram[175] = 48;
    exp_54_ram[176] = 0;
    exp_54_ram[177] = 102;
    exp_54_ram[178] = 0;
    exp_54_ram[179] = 102;
    exp_54_ram[180] = 0;
    exp_54_ram[181] = 102;
    exp_54_ram[182] = 0;
    exp_54_ram[183] = 116;
    exp_54_ram[184] = 105;
    exp_54_ram[185] = 32;
    exp_54_ram[186] = 0;
    exp_54_ram[187] = 0;
    exp_54_ram[188] = 46;
    exp_54_ram[189] = 10;
    exp_54_ram[190] = 0;
    exp_54_ram[191] = 0;
    exp_54_ram[192] = 116;
    exp_54_ram[193] = 48;
    exp_54_ram[194] = 48;
    exp_54_ram[195] = 10;
    exp_54_ram[196] = 0;
    exp_54_ram[197] = 0;
    exp_54_ram[198] = 0;
    exp_54_ram[199] = 0;
    exp_54_ram[200] = 160;
    exp_54_ram[201] = 62;
    exp_54_ram[202] = 136;
    exp_54_ram[203] = 62;
    exp_54_ram[204] = 235;
    exp_54_ram[205] = 63;
    exp_54_ram[206] = 210;
    exp_54_ram[207] = 63;
    exp_54_ram[208] = 71;
    exp_54_ram[209] = 63;
    exp_54_ram[210] = 153;
    exp_54_ram[211] = 63;
    exp_54_ram[212] = 0;
    exp_54_ram[213] = 63;
    exp_54_ram[214] = 0;
    exp_54_ram[215] = 64;
    exp_54_ram[216] = 0;
    exp_54_ram[217] = 64;
    exp_54_ram[218] = 0;
    exp_54_ram[219] = 64;
    exp_54_ram[220] = 0;
    exp_54_ram[221] = 64;
    exp_54_ram[222] = 0;
    exp_54_ram[223] = 64;
    exp_54_ram[224] = 0;
    exp_54_ram[225] = 65;
    exp_54_ram[226] = 0;
    exp_54_ram[227] = 65;
    exp_54_ram[228] = 0;
    exp_54_ram[229] = 65;
    exp_54_ram[230] = 0;
    exp_54_ram[231] = 65;
    exp_54_ram[232] = 0;
    exp_54_ram[233] = 127;
    exp_54_ram[234] = 0;
    exp_54_ram[235] = 255;
    exp_54_ram[236] = 0;
    exp_54_ram[237] = 127;
    exp_54_ram[238] = 0;
    exp_54_ram[239] = 255;
    exp_54_ram[240] = 0;
    exp_54_ram[241] = 0;
    exp_54_ram[242] = 0;
    exp_54_ram[243] = 0;
    exp_54_ram[244] = 0;
    exp_54_ram[245] = 0;
    exp_54_ram[246] = 0;
    exp_54_ram[247] = 0;
    exp_54_ram[248] = 0;
    exp_54_ram[249] = 0;
    exp_54_ram[250] = 254;
    exp_54_ram[251] = 255;
    exp_54_ram[252] = 0;
    exp_54_ram[253] = 0;
    exp_54_ram[254] = 219;
    exp_54_ram[255] = 0;
    exp_54_ram[256] = 0;
    exp_54_ram[257] = 252;
    exp_54_ram[258] = 0;
    exp_54_ram[259] = 0;
    exp_54_ram[260] = 0;
    exp_54_ram[261] = 0;
    exp_54_ram[262] = 0;
    exp_54_ram[263] = 1;
    exp_54_ram[264] = 0;
    exp_54_ram[265] = 254;
    exp_54_ram[266] = 0;
    exp_54_ram[267] = 2;
    exp_54_ram[268] = 0;
    exp_54_ram[269] = 254;
    exp_54_ram[270] = 254;
    exp_54_ram[271] = 254;
    exp_54_ram[272] = 254;
    exp_54_ram[273] = 0;
    exp_54_ram[274] = 1;
    exp_54_ram[275] = 2;
    exp_54_ram[276] = 0;
    exp_54_ram[277] = 254;
    exp_54_ram[278] = 0;
    exp_54_ram[279] = 0;
    exp_54_ram[280] = 2;
    exp_54_ram[281] = 0;
    exp_54_ram[282] = 254;
    exp_54_ram[283] = 254;
    exp_54_ram[284] = 254;
    exp_54_ram[285] = 254;
    exp_54_ram[286] = 254;
    exp_54_ram[287] = 0;
    exp_54_ram[288] = 254;
    exp_54_ram[289] = 0;
    exp_54_ram[290] = 31;
    exp_54_ram[291] = 0;
    exp_54_ram[292] = 1;
    exp_54_ram[293] = 1;
    exp_54_ram[294] = 2;
    exp_54_ram[295] = 0;
    exp_54_ram[296] = 253;
    exp_54_ram[297] = 2;
    exp_54_ram[298] = 3;
    exp_54_ram[299] = 252;
    exp_54_ram[300] = 252;
    exp_54_ram[301] = 253;
    exp_54_ram[302] = 254;
    exp_54_ram[303] = 1;
    exp_54_ram[304] = 254;
    exp_54_ram[305] = 0;
    exp_54_ram[306] = 254;
    exp_54_ram[307] = 254;
    exp_54_ram[308] = 0;
    exp_54_ram[309] = 0;
    exp_54_ram[310] = 253;
    exp_54_ram[311] = 255;
    exp_54_ram[312] = 252;
    exp_54_ram[313] = 252;
    exp_54_ram[314] = 254;
    exp_54_ram[315] = 253;
    exp_54_ram[316] = 64;
    exp_54_ram[317] = 0;
    exp_54_ram[318] = 2;
    exp_54_ram[319] = 3;
    exp_54_ram[320] = 0;
    exp_54_ram[321] = 254;
    exp_54_ram[322] = 0;
    exp_54_ram[323] = 2;
    exp_54_ram[324] = 0;
    exp_54_ram[325] = 254;
    exp_54_ram[326] = 254;
    exp_54_ram[327] = 2;
    exp_54_ram[328] = 0;
    exp_54_ram[329] = 254;
    exp_54_ram[330] = 3;
    exp_54_ram[331] = 0;
    exp_54_ram[332] = 0;
    exp_54_ram[333] = 0;
    exp_54_ram[334] = 0;
    exp_54_ram[335] = 0;
    exp_54_ram[336] = 15;
    exp_54_ram[337] = 0;
    exp_54_ram[338] = 1;
    exp_54_ram[339] = 2;
    exp_54_ram[340] = 0;
    exp_54_ram[341] = 253;
    exp_54_ram[342] = 2;
    exp_54_ram[343] = 2;
    exp_54_ram[344] = 3;
    exp_54_ram[345] = 252;
    exp_54_ram[346] = 254;
    exp_54_ram[347] = 4;
    exp_54_ram[348] = 254;
    exp_54_ram[349] = 0;
    exp_54_ram[350] = 0;
    exp_54_ram[351] = 0;
    exp_54_ram[352] = 0;
    exp_54_ram[353] = 0;
    exp_54_ram[354] = 253;
    exp_54_ram[355] = 0;
    exp_54_ram[356] = 0;
    exp_54_ram[357] = 253;
    exp_54_ram[358] = 0;
    exp_54_ram[359] = 0;
    exp_54_ram[360] = 0;
    exp_54_ram[361] = 253;
    exp_54_ram[362] = 254;
    exp_54_ram[363] = 253;
    exp_54_ram[364] = 0;
    exp_54_ram[365] = 0;
    exp_54_ram[366] = 0;
    exp_54_ram[367] = 244;
    exp_54_ram[368] = 0;
    exp_54_ram[369] = 250;
    exp_54_ram[370] = 254;
    exp_54_ram[371] = 0;
    exp_54_ram[372] = 2;
    exp_54_ram[373] = 2;
    exp_54_ram[374] = 3;
    exp_54_ram[375] = 0;
    exp_54_ram[376] = 252;
    exp_54_ram[377] = 2;
    exp_54_ram[378] = 2;
    exp_54_ram[379] = 4;
    exp_54_ram[380] = 252;
    exp_54_ram[381] = 252;
    exp_54_ram[382] = 252;
    exp_54_ram[383] = 252;
    exp_54_ram[384] = 252;
    exp_54_ram[385] = 252;
    exp_54_ram[386] = 253;
    exp_54_ram[387] = 253;
    exp_54_ram[388] = 253;
    exp_54_ram[389] = 254;
    exp_54_ram[390] = 252;
    exp_54_ram[391] = 0;
    exp_54_ram[392] = 8;
    exp_54_ram[393] = 252;
    exp_54_ram[394] = 0;
    exp_54_ram[395] = 8;
    exp_54_ram[396] = 252;
    exp_54_ram[397] = 254;
    exp_54_ram[398] = 3;
    exp_54_ram[399] = 253;
    exp_54_ram[400] = 0;
    exp_54_ram[401] = 252;
    exp_54_ram[402] = 253;
    exp_54_ram[403] = 253;
    exp_54_ram[404] = 0;
    exp_54_ram[405] = 253;
    exp_54_ram[406] = 2;
    exp_54_ram[407] = 0;
    exp_54_ram[408] = 254;
    exp_54_ram[409] = 0;
    exp_54_ram[410] = 254;
    exp_54_ram[411] = 254;
    exp_54_ram[412] = 252;
    exp_54_ram[413] = 252;
    exp_54_ram[414] = 4;
    exp_54_ram[415] = 252;
    exp_54_ram[416] = 255;
    exp_54_ram[417] = 252;
    exp_54_ram[418] = 252;
    exp_54_ram[419] = 252;
    exp_54_ram[420] = 0;
    exp_54_ram[421] = 0;
    exp_54_ram[422] = 253;
    exp_54_ram[423] = 0;
    exp_54_ram[424] = 252;
    exp_54_ram[425] = 253;
    exp_54_ram[426] = 253;
    exp_54_ram[427] = 0;
    exp_54_ram[428] = 253;
    exp_54_ram[429] = 0;
    exp_54_ram[430] = 252;
    exp_54_ram[431] = 252;
    exp_54_ram[432] = 252;
    exp_54_ram[433] = 0;
    exp_54_ram[434] = 4;
    exp_54_ram[435] = 2;
    exp_54_ram[436] = 253;
    exp_54_ram[437] = 0;
    exp_54_ram[438] = 252;
    exp_54_ram[439] = 253;
    exp_54_ram[440] = 253;
    exp_54_ram[441] = 0;
    exp_54_ram[442] = 253;
    exp_54_ram[443] = 2;
    exp_54_ram[444] = 0;
    exp_54_ram[445] = 253;
    exp_54_ram[446] = 254;
    exp_54_ram[447] = 64;
    exp_54_ram[448] = 252;
    exp_54_ram[449] = 252;
    exp_54_ram[450] = 253;
    exp_54_ram[451] = 0;
    exp_54_ram[452] = 3;
    exp_54_ram[453] = 3;
    exp_54_ram[454] = 4;
    exp_54_ram[455] = 0;
    exp_54_ram[456] = 253;
    exp_54_ram[457] = 2;
    exp_54_ram[458] = 2;
    exp_54_ram[459] = 3;
    exp_54_ram[460] = 254;
    exp_54_ram[461] = 254;
    exp_54_ram[462] = 254;
    exp_54_ram[463] = 254;
    exp_54_ram[464] = 252;
    exp_54_ram[465] = 252;
    exp_54_ram[466] = 0;
    exp_54_ram[467] = 253;
    exp_54_ram[468] = 252;
    exp_54_ram[469] = 0;
    exp_54_ram[470] = 0;
    exp_54_ram[471] = 10;
    exp_54_ram[472] = 0;
    exp_54_ram[473] = 4;
    exp_54_ram[474] = 0;
    exp_54_ram[475] = 0;
    exp_54_ram[476] = 4;
    exp_54_ram[477] = 253;
    exp_54_ram[478] = 0;
    exp_54_ram[479] = 0;
    exp_54_ram[480] = 0;
    exp_54_ram[481] = 2;
    exp_54_ram[482] = 0;
    exp_54_ram[483] = 255;
    exp_54_ram[484] = 0;
    exp_54_ram[485] = 2;
    exp_54_ram[486] = 253;
    exp_54_ram[487] = 0;
    exp_54_ram[488] = 252;
    exp_54_ram[489] = 253;
    exp_54_ram[490] = 0;
    exp_54_ram[491] = 3;
    exp_54_ram[492] = 0;
    exp_54_ram[493] = 253;
    exp_54_ram[494] = 0;
    exp_54_ram[495] = 2;
    exp_54_ram[496] = 253;
    exp_54_ram[497] = 1;
    exp_54_ram[498] = 252;
    exp_54_ram[499] = 2;
    exp_54_ram[500] = 253;
    exp_54_ram[501] = 0;
    exp_54_ram[502] = 252;
    exp_54_ram[503] = 253;
    exp_54_ram[504] = 0;
    exp_54_ram[505] = 3;
    exp_54_ram[506] = 0;
    exp_54_ram[507] = 0;
    exp_54_ram[508] = 0;
    exp_54_ram[509] = 0;
    exp_54_ram[510] = 253;
    exp_54_ram[511] = 0;
    exp_54_ram[512] = 0;
    exp_54_ram[513] = 253;
    exp_54_ram[514] = 1;
    exp_54_ram[515] = 252;
    exp_54_ram[516] = 0;
    exp_54_ram[517] = 1;
    exp_54_ram[518] = 20;
    exp_54_ram[519] = 0;
    exp_54_ram[520] = 64;
    exp_54_ram[521] = 4;
    exp_54_ram[522] = 253;
    exp_54_ram[523] = 4;
    exp_54_ram[524] = 253;
    exp_54_ram[525] = 0;
    exp_54_ram[526] = 0;
    exp_54_ram[527] = 253;
    exp_54_ram[528] = 0;
    exp_54_ram[529] = 2;
    exp_54_ram[530] = 253;
    exp_54_ram[531] = 255;
    exp_54_ram[532] = 252;
    exp_54_ram[533] = 253;
    exp_54_ram[534] = 0;
    exp_54_ram[535] = 253;
    exp_54_ram[536] = 1;
    exp_54_ram[537] = 0;
    exp_54_ram[538] = 253;
    exp_54_ram[539] = 255;
    exp_54_ram[540] = 252;
    exp_54_ram[541] = 253;
    exp_54_ram[542] = 1;
    exp_54_ram[543] = 2;
    exp_54_ram[544] = 0;
    exp_54_ram[545] = 2;
    exp_54_ram[546] = 2;
    exp_54_ram[547] = 253;
    exp_54_ram[548] = 1;
    exp_54_ram[549] = 2;
    exp_54_ram[550] = 253;
    exp_54_ram[551] = 0;
    exp_54_ram[552] = 252;
    exp_54_ram[553] = 253;
    exp_54_ram[554] = 0;
    exp_54_ram[555] = 7;
    exp_54_ram[556] = 0;
    exp_54_ram[557] = 7;
    exp_54_ram[558] = 253;
    exp_54_ram[559] = 1;
    exp_54_ram[560] = 2;
    exp_54_ram[561] = 0;
    exp_54_ram[562] = 2;
    exp_54_ram[563] = 2;
    exp_54_ram[564] = 253;
    exp_54_ram[565] = 1;
    exp_54_ram[566] = 2;
    exp_54_ram[567] = 253;
    exp_54_ram[568] = 0;
    exp_54_ram[569] = 252;
    exp_54_ram[570] = 253;
    exp_54_ram[571] = 0;
    exp_54_ram[572] = 5;
    exp_54_ram[573] = 0;
    exp_54_ram[574] = 3;
    exp_54_ram[575] = 253;
    exp_54_ram[576] = 0;
    exp_54_ram[577] = 2;
    exp_54_ram[578] = 253;
    exp_54_ram[579] = 1;
    exp_54_ram[580] = 2;
    exp_54_ram[581] = 253;
    exp_54_ram[582] = 0;
    exp_54_ram[583] = 252;
    exp_54_ram[584] = 253;
    exp_54_ram[585] = 0;
    exp_54_ram[586] = 6;
    exp_54_ram[587] = 0;
    exp_54_ram[588] = 253;
    exp_54_ram[589] = 1;
    exp_54_ram[590] = 2;
    exp_54_ram[591] = 253;
    exp_54_ram[592] = 0;
    exp_54_ram[593] = 252;
    exp_54_ram[594] = 253;
    exp_54_ram[595] = 0;
    exp_54_ram[596] = 3;
    exp_54_ram[597] = 0;
    exp_54_ram[598] = 253;
    exp_54_ram[599] = 1;
    exp_54_ram[600] = 8;
    exp_54_ram[601] = 253;
    exp_54_ram[602] = 2;
    exp_54_ram[603] = 253;
    exp_54_ram[604] = 0;
    exp_54_ram[605] = 252;
    exp_54_ram[606] = 253;
    exp_54_ram[607] = 0;
    exp_54_ram[608] = 2;
    exp_54_ram[609] = 0;
    exp_54_ram[610] = 5;
    exp_54_ram[611] = 0;
    exp_54_ram[612] = 0;
    exp_54_ram[613] = 2;
    exp_54_ram[614] = 253;
    exp_54_ram[615] = 0;
    exp_54_ram[616] = 252;
    exp_54_ram[617] = 253;
    exp_54_ram[618] = 0;
    exp_54_ram[619] = 2;
    exp_54_ram[620] = 0;
    exp_54_ram[621] = 2;
    exp_54_ram[622] = 0;
    exp_54_ram[623] = 0;
    exp_54_ram[624] = 2;
    exp_54_ram[625] = 253;
    exp_54_ram[626] = 0;
    exp_54_ram[627] = 252;
    exp_54_ram[628] = 253;
    exp_54_ram[629] = 0;
    exp_54_ram[630] = 2;
    exp_54_ram[631] = 0;
    exp_54_ram[632] = 0;
    exp_54_ram[633] = 0;
    exp_54_ram[634] = 253;
    exp_54_ram[635] = 253;
    exp_54_ram[636] = 254;
    exp_54_ram[637] = 254;
    exp_54_ram[638] = 254;
    exp_54_ram[639] = 254;
    exp_54_ram[640] = 190;
    exp_54_ram[641] = 0;
    exp_54_ram[642] = 0;
    exp_54_ram[643] = 2;
    exp_54_ram[644] = 2;
    exp_54_ram[645] = 3;
    exp_54_ram[646] = 0;
    exp_54_ram[647] = 249;
    exp_54_ram[648] = 6;
    exp_54_ram[649] = 6;
    exp_54_ram[650] = 7;
    exp_54_ram[651] = 250;
    exp_54_ram[652] = 250;
    exp_54_ram[653] = 250;
    exp_54_ram[654] = 250;
    exp_54_ram[655] = 250;
    exp_54_ram[656] = 251;
    exp_54_ram[657] = 251;
    exp_54_ram[658] = 250;
    exp_54_ram[659] = 254;
    exp_54_ram[660] = 250;
    exp_54_ram[661] = 0;
    exp_54_ram[662] = 0;
    exp_54_ram[663] = 254;
    exp_54_ram[664] = 0;
    exp_54_ram[665] = 0;
    exp_54_ram[666] = 64;
    exp_54_ram[667] = 0;
    exp_54_ram[668] = 250;
    exp_54_ram[669] = 8;
    exp_54_ram[670] = 250;
    exp_54_ram[671] = 250;
    exp_54_ram[672] = 2;
    exp_54_ram[673] = 254;
    exp_54_ram[674] = 254;
    exp_54_ram[675] = 0;
    exp_54_ram[676] = 0;
    exp_54_ram[677] = 254;
    exp_54_ram[678] = 3;
    exp_54_ram[679] = 15;
    exp_54_ram[680] = 3;
    exp_54_ram[681] = 0;
    exp_54_ram[682] = 2;
    exp_54_ram[683] = 0;
    exp_54_ram[684] = 4;
    exp_54_ram[685] = 0;
    exp_54_ram[686] = 6;
    exp_54_ram[687] = 254;
    exp_54_ram[688] = 0;
    exp_54_ram[689] = 15;
    exp_54_ram[690] = 255;
    exp_54_ram[691] = 15;
    exp_54_ram[692] = 254;
    exp_54_ram[693] = 0;
    exp_54_ram[694] = 254;
    exp_54_ram[695] = 255;
    exp_54_ram[696] = 0;
    exp_54_ram[697] = 252;
    exp_54_ram[698] = 250;
    exp_54_ram[699] = 250;
    exp_54_ram[700] = 2;
    exp_54_ram[701] = 250;
    exp_54_ram[702] = 250;
    exp_54_ram[703] = 0;
    exp_54_ram[704] = 254;
    exp_54_ram[705] = 1;
    exp_54_ram[706] = 246;
    exp_54_ram[707] = 250;
    exp_54_ram[708] = 252;
    exp_54_ram[709] = 0;
    exp_54_ram[710] = 0;
    exp_54_ram[711] = 0;
    exp_54_ram[712] = 0;
    exp_54_ram[713] = 250;
    exp_54_ram[714] = 0;
    exp_54_ram[715] = 250;
    exp_54_ram[716] = 0;
    exp_54_ram[717] = 254;
    exp_54_ram[718] = 251;
    exp_54_ram[719] = 251;
    exp_54_ram[720] = 251;
    exp_54_ram[721] = 251;
    exp_54_ram[722] = 189;
    exp_54_ram[723] = 0;
    exp_54_ram[724] = 0;
    exp_54_ram[725] = 6;
    exp_54_ram[726] = 6;
    exp_54_ram[727] = 7;
    exp_54_ram[728] = 0;
    exp_54_ram[729] = 248;
    exp_54_ram[730] = 6;
    exp_54_ram[731] = 6;
    exp_54_ram[732] = 8;
    exp_54_ram[733] = 250;
    exp_54_ram[734] = 250;
    exp_54_ram[735] = 250;
    exp_54_ram[736] = 250;
    exp_54_ram[737] = 248;
    exp_54_ram[738] = 252;
    exp_54_ram[739] = 250;
    exp_54_ram[740] = 32;
    exp_54_ram[741] = 66;
    exp_54_ram[742] = 250;
    exp_54_ram[743] = 32;
    exp_54_ram[744] = 250;
    exp_54_ram[745] = 0;
    exp_54_ram[746] = 2;
    exp_54_ram[747] = 2;
    exp_54_ram[748] = 250;
    exp_54_ram[749] = 0;
    exp_54_ram[750] = 253;
    exp_54_ram[751] = 0;
    exp_54_ram[752] = 252;
    exp_54_ram[753] = 250;
    exp_54_ram[754] = 250;
    exp_54_ram[755] = 0;
    exp_54_ram[756] = 250;
    exp_54_ram[757] = 0;
    exp_54_ram[758] = 250;
    exp_54_ram[759] = 0;
    exp_54_ram[760] = 250;
    exp_54_ram[761] = 28;
    exp_54_ram[762] = 250;
    exp_54_ram[763] = 0;
    exp_54_ram[764] = 250;
    exp_54_ram[765] = 254;
    exp_54_ram[766] = 250;
    exp_54_ram[767] = 0;
    exp_54_ram[768] = 254;
    exp_54_ram[769] = 1;
    exp_54_ram[770] = 12;
    exp_54_ram[771] = 0;
    exp_54_ram[772] = 0;
    exp_54_ram[773] = 220;
    exp_54_ram[774] = 0;
    exp_54_ram[775] = 0;
    exp_54_ram[776] = 0;
    exp_54_ram[777] = 254;
    exp_54_ram[778] = 0;
    exp_54_ram[779] = 254;
    exp_54_ram[780] = 250;
    exp_54_ram[781] = 0;
    exp_54_ram[782] = 250;
    exp_54_ram[783] = 0;
    exp_54_ram[784] = 254;
    exp_54_ram[785] = 9;
    exp_54_ram[786] = 254;
    exp_54_ram[787] = 0;
    exp_54_ram[788] = 254;
    exp_54_ram[789] = 250;
    exp_54_ram[790] = 0;
    exp_54_ram[791] = 250;
    exp_54_ram[792] = 0;
    exp_54_ram[793] = 254;
    exp_54_ram[794] = 7;
    exp_54_ram[795] = 254;
    exp_54_ram[796] = 0;
    exp_54_ram[797] = 254;
    exp_54_ram[798] = 250;
    exp_54_ram[799] = 0;
    exp_54_ram[800] = 250;
    exp_54_ram[801] = 0;
    exp_54_ram[802] = 254;
    exp_54_ram[803] = 5;
    exp_54_ram[804] = 254;
    exp_54_ram[805] = 0;
    exp_54_ram[806] = 254;
    exp_54_ram[807] = 250;
    exp_54_ram[808] = 0;
    exp_54_ram[809] = 250;
    exp_54_ram[810] = 0;
    exp_54_ram[811] = 254;
    exp_54_ram[812] = 3;
    exp_54_ram[813] = 254;
    exp_54_ram[814] = 1;
    exp_54_ram[815] = 254;
    exp_54_ram[816] = 250;
    exp_54_ram[817] = 0;
    exp_54_ram[818] = 250;
    exp_54_ram[819] = 0;
    exp_54_ram[820] = 254;
    exp_54_ram[821] = 0;
    exp_54_ram[822] = 254;
    exp_54_ram[823] = 0;
    exp_54_ram[824] = 254;
    exp_54_ram[825] = 240;
    exp_54_ram[826] = 254;
    exp_54_ram[827] = 250;
    exp_54_ram[828] = 0;
    exp_54_ram[829] = 0;
    exp_54_ram[830] = 128;
    exp_54_ram[831] = 0;
    exp_54_ram[832] = 0;
    exp_54_ram[833] = 250;
    exp_54_ram[834] = 0;
    exp_54_ram[835] = 132;
    exp_54_ram[836] = 254;
    exp_54_ram[837] = 6;
    exp_54_ram[838] = 250;
    exp_54_ram[839] = 0;
    exp_54_ram[840] = 2;
    exp_54_ram[841] = 4;
    exp_54_ram[842] = 249;
    exp_54_ram[843] = 0;
    exp_54_ram[844] = 248;
    exp_54_ram[845] = 0;
    exp_54_ram[846] = 252;
    exp_54_ram[847] = 252;
    exp_54_ram[848] = 2;
    exp_54_ram[849] = 254;
    exp_54_ram[850] = 0;
    exp_54_ram[851] = 254;
    exp_54_ram[852] = 252;
    exp_54_ram[853] = 64;
    exp_54_ram[854] = 254;
    exp_54_ram[855] = 0;
    exp_54_ram[856] = 252;
    exp_54_ram[857] = 254;
    exp_54_ram[858] = 250;
    exp_54_ram[859] = 0;
    exp_54_ram[860] = 250;
    exp_54_ram[861] = 254;
    exp_54_ram[862] = 250;
    exp_54_ram[863] = 0;
    exp_54_ram[864] = 2;
    exp_54_ram[865] = 8;
    exp_54_ram[866] = 254;
    exp_54_ram[867] = 64;
    exp_54_ram[868] = 254;
    exp_54_ram[869] = 250;
    exp_54_ram[870] = 0;
    exp_54_ram[871] = 250;
    exp_54_ram[872] = 250;
    exp_54_ram[873] = 0;
    exp_54_ram[874] = 0;
    exp_54_ram[875] = 245;
    exp_54_ram[876] = 0;
    exp_54_ram[877] = 0;
    exp_54_ram[878] = 250;
    exp_54_ram[879] = 0;
    exp_54_ram[880] = 249;
    exp_54_ram[881] = 254;
    exp_54_ram[882] = 4;
    exp_54_ram[883] = 250;
    exp_54_ram[884] = 0;
    exp_54_ram[885] = 2;
    exp_54_ram[886] = 2;
    exp_54_ram[887] = 249;
    exp_54_ram[888] = 0;
    exp_54_ram[889] = 248;
    exp_54_ram[890] = 0;
    exp_54_ram[891] = 252;
    exp_54_ram[892] = 252;
    exp_54_ram[893] = 0;
    exp_54_ram[894] = 0;
    exp_54_ram[895] = 254;
    exp_54_ram[896] = 250;
    exp_54_ram[897] = 0;
    exp_54_ram[898] = 250;
    exp_54_ram[899] = 250;
    exp_54_ram[900] = 0;
    exp_54_ram[901] = 249;
    exp_54_ram[902] = 1;
    exp_54_ram[903] = 14;
    exp_54_ram[904] = 0;
    exp_54_ram[905] = 0;
    exp_54_ram[906] = 224;
    exp_54_ram[907] = 0;
    exp_54_ram[908] = 0;
    exp_54_ram[909] = 0;
    exp_54_ram[910] = 254;
    exp_54_ram[911] = 16;
    exp_54_ram[912] = 254;
    exp_54_ram[913] = 250;
    exp_54_ram[914] = 0;
    exp_54_ram[915] = 250;
    exp_54_ram[916] = 250;
    exp_54_ram[917] = 0;
    exp_54_ram[918] = 6;
    exp_54_ram[919] = 12;
    exp_54_ram[920] = 254;
    exp_54_ram[921] = 32;
    exp_54_ram[922] = 254;
    exp_54_ram[923] = 250;
    exp_54_ram[924] = 0;
    exp_54_ram[925] = 250;
    exp_54_ram[926] = 10;
    exp_54_ram[927] = 254;
    exp_54_ram[928] = 8;
    exp_54_ram[929] = 254;
    exp_54_ram[930] = 250;
    exp_54_ram[931] = 0;
    exp_54_ram[932] = 250;
    exp_54_ram[933] = 250;
    exp_54_ram[934] = 0;
    exp_54_ram[935] = 6;
    exp_54_ram[936] = 8;
    exp_54_ram[937] = 254;
    exp_54_ram[938] = 4;
    exp_54_ram[939] = 254;
    exp_54_ram[940] = 250;
    exp_54_ram[941] = 0;
    exp_54_ram[942] = 250;
    exp_54_ram[943] = 6;
    exp_54_ram[944] = 254;
    exp_54_ram[945] = 16;
    exp_54_ram[946] = 254;
    exp_54_ram[947] = 250;
    exp_54_ram[948] = 0;
    exp_54_ram[949] = 250;
    exp_54_ram[950] = 5;
    exp_54_ram[951] = 254;
    exp_54_ram[952] = 32;
    exp_54_ram[953] = 254;
    exp_54_ram[954] = 250;
    exp_54_ram[955] = 0;
    exp_54_ram[956] = 250;
    exp_54_ram[957] = 3;
    exp_54_ram[958] = 254;
    exp_54_ram[959] = 16;
    exp_54_ram[960] = 254;
    exp_54_ram[961] = 250;
    exp_54_ram[962] = 0;
    exp_54_ram[963] = 250;
    exp_54_ram[964] = 1;
    exp_54_ram[965] = 0;
    exp_54_ram[966] = 1;
    exp_54_ram[967] = 0;
    exp_54_ram[968] = 0;
    exp_54_ram[969] = 0;
    exp_54_ram[970] = 250;
    exp_54_ram[971] = 0;
    exp_54_ram[972] = 253;
    exp_54_ram[973] = 5;
    exp_54_ram[974] = 98;
    exp_54_ram[975] = 0;
    exp_54_ram[976] = 0;
    exp_54_ram[977] = 229;
    exp_54_ram[978] = 0;
    exp_54_ram[979] = 0;
    exp_54_ram[980] = 0;
    exp_54_ram[981] = 250;
    exp_54_ram[982] = 0;
    exp_54_ram[983] = 7;
    exp_54_ram[984] = 0;
    exp_54_ram[985] = 250;
    exp_54_ram[986] = 0;
    exp_54_ram[987] = 5;
    exp_54_ram[988] = 0;
    exp_54_ram[989] = 1;
    exp_54_ram[990] = 252;
    exp_54_ram[991] = 5;
    exp_54_ram[992] = 250;
    exp_54_ram[993] = 0;
    exp_54_ram[994] = 6;
    exp_54_ram[995] = 0;
    exp_54_ram[996] = 0;
    exp_54_ram[997] = 252;
    exp_54_ram[998] = 3;
    exp_54_ram[999] = 250;
    exp_54_ram[1000] = 0;
    exp_54_ram[1001] = 6;
    exp_54_ram[1002] = 0;
    exp_54_ram[1003] = 0;
    exp_54_ram[1004] = 252;
    exp_54_ram[1005] = 1;
    exp_54_ram[1006] = 0;
    exp_54_ram[1007] = 252;
    exp_54_ram[1008] = 254;
    exp_54_ram[1009] = 254;
    exp_54_ram[1010] = 254;
    exp_54_ram[1011] = 250;
    exp_54_ram[1012] = 0;
    exp_54_ram[1013] = 5;
    exp_54_ram[1014] = 0;
    exp_54_ram[1015] = 254;
    exp_54_ram[1016] = 2;
    exp_54_ram[1017] = 254;
    exp_54_ram[1018] = 250;
    exp_54_ram[1019] = 0;
    exp_54_ram[1020] = 6;
    exp_54_ram[1021] = 2;
    exp_54_ram[1022] = 250;
    exp_54_ram[1023] = 0;
    exp_54_ram[1024] = 6;
    exp_54_ram[1025] = 0;
    exp_54_ram[1026] = 254;
    exp_54_ram[1027] = 255;
    exp_54_ram[1028] = 254;
    exp_54_ram[1029] = 254;
    exp_54_ram[1030] = 64;
    exp_54_ram[1031] = 0;
    exp_54_ram[1032] = 254;
    exp_54_ram[1033] = 255;
    exp_54_ram[1034] = 254;
    exp_54_ram[1035] = 250;
    exp_54_ram[1036] = 0;
    exp_54_ram[1037] = 6;
    exp_54_ram[1038] = 0;
    exp_54_ram[1039] = 250;
    exp_54_ram[1040] = 0;
    exp_54_ram[1041] = 6;
    exp_54_ram[1042] = 20;
    exp_54_ram[1043] = 254;
    exp_54_ram[1044] = 32;
    exp_54_ram[1045] = 34;
    exp_54_ram[1046] = 254;
    exp_54_ram[1047] = 16;
    exp_54_ram[1048] = 6;
    exp_54_ram[1049] = 249;
    exp_54_ram[1050] = 0;
    exp_54_ram[1051] = 248;
    exp_54_ram[1052] = 0;
    exp_54_ram[1053] = 250;
    exp_54_ram[1054] = 251;
    exp_54_ram[1055] = 65;
    exp_54_ram[1056] = 251;
    exp_54_ram[1057] = 0;
    exp_54_ram[1058] = 64;
    exp_54_ram[1059] = 0;
    exp_54_ram[1060] = 251;
    exp_54_ram[1061] = 1;
    exp_54_ram[1062] = 15;
    exp_54_ram[1063] = 254;
    exp_54_ram[1064] = 0;
    exp_54_ram[1065] = 254;
    exp_54_ram[1066] = 0;
    exp_54_ram[1067] = 254;
    exp_54_ram[1068] = 253;
    exp_54_ram[1069] = 0;
    exp_54_ram[1070] = 0;
    exp_54_ram[1071] = 250;
    exp_54_ram[1072] = 253;
    exp_54_ram[1073] = 250;
    exp_54_ram[1074] = 250;
    exp_54_ram[1075] = 149;
    exp_54_ram[1076] = 252;
    exp_54_ram[1077] = 27;
    exp_54_ram[1078] = 254;
    exp_54_ram[1079] = 4;
    exp_54_ram[1080] = 0;
    exp_54_ram[1081] = 249;
    exp_54_ram[1082] = 0;
    exp_54_ram[1083] = 248;
    exp_54_ram[1084] = 0;
    exp_54_ram[1085] = 15;
    exp_54_ram[1086] = 3;
    exp_54_ram[1087] = 254;
    exp_54_ram[1088] = 8;
    exp_54_ram[1089] = 2;
    exp_54_ram[1090] = 249;
    exp_54_ram[1091] = 0;
    exp_54_ram[1092] = 248;
    exp_54_ram[1093] = 0;
    exp_54_ram[1094] = 1;
    exp_54_ram[1095] = 65;
    exp_54_ram[1096] = 1;
    exp_54_ram[1097] = 249;
    exp_54_ram[1098] = 0;
    exp_54_ram[1099] = 248;
    exp_54_ram[1100] = 0;
    exp_54_ram[1101] = 250;
    exp_54_ram[1102] = 251;
    exp_54_ram[1103] = 65;
    exp_54_ram[1104] = 251;
    exp_54_ram[1105] = 0;
    exp_54_ram[1106] = 64;
    exp_54_ram[1107] = 0;
    exp_54_ram[1108] = 251;
    exp_54_ram[1109] = 1;
    exp_54_ram[1110] = 15;
    exp_54_ram[1111] = 254;
    exp_54_ram[1112] = 0;
    exp_54_ram[1113] = 254;
    exp_54_ram[1114] = 0;
    exp_54_ram[1115] = 254;
    exp_54_ram[1116] = 253;
    exp_54_ram[1117] = 0;
    exp_54_ram[1118] = 0;
    exp_54_ram[1119] = 250;
    exp_54_ram[1120] = 253;
    exp_54_ram[1121] = 250;
    exp_54_ram[1122] = 250;
    exp_54_ram[1123] = 137;
    exp_54_ram[1124] = 252;
    exp_54_ram[1125] = 15;
    exp_54_ram[1126] = 254;
    exp_54_ram[1127] = 32;
    exp_54_ram[1128] = 14;
    exp_54_ram[1129] = 254;
    exp_54_ram[1130] = 16;
    exp_54_ram[1131] = 4;
    exp_54_ram[1132] = 249;
    exp_54_ram[1133] = 0;
    exp_54_ram[1134] = 248;
    exp_54_ram[1135] = 0;
    exp_54_ram[1136] = 254;
    exp_54_ram[1137] = 0;
    exp_54_ram[1138] = 254;
    exp_54_ram[1139] = 0;
    exp_54_ram[1140] = 254;
    exp_54_ram[1141] = 253;
    exp_54_ram[1142] = 0;
    exp_54_ram[1143] = 250;
    exp_54_ram[1144] = 253;
    exp_54_ram[1145] = 250;
    exp_54_ram[1146] = 250;
    exp_54_ram[1147] = 131;
    exp_54_ram[1148] = 252;
    exp_54_ram[1149] = 9;
    exp_54_ram[1150] = 254;
    exp_54_ram[1151] = 4;
    exp_54_ram[1152] = 0;
    exp_54_ram[1153] = 249;
    exp_54_ram[1154] = 0;
    exp_54_ram[1155] = 248;
    exp_54_ram[1156] = 0;
    exp_54_ram[1157] = 15;
    exp_54_ram[1158] = 3;
    exp_54_ram[1159] = 254;
    exp_54_ram[1160] = 8;
    exp_54_ram[1161] = 2;
    exp_54_ram[1162] = 249;
    exp_54_ram[1163] = 0;
    exp_54_ram[1164] = 248;
    exp_54_ram[1165] = 0;
    exp_54_ram[1166] = 1;
    exp_54_ram[1167] = 1;
    exp_54_ram[1168] = 1;
    exp_54_ram[1169] = 249;
    exp_54_ram[1170] = 0;
    exp_54_ram[1171] = 248;
    exp_54_ram[1172] = 0;
    exp_54_ram[1173] = 252;
    exp_54_ram[1174] = 254;
    exp_54_ram[1175] = 0;
    exp_54_ram[1176] = 254;
    exp_54_ram[1177] = 0;
    exp_54_ram[1178] = 254;
    exp_54_ram[1179] = 253;
    exp_54_ram[1180] = 0;
    exp_54_ram[1181] = 252;
    exp_54_ram[1182] = 250;
    exp_54_ram[1183] = 253;
    exp_54_ram[1184] = 250;
    exp_54_ram[1185] = 250;
    exp_54_ram[1186] = 249;
    exp_54_ram[1187] = 252;
    exp_54_ram[1188] = 250;
    exp_54_ram[1189] = 0;
    exp_54_ram[1190] = 250;
    exp_54_ram[1191] = 48;
    exp_54_ram[1192] = 0;
    exp_54_ram[1193] = 252;
    exp_54_ram[1194] = 254;
    exp_54_ram[1195] = 0;
    exp_54_ram[1196] = 4;
    exp_54_ram[1197] = 2;
    exp_54_ram[1198] = 253;
    exp_54_ram[1199] = 0;
    exp_54_ram[1200] = 252;
    exp_54_ram[1201] = 250;
    exp_54_ram[1202] = 250;
    exp_54_ram[1203] = 0;
    exp_54_ram[1204] = 250;
    exp_54_ram[1205] = 2;
    exp_54_ram[1206] = 0;
    exp_54_ram[1207] = 253;
    exp_54_ram[1208] = 0;
    exp_54_ram[1209] = 252;
    exp_54_ram[1210] = 254;
    exp_54_ram[1211] = 252;
    exp_54_ram[1212] = 249;
    exp_54_ram[1213] = 0;
    exp_54_ram[1214] = 248;
    exp_54_ram[1215] = 0;
    exp_54_ram[1216] = 15;
    exp_54_ram[1217] = 253;
    exp_54_ram[1218] = 0;
    exp_54_ram[1219] = 252;
    exp_54_ram[1220] = 250;
    exp_54_ram[1221] = 250;
    exp_54_ram[1222] = 0;
    exp_54_ram[1223] = 250;
    exp_54_ram[1224] = 0;
    exp_54_ram[1225] = 254;
    exp_54_ram[1226] = 0;
    exp_54_ram[1227] = 4;
    exp_54_ram[1228] = 2;
    exp_54_ram[1229] = 253;
    exp_54_ram[1230] = 0;
    exp_54_ram[1231] = 252;
    exp_54_ram[1232] = 250;
    exp_54_ram[1233] = 250;
    exp_54_ram[1234] = 0;
    exp_54_ram[1235] = 250;
    exp_54_ram[1236] = 2;
    exp_54_ram[1237] = 0;
    exp_54_ram[1238] = 253;
    exp_54_ram[1239] = 0;
    exp_54_ram[1240] = 252;
    exp_54_ram[1241] = 254;
    exp_54_ram[1242] = 252;
    exp_54_ram[1243] = 250;
    exp_54_ram[1244] = 0;
    exp_54_ram[1245] = 250;
    exp_54_ram[1246] = 35;
    exp_54_ram[1247] = 249;
    exp_54_ram[1248] = 0;
    exp_54_ram[1249] = 248;
    exp_54_ram[1250] = 0;
    exp_54_ram[1251] = 252;
    exp_54_ram[1252] = 254;
    exp_54_ram[1253] = 0;
    exp_54_ram[1254] = 254;
    exp_54_ram[1255] = 0;
    exp_54_ram[1256] = 255;
    exp_54_ram[1257] = 0;
    exp_54_ram[1258] = 253;
    exp_54_ram[1259] = 143;
    exp_54_ram[1260] = 252;
    exp_54_ram[1261] = 254;
    exp_54_ram[1262] = 64;
    exp_54_ram[1263] = 0;
    exp_54_ram[1264] = 252;
    exp_54_ram[1265] = 254;
    exp_54_ram[1266] = 0;
    exp_54_ram[1267] = 0;
    exp_54_ram[1268] = 252;
    exp_54_ram[1269] = 254;
    exp_54_ram[1270] = 0;
    exp_54_ram[1271] = 6;
    exp_54_ram[1272] = 2;
    exp_54_ram[1273] = 253;
    exp_54_ram[1274] = 0;
    exp_54_ram[1275] = 252;
    exp_54_ram[1276] = 250;
    exp_54_ram[1277] = 250;
    exp_54_ram[1278] = 0;
    exp_54_ram[1279] = 250;
    exp_54_ram[1280] = 2;
    exp_54_ram[1281] = 0;
    exp_54_ram[1282] = 252;
    exp_54_ram[1283] = 0;
    exp_54_ram[1284] = 252;
    exp_54_ram[1285] = 254;
    exp_54_ram[1286] = 252;
    exp_54_ram[1287] = 3;
    exp_54_ram[1288] = 253;
    exp_54_ram[1289] = 0;
    exp_54_ram[1290] = 252;
    exp_54_ram[1291] = 0;
    exp_54_ram[1292] = 253;
    exp_54_ram[1293] = 0;
    exp_54_ram[1294] = 252;
    exp_54_ram[1295] = 250;
    exp_54_ram[1296] = 250;
    exp_54_ram[1297] = 0;
    exp_54_ram[1298] = 250;
    exp_54_ram[1299] = 0;
    exp_54_ram[1300] = 253;
    exp_54_ram[1301] = 0;
    exp_54_ram[1302] = 2;
    exp_54_ram[1303] = 254;
    exp_54_ram[1304] = 64;
    exp_54_ram[1305] = 250;
    exp_54_ram[1306] = 254;
    exp_54_ram[1307] = 255;
    exp_54_ram[1308] = 254;
    exp_54_ram[1309] = 250;
    exp_54_ram[1310] = 254;
    exp_54_ram[1311] = 0;
    exp_54_ram[1312] = 4;
    exp_54_ram[1313] = 2;
    exp_54_ram[1314] = 253;
    exp_54_ram[1315] = 0;
    exp_54_ram[1316] = 252;
    exp_54_ram[1317] = 250;
    exp_54_ram[1318] = 250;
    exp_54_ram[1319] = 0;
    exp_54_ram[1320] = 250;
    exp_54_ram[1321] = 2;
    exp_54_ram[1322] = 0;
    exp_54_ram[1323] = 252;
    exp_54_ram[1324] = 0;
    exp_54_ram[1325] = 252;
    exp_54_ram[1326] = 254;
    exp_54_ram[1327] = 252;
    exp_54_ram[1328] = 250;
    exp_54_ram[1329] = 0;
    exp_54_ram[1330] = 250;
    exp_54_ram[1331] = 13;
    exp_54_ram[1332] = 0;
    exp_54_ram[1333] = 254;
    exp_54_ram[1334] = 254;
    exp_54_ram[1335] = 2;
    exp_54_ram[1336] = 254;
    exp_54_ram[1337] = 249;
    exp_54_ram[1338] = 0;
    exp_54_ram[1339] = 248;
    exp_54_ram[1340] = 0;
    exp_54_ram[1341] = 0;
    exp_54_ram[1342] = 254;
    exp_54_ram[1343] = 0;
    exp_54_ram[1344] = 254;
    exp_54_ram[1345] = 0;
    exp_54_ram[1346] = 254;
    exp_54_ram[1347] = 1;
    exp_54_ram[1348] = 0;
    exp_54_ram[1349] = 250;
    exp_54_ram[1350] = 253;
    exp_54_ram[1351] = 250;
    exp_54_ram[1352] = 250;
    exp_54_ram[1353] = 207;
    exp_54_ram[1354] = 252;
    exp_54_ram[1355] = 250;
    exp_54_ram[1356] = 0;
    exp_54_ram[1357] = 250;
    exp_54_ram[1358] = 7;
    exp_54_ram[1359] = 253;
    exp_54_ram[1360] = 0;
    exp_54_ram[1361] = 252;
    exp_54_ram[1362] = 250;
    exp_54_ram[1363] = 250;
    exp_54_ram[1364] = 0;
    exp_54_ram[1365] = 250;
    exp_54_ram[1366] = 2;
    exp_54_ram[1367] = 0;
    exp_54_ram[1368] = 250;
    exp_54_ram[1369] = 0;
    exp_54_ram[1370] = 250;
    exp_54_ram[1371] = 3;
    exp_54_ram[1372] = 250;
    exp_54_ram[1373] = 0;
    exp_54_ram[1374] = 253;
    exp_54_ram[1375] = 0;
    exp_54_ram[1376] = 252;
    exp_54_ram[1377] = 250;
    exp_54_ram[1378] = 250;
    exp_54_ram[1379] = 0;
    exp_54_ram[1380] = 250;
    exp_54_ram[1381] = 0;
    exp_54_ram[1382] = 250;
    exp_54_ram[1383] = 0;
    exp_54_ram[1384] = 250;
    exp_54_ram[1385] = 0;
    exp_54_ram[1386] = 250;
    exp_54_ram[1387] = 0;
    exp_54_ram[1388] = 222;
    exp_54_ram[1389] = 253;
    exp_54_ram[1390] = 250;
    exp_54_ram[1391] = 0;
    exp_54_ram[1392] = 250;
    exp_54_ram[1393] = 255;
    exp_54_ram[1394] = 0;
    exp_54_ram[1395] = 253;
    exp_54_ram[1396] = 250;
    exp_54_ram[1397] = 250;
    exp_54_ram[1398] = 0;
    exp_54_ram[1399] = 250;
    exp_54_ram[1400] = 0;
    exp_54_ram[1401] = 0;
    exp_54_ram[1402] = 253;
    exp_54_ram[1403] = 0;
    exp_54_ram[1404] = 7;
    exp_54_ram[1405] = 7;
    exp_54_ram[1406] = 8;
    exp_54_ram[1407] = 0;
    exp_54_ram[1408] = 251;
    exp_54_ram[1409] = 2;
    exp_54_ram[1410] = 2;
    exp_54_ram[1411] = 3;
    exp_54_ram[1412] = 252;
    exp_54_ram[1413] = 0;
    exp_54_ram[1414] = 0;
    exp_54_ram[1415] = 0;
    exp_54_ram[1416] = 0;
    exp_54_ram[1417] = 0;
    exp_54_ram[1418] = 1;
    exp_54_ram[1419] = 1;
    exp_54_ram[1420] = 2;
    exp_54_ram[1421] = 252;
    exp_54_ram[1422] = 253;
    exp_54_ram[1423] = 254;
    exp_54_ram[1424] = 254;
    exp_54_ram[1425] = 254;
    exp_54_ram[1426] = 254;
    exp_54_ram[1427] = 253;
    exp_54_ram[1428] = 255;
    exp_54_ram[1429] = 0;
    exp_54_ram[1430] = 69;
    exp_54_ram[1431] = 208;
    exp_54_ram[1432] = 254;
    exp_54_ram[1433] = 254;
    exp_54_ram[1434] = 0;
    exp_54_ram[1435] = 2;
    exp_54_ram[1436] = 2;
    exp_54_ram[1437] = 5;
    exp_54_ram[1438] = 0;
    exp_54_ram[1439] = 254;
    exp_54_ram[1440] = 0;
    exp_54_ram[1441] = 0;
    exp_54_ram[1442] = 2;
    exp_54_ram[1443] = 0;
    exp_54_ram[1444] = 254;
    exp_54_ram[1445] = 254;
    exp_54_ram[1446] = 0;
    exp_54_ram[1447] = 219;
    exp_54_ram[1448] = 0;
    exp_54_ram[1449] = 0;
    exp_54_ram[1450] = 209;
    exp_54_ram[1451] = 0;
    exp_54_ram[1452] = 1;
    exp_54_ram[1453] = 1;
    exp_54_ram[1454] = 2;
    exp_54_ram[1455] = 0;
    exp_54_ram[1456] = 255;
    exp_54_ram[1457] = 0;
    exp_54_ram[1458] = 0;
    exp_54_ram[1459] = 1;
    exp_54_ram[1460] = 45;
    exp_54_ram[1461] = 209;
    exp_54_ram[1462] = 50;
    exp_54_ram[1463] = 50;
    exp_54_ram[1464] = 0;
    exp_54_ram[1465] = 0;
    exp_54_ram[1466] = 46;
    exp_54_ram[1467] = 241;
    exp_54_ram[1468] = 50;
    exp_54_ram[1469] = 50;
    exp_54_ram[1470] = 0;
    exp_54_ram[1471] = 0;
    exp_54_ram[1472] = 46;
    exp_54_ram[1473] = 239;
    exp_54_ram[1474] = 51;
    exp_54_ram[1475] = 51;
    exp_54_ram[1476] = 0;
    exp_54_ram[1477] = 0;
    exp_54_ram[1478] = 46;
    exp_54_ram[1479] = 238;
    exp_54_ram[1480] = 51;
    exp_54_ram[1481] = 51;
    exp_54_ram[1482] = 0;
    exp_54_ram[1483] = 0;
    exp_54_ram[1484] = 46;
    exp_54_ram[1485] = 236;
    exp_54_ram[1486] = 52;
    exp_54_ram[1487] = 52;
    exp_54_ram[1488] = 0;
    exp_54_ram[1489] = 0;
    exp_54_ram[1490] = 46;
    exp_54_ram[1491] = 235;
    exp_54_ram[1492] = 52;
    exp_54_ram[1493] = 52;
    exp_54_ram[1494] = 0;
    exp_54_ram[1495] = 0;
    exp_54_ram[1496] = 46;
    exp_54_ram[1497] = 233;
    exp_54_ram[1498] = 0;
    exp_54_ram[1499] = 0;
    exp_54_ram[1500] = 46;
    exp_54_ram[1501] = 232;
    exp_54_ram[1502] = 53;
    exp_54_ram[1503] = 53;
    exp_54_ram[1504] = 0;
    exp_54_ram[1505] = 0;
    exp_54_ram[1506] = 46;
    exp_54_ram[1507] = 231;
    exp_54_ram[1508] = 53;
    exp_54_ram[1509] = 53;
    exp_54_ram[1510] = 0;
    exp_54_ram[1511] = 0;
    exp_54_ram[1512] = 46;
    exp_54_ram[1513] = 229;
    exp_54_ram[1514] = 54;
    exp_54_ram[1515] = 54;
    exp_54_ram[1516] = 0;
    exp_54_ram[1517] = 0;
    exp_54_ram[1518] = 46;
    exp_54_ram[1519] = 228;
    exp_54_ram[1520] = 54;
    exp_54_ram[1521] = 54;
    exp_54_ram[1522] = 0;
    exp_54_ram[1523] = 0;
    exp_54_ram[1524] = 46;
    exp_54_ram[1525] = 226;
    exp_54_ram[1526] = 55;
    exp_54_ram[1527] = 55;
    exp_54_ram[1528] = 0;
    exp_54_ram[1529] = 0;
    exp_54_ram[1530] = 46;
    exp_54_ram[1531] = 225;
    exp_54_ram[1532] = 55;
    exp_54_ram[1533] = 55;
    exp_54_ram[1534] = 0;
    exp_54_ram[1535] = 0;
    exp_54_ram[1536] = 46;
    exp_54_ram[1537] = 223;
    exp_54_ram[1538] = 50;
    exp_54_ram[1539] = 50;
    exp_54_ram[1540] = 0;
    exp_54_ram[1541] = 0;
    exp_54_ram[1542] = 47;
    exp_54_ram[1543] = 222;
    exp_54_ram[1544] = 50;
    exp_54_ram[1545] = 50;
    exp_54_ram[1546] = 0;
    exp_54_ram[1547] = 0;
    exp_54_ram[1548] = 47;
    exp_54_ram[1549] = 220;
    exp_54_ram[1550] = 51;
    exp_54_ram[1551] = 51;
    exp_54_ram[1552] = 0;
    exp_54_ram[1553] = 0;
    exp_54_ram[1554] = 47;
    exp_54_ram[1555] = 219;
    exp_54_ram[1556] = 51;
    exp_54_ram[1557] = 51;
    exp_54_ram[1558] = 0;
    exp_54_ram[1559] = 0;
    exp_54_ram[1560] = 47;
    exp_54_ram[1561] = 217;
    exp_54_ram[1562] = 52;
    exp_54_ram[1563] = 52;
    exp_54_ram[1564] = 0;
    exp_54_ram[1565] = 0;
    exp_54_ram[1566] = 47;
    exp_54_ram[1567] = 216;
    exp_54_ram[1568] = 52;
    exp_54_ram[1569] = 52;
    exp_54_ram[1570] = 0;
    exp_54_ram[1571] = 0;
    exp_54_ram[1572] = 47;
    exp_54_ram[1573] = 214;
    exp_54_ram[1574] = 0;
    exp_54_ram[1575] = 0;
    exp_54_ram[1576] = 47;
    exp_54_ram[1577] = 213;
    exp_54_ram[1578] = 53;
    exp_54_ram[1579] = 53;
    exp_54_ram[1580] = 0;
    exp_54_ram[1581] = 0;
    exp_54_ram[1582] = 47;
    exp_54_ram[1583] = 212;
    exp_54_ram[1584] = 53;
    exp_54_ram[1585] = 53;
    exp_54_ram[1586] = 0;
    exp_54_ram[1587] = 0;
    exp_54_ram[1588] = 47;
    exp_54_ram[1589] = 210;
    exp_54_ram[1590] = 54;
    exp_54_ram[1591] = 54;
    exp_54_ram[1592] = 0;
    exp_54_ram[1593] = 0;
    exp_54_ram[1594] = 47;
    exp_54_ram[1595] = 209;
    exp_54_ram[1596] = 54;
    exp_54_ram[1597] = 54;
    exp_54_ram[1598] = 0;
    exp_54_ram[1599] = 0;
    exp_54_ram[1600] = 47;
    exp_54_ram[1601] = 207;
    exp_54_ram[1602] = 55;
    exp_54_ram[1603] = 55;
    exp_54_ram[1604] = 0;
    exp_54_ram[1605] = 0;
    exp_54_ram[1606] = 47;
    exp_54_ram[1607] = 206;
    exp_54_ram[1608] = 55;
    exp_54_ram[1609] = 55;
    exp_54_ram[1610] = 0;
    exp_54_ram[1611] = 0;
    exp_54_ram[1612] = 47;
    exp_54_ram[1613] = 204;
    exp_54_ram[1614] = 50;
    exp_54_ram[1615] = 50;
    exp_54_ram[1616] = 0;
    exp_54_ram[1617] = 0;
    exp_54_ram[1618] = 47;
    exp_54_ram[1619] = 203;
    exp_54_ram[1620] = 50;
    exp_54_ram[1621] = 50;
    exp_54_ram[1622] = 0;
    exp_54_ram[1623] = 0;
    exp_54_ram[1624] = 47;
    exp_54_ram[1625] = 201;
    exp_54_ram[1626] = 51;
    exp_54_ram[1627] = 51;
    exp_54_ram[1628] = 0;
    exp_54_ram[1629] = 0;
    exp_54_ram[1630] = 47;
    exp_54_ram[1631] = 200;
    exp_54_ram[1632] = 51;
    exp_54_ram[1633] = 51;
    exp_54_ram[1634] = 0;
    exp_54_ram[1635] = 0;
    exp_54_ram[1636] = 47;
    exp_54_ram[1637] = 198;
    exp_54_ram[1638] = 52;
    exp_54_ram[1639] = 52;
    exp_54_ram[1640] = 0;
    exp_54_ram[1641] = 0;
    exp_54_ram[1642] = 47;
    exp_54_ram[1643] = 197;
    exp_54_ram[1644] = 52;
    exp_54_ram[1645] = 52;
    exp_54_ram[1646] = 0;
    exp_54_ram[1647] = 0;
    exp_54_ram[1648] = 47;
    exp_54_ram[1649] = 195;
    exp_54_ram[1650] = 0;
    exp_54_ram[1651] = 0;
    exp_54_ram[1652] = 47;
    exp_54_ram[1653] = 194;
    exp_54_ram[1654] = 53;
    exp_54_ram[1655] = 53;
    exp_54_ram[1656] = 0;
    exp_54_ram[1657] = 0;
    exp_54_ram[1658] = 47;
    exp_54_ram[1659] = 193;
    exp_54_ram[1660] = 53;
    exp_54_ram[1661] = 53;
    exp_54_ram[1662] = 0;
    exp_54_ram[1663] = 0;
    exp_54_ram[1664] = 47;
    exp_54_ram[1665] = 191;
    exp_54_ram[1666] = 54;
    exp_54_ram[1667] = 54;
    exp_54_ram[1668] = 0;
    exp_54_ram[1669] = 0;
    exp_54_ram[1670] = 47;
    exp_54_ram[1671] = 190;
    exp_54_ram[1672] = 54;
    exp_54_ram[1673] = 54;
    exp_54_ram[1674] = 0;
    exp_54_ram[1675] = 0;
    exp_54_ram[1676] = 47;
    exp_54_ram[1677] = 188;
    exp_54_ram[1678] = 55;
    exp_54_ram[1679] = 55;
    exp_54_ram[1680] = 0;
    exp_54_ram[1681] = 0;
    exp_54_ram[1682] = 47;
    exp_54_ram[1683] = 187;
    exp_54_ram[1684] = 55;
    exp_54_ram[1685] = 55;
    exp_54_ram[1686] = 0;
    exp_54_ram[1687] = 0;
    exp_54_ram[1688] = 47;
    exp_54_ram[1689] = 185;
    exp_54_ram[1690] = 50;
    exp_54_ram[1691] = 50;
    exp_54_ram[1692] = 0;
    exp_54_ram[1693] = 0;
    exp_54_ram[1694] = 48;
    exp_54_ram[1695] = 184;
    exp_54_ram[1696] = 50;
    exp_54_ram[1697] = 50;
    exp_54_ram[1698] = 0;
    exp_54_ram[1699] = 0;
    exp_54_ram[1700] = 48;
    exp_54_ram[1701] = 182;
    exp_54_ram[1702] = 51;
    exp_54_ram[1703] = 51;
    exp_54_ram[1704] = 0;
    exp_54_ram[1705] = 0;
    exp_54_ram[1706] = 48;
    exp_54_ram[1707] = 181;
    exp_54_ram[1708] = 51;
    exp_54_ram[1709] = 51;
    exp_54_ram[1710] = 0;
    exp_54_ram[1711] = 0;
    exp_54_ram[1712] = 48;
    exp_54_ram[1713] = 179;
    exp_54_ram[1714] = 52;
    exp_54_ram[1715] = 52;
    exp_54_ram[1716] = 0;
    exp_54_ram[1717] = 0;
    exp_54_ram[1718] = 48;
    exp_54_ram[1719] = 178;
    exp_54_ram[1720] = 52;
    exp_54_ram[1721] = 52;
    exp_54_ram[1722] = 0;
    exp_54_ram[1723] = 0;
    exp_54_ram[1724] = 48;
    exp_54_ram[1725] = 176;
    exp_54_ram[1726] = 0;
    exp_54_ram[1727] = 0;
    exp_54_ram[1728] = 48;
    exp_54_ram[1729] = 175;
    exp_54_ram[1730] = 53;
    exp_54_ram[1731] = 53;
    exp_54_ram[1732] = 0;
    exp_54_ram[1733] = 0;
    exp_54_ram[1734] = 48;
    exp_54_ram[1735] = 174;
    exp_54_ram[1736] = 53;
    exp_54_ram[1737] = 53;
    exp_54_ram[1738] = 0;
    exp_54_ram[1739] = 0;
    exp_54_ram[1740] = 48;
    exp_54_ram[1741] = 172;
    exp_54_ram[1742] = 54;
    exp_54_ram[1743] = 54;
    exp_54_ram[1744] = 0;
    exp_54_ram[1745] = 0;
    exp_54_ram[1746] = 48;
    exp_54_ram[1747] = 171;
    exp_54_ram[1748] = 54;
    exp_54_ram[1749] = 54;
    exp_54_ram[1750] = 0;
    exp_54_ram[1751] = 0;
    exp_54_ram[1752] = 48;
    exp_54_ram[1753] = 169;
    exp_54_ram[1754] = 55;
    exp_54_ram[1755] = 55;
    exp_54_ram[1756] = 0;
    exp_54_ram[1757] = 0;
    exp_54_ram[1758] = 48;
    exp_54_ram[1759] = 168;
    exp_54_ram[1760] = 55;
    exp_54_ram[1761] = 55;
    exp_54_ram[1762] = 0;
    exp_54_ram[1763] = 0;
    exp_54_ram[1764] = 48;
    exp_54_ram[1765] = 166;
    exp_54_ram[1766] = 56;
    exp_54_ram[1767] = 56;
    exp_54_ram[1768] = 0;
    exp_54_ram[1769] = 0;
    exp_54_ram[1770] = 48;
    exp_54_ram[1771] = 165;
    exp_54_ram[1772] = 56;
    exp_54_ram[1773] = 56;
    exp_54_ram[1774] = 0;
    exp_54_ram[1775] = 0;
    exp_54_ram[1776] = 48;
    exp_54_ram[1777] = 163;
    exp_54_ram[1778] = 57;
    exp_54_ram[1779] = 57;
    exp_54_ram[1780] = 0;
    exp_54_ram[1781] = 0;
    exp_54_ram[1782] = 48;
    exp_54_ram[1783] = 162;
    exp_54_ram[1784] = 57;
    exp_54_ram[1785] = 57;
    exp_54_ram[1786] = 0;
    exp_54_ram[1787] = 0;
    exp_54_ram[1788] = 48;
    exp_54_ram[1789] = 160;
    exp_54_ram[1790] = 58;
    exp_54_ram[1791] = 58;
    exp_54_ram[1792] = 0;
    exp_54_ram[1793] = 0;
    exp_54_ram[1794] = 47;
    exp_54_ram[1795] = 159;
    exp_54_ram[1796] = 58;
    exp_54_ram[1797] = 58;
    exp_54_ram[1798] = 0;
    exp_54_ram[1799] = 0;
    exp_54_ram[1800] = 49;
    exp_54_ram[1801] = 157;
    exp_54_ram[1802] = 58;
    exp_54_ram[1803] = 58;
    exp_54_ram[1804] = 0;
    exp_54_ram[1805] = 0;
    exp_54_ram[1806] = 49;
    exp_54_ram[1807] = 156;
    exp_54_ram[1808] = 58;
    exp_54_ram[1809] = 58;
    exp_54_ram[1810] = 0;
    exp_54_ram[1811] = 0;
    exp_54_ram[1812] = 49;
    exp_54_ram[1813] = 154;
    exp_54_ram[1814] = 58;
    exp_54_ram[1815] = 58;
    exp_54_ram[1816] = 0;
    exp_54_ram[1817] = 0;
    exp_54_ram[1818] = 47;
    exp_54_ram[1819] = 153;
    exp_54_ram[1820] = 58;
    exp_54_ram[1821] = 58;
    exp_54_ram[1822] = 0;
    exp_54_ram[1823] = 0;
    exp_54_ram[1824] = 49;
    exp_54_ram[1825] = 151;
    exp_54_ram[1826] = 58;
    exp_54_ram[1827] = 58;
    exp_54_ram[1828] = 0;
    exp_54_ram[1829] = 0;
    exp_54_ram[1830] = 49;
    exp_54_ram[1831] = 150;
    exp_54_ram[1832] = 58;
    exp_54_ram[1833] = 58;
    exp_54_ram[1834] = 0;
    exp_54_ram[1835] = 0;
    exp_54_ram[1836] = 49;
    exp_54_ram[1837] = 148;
    exp_54_ram[1838] = 59;
    exp_54_ram[1839] = 59;
    exp_54_ram[1840] = 0;
    exp_54_ram[1841] = 0;
    exp_54_ram[1842] = 47;
    exp_54_ram[1843] = 147;
    exp_54_ram[1844] = 59;
    exp_54_ram[1845] = 59;
    exp_54_ram[1846] = 0;
    exp_54_ram[1847] = 0;
    exp_54_ram[1848] = 49;
    exp_54_ram[1849] = 145;
    exp_54_ram[1850] = 59;
    exp_54_ram[1851] = 59;
    exp_54_ram[1852] = 0;
    exp_54_ram[1853] = 0;
    exp_54_ram[1854] = 49;
    exp_54_ram[1855] = 144;
    exp_54_ram[1856] = 59;
    exp_54_ram[1857] = 59;
    exp_54_ram[1858] = 0;
    exp_54_ram[1859] = 0;
    exp_54_ram[1860] = 49;
    exp_54_ram[1861] = 142;
    exp_54_ram[1862] = 59;
    exp_54_ram[1863] = 59;
    exp_54_ram[1864] = 0;
    exp_54_ram[1865] = 0;
    exp_54_ram[1866] = 47;
    exp_54_ram[1867] = 141;
    exp_54_ram[1868] = 59;
    exp_54_ram[1869] = 59;
    exp_54_ram[1870] = 0;
    exp_54_ram[1871] = 0;
    exp_54_ram[1872] = 49;
    exp_54_ram[1873] = 139;
    exp_54_ram[1874] = 59;
    exp_54_ram[1875] = 59;
    exp_54_ram[1876] = 0;
    exp_54_ram[1877] = 0;
    exp_54_ram[1878] = 49;
    exp_54_ram[1879] = 138;
    exp_54_ram[1880] = 59;
    exp_54_ram[1881] = 59;
    exp_54_ram[1882] = 0;
    exp_54_ram[1883] = 0;
    exp_54_ram[1884] = 49;
    exp_54_ram[1885] = 136;
    exp_54_ram[1886] = 12;
    exp_54_ram[1887] = 231;
    exp_54_ram[1888] = 0;
    exp_54_ram[1889] = 0;
    exp_54_ram[1890] = 0;
    exp_54_ram[1891] = 1;
    exp_54_ram[1892] = 0;
    exp_54_ram[1893] = 255;
    exp_54_ram[1894] = 0;
    exp_54_ram[1895] = 0;
    exp_54_ram[1896] = 1;
    exp_54_ram[1897] = 145;
    exp_54_ram[1898] = 0;
    exp_54_ram[1899] = 0;
    exp_54_ram[1900] = 0;
    exp_54_ram[1901] = 1;
    exp_54_ram[1902] = 0;
    exp_54_ram[1903] = 128;
    exp_54_ram[1904] = 0;
    exp_54_ram[1905] = 0;
    exp_54_ram[1906] = 0;
    exp_54_ram[1907] = 0;
    exp_54_ram[1908] = 0;
    exp_54_ram[1909] = 0;
    exp_54_ram[1910] = 0;
    exp_54_ram[1911] = 0;
    exp_54_ram[1912] = 0;
    exp_54_ram[1913] = 0;
    exp_54_ram[1914] = 0;
    exp_54_ram[1915] = 0;
    exp_54_ram[1916] = 0;
    exp_54_ram[1917] = 0;
    exp_54_ram[1918] = 0;
    exp_54_ram[1919] = 0;
    exp_54_ram[1920] = 0;
    exp_54_ram[1921] = 0;
    exp_54_ram[1922] = 0;
    exp_54_ram[1923] = 0;
    exp_54_ram[1924] = 0;
    exp_54_ram[1925] = 0;
    exp_54_ram[1926] = 0;
    exp_54_ram[1927] = 0;
    exp_54_ram[1928] = 0;
    exp_54_ram[1929] = 0;
    exp_54_ram[1930] = 0;
    exp_54_ram[1931] = 0;
    exp_54_ram[1932] = 0;
    exp_54_ram[1933] = 0;
    exp_54_ram[1934] = 0;
    exp_54_ram[1935] = 0;
    exp_54_ram[1936] = 0;
    exp_54_ram[1937] = 0;
    exp_54_ram[1938] = 0;
    exp_54_ram[1939] = 0;
    exp_54_ram[1940] = 0;
    exp_54_ram[1941] = 0;
    exp_54_ram[1942] = 0;
    exp_54_ram[1943] = 0;
    exp_54_ram[1944] = 0;
    exp_54_ram[1945] = 0;
    exp_54_ram[1946] = 0;
    exp_54_ram[1947] = 0;
    exp_54_ram[1948] = 0;
    exp_54_ram[1949] = 0;
    exp_54_ram[1950] = 0;
    exp_54_ram[1951] = 0;
    exp_54_ram[1952] = 0;
    exp_54_ram[1953] = 0;
    exp_54_ram[1954] = 0;
    exp_54_ram[1955] = 0;
    exp_54_ram[1956] = 0;
    exp_54_ram[1957] = 0;
    exp_54_ram[1958] = 0;
    exp_54_ram[1959] = 0;
    exp_54_ram[1960] = 0;
    exp_54_ram[1961] = 0;
    exp_54_ram[1962] = 0;
    exp_54_ram[1963] = 0;
    exp_54_ram[1964] = 0;
    exp_54_ram[1965] = 0;
    exp_54_ram[1966] = 0;
    exp_54_ram[1967] = 0;
    exp_54_ram[1968] = 0;
    exp_54_ram[1969] = 0;
    exp_54_ram[1970] = 0;
    exp_54_ram[1971] = 0;
    exp_54_ram[1972] = 0;
    exp_54_ram[1973] = 0;
    exp_54_ram[1974] = 0;
    exp_54_ram[1975] = 0;
    exp_54_ram[1976] = 0;
    exp_54_ram[1977] = 0;
    exp_54_ram[1978] = 0;
    exp_54_ram[1979] = 0;
    exp_54_ram[1980] = 0;
    exp_54_ram[1981] = 0;
    exp_54_ram[1982] = 0;
    exp_54_ram[1983] = 0;
    exp_54_ram[1984] = 0;
    exp_54_ram[1985] = 0;
    exp_54_ram[1986] = 0;
    exp_54_ram[1987] = 0;
    exp_54_ram[1988] = 0;
    exp_54_ram[1989] = 0;
    exp_54_ram[1990] = 0;
    exp_54_ram[1991] = 0;
    exp_54_ram[1992] = 0;
    exp_54_ram[1993] = 0;
    exp_54_ram[1994] = 0;
    exp_54_ram[1995] = 0;
    exp_54_ram[1996] = 0;
    exp_54_ram[1997] = 0;
    exp_54_ram[1998] = 0;
    exp_54_ram[1999] = 0;
    exp_54_ram[2000] = 0;
    exp_54_ram[2001] = 0;
    exp_54_ram[2002] = 0;
    exp_54_ram[2003] = 0;
    exp_54_ram[2004] = 0;
    exp_54_ram[2005] = 0;
    exp_54_ram[2006] = 0;
    exp_54_ram[2007] = 0;
    exp_54_ram[2008] = 0;
    exp_54_ram[2009] = 0;
    exp_54_ram[2010] = 0;
    exp_54_ram[2011] = 0;
    exp_54_ram[2012] = 0;
    exp_54_ram[2013] = 0;
    exp_54_ram[2014] = 0;
    exp_54_ram[2015] = 0;
    exp_54_ram[2016] = 0;
    exp_54_ram[2017] = 0;
    exp_54_ram[2018] = 0;
    exp_54_ram[2019] = 0;
    exp_54_ram[2020] = 0;
    exp_54_ram[2021] = 0;
    exp_54_ram[2022] = 0;
    exp_54_ram[2023] = 0;
    exp_54_ram[2024] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_252;
  assign exp_252 = exp_533;

  reg [3:0] exp_533_reg;
  always@(*) begin
    case (exp_385)
      0:exp_533_reg <= exp_520;
      1:exp_533_reg <= exp_525;
      2:exp_533_reg <= exp_526;
      3:exp_533_reg <= exp_527;
      4:exp_533_reg <= exp_528;
      5:exp_533_reg <= exp_529;
      6:exp_533_reg <= exp_530;
      7:exp_533_reg <= exp_531;
      default:exp_533_reg <= exp_532;
    endcase
  end
  assign exp_533 = exp_533_reg;
  assign exp_532 = 0;
  assign exp_520 = exp_516 << exp_519;
  assign exp_516 = 1;
  assign exp_519 = exp_518 + exp_517;
  assign exp_518 = 0;
  assign exp_517 = exp_453[1:0];
  assign exp_525 = exp_521 << exp_524;
  assign exp_521 = 3;
  assign exp_524 = exp_523 + exp_522;
  assign exp_523 = 0;
  assign exp_522 = exp_453[1:1];
  assign exp_526 = 15;
  assign exp_527 = 0;
  assign exp_528 = 0;
  assign exp_529 = 0;
  assign exp_530 = 0;
  assign exp_531 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_247;
  assign exp_247 = exp_515;

  reg [31:0] exp_515_reg;
  always@(*) begin
    case (exp_385)
      0:exp_515_reg <= exp_502;
      1:exp_515_reg <= exp_506;
      2:exp_515_reg <= exp_508;
      3:exp_515_reg <= exp_509;
      4:exp_515_reg <= exp_510;
      5:exp_515_reg <= exp_511;
      6:exp_515_reg <= exp_512;
      7:exp_515_reg <= exp_513;
      default:exp_515_reg <= exp_514;
    endcase
  end
  assign exp_515 = exp_515_reg;
  assign exp_514 = 0;

  reg [31:0] exp_502_reg;
  always@(*) begin
    case (exp_456)
      0:exp_502_reg <= exp_488;
      1:exp_502_reg <= exp_496;
      2:exp_502_reg <= exp_498;
      3:exp_502_reg <= exp_500;
      default:exp_502_reg <= exp_501;
    endcase
  end
  assign exp_502 = exp_502_reg;
  assign exp_501 = 0;
  assign exp_488 = exp_487;
  assign exp_487 = exp_486 + exp_485;
  assign exp_486 = 0;
  assign exp_485 = exp_375[7:0];

      reg [31:0] exp_375_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_375_reg <= exp_318;
        end
      end
      assign exp_375 = exp_375_reg;
      assign exp_496 = exp_488 << exp_495;
  assign exp_495 = 8;
  assign exp_498 = exp_488 << exp_497;
  assign exp_497 = 16;
  assign exp_500 = exp_488 << exp_499;
  assign exp_499 = 24;

  reg [31:0] exp_506_reg;
  always@(*) begin
    case (exp_459)
      0:exp_506_reg <= exp_492;
      1:exp_506_reg <= exp_504;
      default:exp_506_reg <= exp_505;
    endcase
  end
  assign exp_506 = exp_506_reg;
  assign exp_459 = exp_458 + exp_457;
  assign exp_458 = 0;
  assign exp_457 = exp_453[1:1];
  assign exp_505 = 0;
  assign exp_492 = exp_491;
  assign exp_491 = exp_490 + exp_489;
  assign exp_490 = 0;
  assign exp_489 = exp_375[15:0];
  assign exp_504 = exp_492 << exp_503;
  assign exp_503 = 16;
  assign exp_508 = exp_507 + exp_494;
  assign exp_507 = 0;
  assign exp_494 = exp_493 + exp_375;
  assign exp_493 = 0;
  assign exp_509 = 0;
  assign exp_510 = 0;
  assign exp_511 = 0;
  assign exp_512 = 0;
  assign exp_513 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 0;
    exp_47_ram[32] = 1;
    exp_47_ram[33] = 16;
    exp_47_ram[34] = 0;
    exp_47_ram[35] = 0;
    exp_47_ram[36] = 114;
    exp_47_ram[37] = 46;
    exp_47_ram[38] = 0;
    exp_47_ram[39] = 111;
    exp_47_ram[40] = 108;
    exp_47_ram[41] = 0;
    exp_47_ram[42] = 102;
    exp_47_ram[43] = 0;
    exp_47_ram[44] = 102;
    exp_47_ram[45] = 0;
    exp_47_ram[46] = 0;
    exp_47_ram[47] = 102;
    exp_47_ram[48] = 0;
    exp_47_ram[49] = 102;
    exp_47_ram[50] = 0;
    exp_47_ram[51] = 115;
    exp_47_ram[52] = 0;
    exp_47_ram[53] = 114;
    exp_47_ram[54] = 116;
    exp_47_ram[55] = 0;
    exp_47_ram[56] = 111;
    exp_47_ram[57] = 0;
    exp_47_ram[58] = 109;
    exp_47_ram[59] = 46;
    exp_47_ram[60] = 0;
    exp_47_ram[61] = 114;
    exp_47_ram[62] = 46;
    exp_47_ram[63] = 0;
    exp_47_ram[64] = 114;
    exp_47_ram[65] = 112;
    exp_47_ram[66] = 0;
    exp_47_ram[67] = 109;
    exp_47_ram[68] = 46;
    exp_47_ram[69] = 0;
    exp_47_ram[70] = 102;
    exp_47_ram[71] = 0;
    exp_47_ram[72] = 114;
    exp_47_ram[73] = 46;
    exp_47_ram[74] = 0;
    exp_47_ram[75] = 102;
    exp_47_ram[76] = 0;
    exp_47_ram[77] = 114;
    exp_47_ram[78] = 110;
    exp_47_ram[79] = 0;
    exp_47_ram[80] = 100;
    exp_47_ram[81] = 0;
    exp_47_ram[82] = 100;
    exp_47_ram[83] = 100;
    exp_47_ram[84] = 0;
    exp_47_ram[85] = 100;
    exp_47_ram[86] = 100;
    exp_47_ram[87] = 0;
    exp_47_ram[88] = 100;
    exp_47_ram[89] = 102;
    exp_47_ram[90] = 0;
    exp_47_ram[91] = 100;
    exp_47_ram[92] = 103;
    exp_47_ram[93] = 0;
    exp_47_ram[94] = 114;
    exp_47_ram[95] = 107;
    exp_47_ram[96] = 0;
    exp_47_ram[97] = 100;
    exp_47_ram[98] = 100;
    exp_47_ram[99] = 0;
    exp_47_ram[100] = 115;
    exp_47_ram[101] = 100;
    exp_47_ram[102] = 106;
    exp_47_ram[103] = 106;
    exp_47_ram[104] = 115;
    exp_47_ram[105] = 0;
    exp_47_ram[106] = 100;
    exp_47_ram[107] = 100;
    exp_47_ram[108] = 0;
    exp_47_ram[109] = 114;
    exp_47_ram[110] = 114;
    exp_47_ram[111] = 0;
    exp_47_ram[112] = 114;
    exp_47_ram[113] = 46;
    exp_47_ram[114] = 0;
    exp_47_ram[115] = 51;
    exp_47_ram[116] = 49;
    exp_47_ram[117] = 52;
    exp_47_ram[118] = 97;
    exp_47_ram[119] = 50;
    exp_47_ram[120] = 100;
    exp_47_ram[121] = 115;
    exp_47_ram[122] = 51;
    exp_47_ram[123] = 49;
    exp_47_ram[124] = 97;
    exp_47_ram[125] = 103;
    exp_47_ram[126] = 0;
    exp_47_ram[127] = 114;
    exp_47_ram[128] = 46;
    exp_47_ram[129] = 0;
    exp_47_ram[130] = 51;
    exp_47_ram[131] = 0;
    exp_47_ram[132] = 52;
    exp_47_ram[133] = 0;
    exp_47_ram[134] = 109;
    exp_47_ram[135] = 46;
    exp_47_ram[136] = 0;
    exp_47_ram[137] = 51;
    exp_47_ram[138] = 0;
    exp_47_ram[139] = 51;
    exp_47_ram[140] = 0;
    exp_47_ram[141] = 99;
    exp_47_ram[142] = 0;
    exp_47_ram[143] = 100;
    exp_47_ram[144] = 0;
    exp_47_ram[145] = 114;
    exp_47_ram[146] = 46;
    exp_47_ram[147] = 0;
    exp_47_ram[148] = 109;
    exp_47_ram[149] = 46;
    exp_47_ram[150] = 117;
    exp_47_ram[151] = 112;
    exp_47_ram[152] = 32;
    exp_47_ram[153] = 50;
    exp_47_ram[154] = 48;
    exp_47_ram[155] = 50;
    exp_47_ram[156] = 0;
    exp_47_ram[157] = 117;
    exp_47_ram[158] = 112;
    exp_47_ram[159] = 32;
    exp_47_ram[160] = 50;
    exp_47_ram[161] = 48;
    exp_47_ram[162] = 50;
    exp_47_ram[163] = 0;
    exp_47_ram[164] = 102;
    exp_47_ram[165] = 0;
    exp_47_ram[166] = 102;
    exp_47_ram[167] = 0;
    exp_47_ram[168] = 102;
    exp_47_ram[169] = 0;
    exp_47_ram[170] = 117;
    exp_47_ram[171] = 112;
    exp_47_ram[172] = 32;
    exp_47_ram[173] = 50;
    exp_47_ram[174] = 48;
    exp_47_ram[175] = 50;
    exp_47_ram[176] = 0;
    exp_47_ram[177] = 32;
    exp_47_ram[178] = 108;
    exp_47_ram[179] = 32;
    exp_47_ram[180] = 108;
    exp_47_ram[181] = 32;
    exp_47_ram[182] = 108;
    exp_47_ram[183] = 115;
    exp_47_ram[184] = 114;
    exp_47_ram[185] = 102;
    exp_47_ram[186] = 46;
    exp_47_ram[187] = 10;
    exp_47_ram[188] = 48;
    exp_47_ram[189] = 102;
    exp_47_ram[190] = 0;
    exp_47_ram[191] = 10;
    exp_47_ram[192] = 100;
    exp_47_ram[193] = 50;
    exp_47_ram[194] = 50;
    exp_47_ram[195] = 103;
    exp_47_ram[196] = 0;
    exp_47_ram[197] = 10;
    exp_47_ram[198] = 10;
    exp_47_ram[199] = 10;
    exp_47_ram[200] = 181;
    exp_47_ram[201] = 176;
    exp_47_ram[202] = 227;
    exp_47_ram[203] = 228;
    exp_47_ram[204] = 28;
    exp_47_ram[205] = 26;
    exp_47_ram[206] = 241;
    exp_47_ram[207] = 80;
    exp_47_ram[208] = 174;
    exp_47_ram[209] = 132;
    exp_47_ram[210] = 153;
    exp_47_ram[211] = 185;
    exp_47_ram[212] = 0;
    exp_47_ram[213] = 240;
    exp_47_ram[214] = 0;
    exp_47_ram[215] = 36;
    exp_47_ram[216] = 0;
    exp_47_ram[217] = 89;
    exp_47_ram[218] = 0;
    exp_47_ram[219] = 143;
    exp_47_ram[220] = 0;
    exp_47_ram[221] = 195;
    exp_47_ram[222] = 0;
    exp_47_ram[223] = 248;
    exp_47_ram[224] = 0;
    exp_47_ram[225] = 46;
    exp_47_ram[226] = 0;
    exp_47_ram[227] = 99;
    exp_47_ram[228] = 0;
    exp_47_ram[229] = 151;
    exp_47_ram[230] = 0;
    exp_47_ram[231] = 205;
    exp_47_ram[232] = 0;
    exp_47_ram[233] = 248;
    exp_47_ram[234] = 0;
    exp_47_ram[235] = 248;
    exp_47_ram[236] = 0;
    exp_47_ram[237] = 240;
    exp_47_ram[238] = 0;
    exp_47_ram[239] = 240;
    exp_47_ram[240] = 165;
    exp_47_ram[241] = 0;
    exp_47_ram[242] = 5;
    exp_47_ram[243] = 0;
    exp_47_ram[244] = 167;
    exp_47_ram[245] = 7;
    exp_47_ram[246] = 7;
    exp_47_ram[247] = 0;
    exp_47_ram[248] = 21;
    exp_47_ram[249] = 229;
    exp_47_ram[250] = 159;
    exp_47_ram[251] = 1;
    exp_47_ram[252] = 0;
    exp_47_ram[253] = 129;
    exp_47_ram[254] = 199;
    exp_47_ram[255] = 17;
    exp_47_ram[256] = 4;
    exp_47_ram[257] = 95;
    exp_47_ram[258] = 160;
    exp_47_ram[259] = 193;
    exp_47_ram[260] = 244;
    exp_47_ram[261] = 129;
    exp_47_ram[262] = 0;
    exp_47_ram[263] = 1;
    exp_47_ram[264] = 0;
    exp_47_ram[265] = 1;
    exp_47_ram[266] = 129;
    exp_47_ram[267] = 1;
    exp_47_ram[268] = 5;
    exp_47_ram[269] = 180;
    exp_47_ram[270] = 196;
    exp_47_ram[271] = 212;
    exp_47_ram[272] = 244;
    exp_47_ram[273] = 0;
    exp_47_ram[274] = 193;
    exp_47_ram[275] = 1;
    exp_47_ram[276] = 0;
    exp_47_ram[277] = 1;
    exp_47_ram[278] = 17;
    exp_47_ram[279] = 129;
    exp_47_ram[280] = 1;
    exp_47_ram[281] = 5;
    exp_47_ram[282] = 180;
    exp_47_ram[283] = 196;
    exp_47_ram[284] = 212;
    exp_47_ram[285] = 244;
    exp_47_ram[286] = 244;
    exp_47_ram[287] = 7;
    exp_47_ram[288] = 244;
    exp_47_ram[289] = 7;
    exp_47_ram[290] = 64;
    exp_47_ram[291] = 0;
    exp_47_ram[292] = 193;
    exp_47_ram[293] = 129;
    exp_47_ram[294] = 1;
    exp_47_ram[295] = 0;
    exp_47_ram[296] = 1;
    exp_47_ram[297] = 129;
    exp_47_ram[298] = 1;
    exp_47_ram[299] = 164;
    exp_47_ram[300] = 180;
    exp_47_ram[301] = 196;
    exp_47_ram[302] = 244;
    exp_47_ram[303] = 0;
    exp_47_ram[304] = 196;
    exp_47_ram[305] = 23;
    exp_47_ram[306] = 244;
    exp_47_ram[307] = 196;
    exp_47_ram[308] = 7;
    exp_47_ram[309] = 7;
    exp_47_ram[310] = 132;
    exp_47_ram[311] = 247;
    exp_47_ram[312] = 228;
    exp_47_ram[313] = 7;
    exp_47_ram[314] = 196;
    exp_47_ram[315] = 196;
    exp_47_ram[316] = 247;
    exp_47_ram[317] = 7;
    exp_47_ram[318] = 193;
    exp_47_ram[319] = 1;
    exp_47_ram[320] = 0;
    exp_47_ram[321] = 1;
    exp_47_ram[322] = 129;
    exp_47_ram[323] = 1;
    exp_47_ram[324] = 5;
    exp_47_ram[325] = 244;
    exp_47_ram[326] = 244;
    exp_47_ram[327] = 240;
    exp_47_ram[328] = 231;
    exp_47_ram[329] = 244;
    exp_47_ram[330] = 144;
    exp_47_ram[331] = 231;
    exp_47_ram[332] = 16;
    exp_47_ram[333] = 128;
    exp_47_ram[334] = 0;
    exp_47_ram[335] = 23;
    exp_47_ram[336] = 247;
    exp_47_ram[337] = 7;
    exp_47_ram[338] = 193;
    exp_47_ram[339] = 1;
    exp_47_ram[340] = 0;
    exp_47_ram[341] = 1;
    exp_47_ram[342] = 17;
    exp_47_ram[343] = 129;
    exp_47_ram[344] = 1;
    exp_47_ram[345] = 164;
    exp_47_ram[346] = 4;
    exp_47_ram[347] = 0;
    exp_47_ram[348] = 196;
    exp_47_ram[349] = 7;
    exp_47_ram[350] = 39;
    exp_47_ram[351] = 231;
    exp_47_ram[352] = 23;
    exp_47_ram[353] = 7;
    exp_47_ram[354] = 196;
    exp_47_ram[355] = 7;
    exp_47_ram[356] = 23;
    exp_47_ram[357] = 196;
    exp_47_ram[358] = 215;
    exp_47_ram[359] = 7;
    exp_47_ram[360] = 246;
    exp_47_ram[361] = 7;
    exp_47_ram[362] = 244;
    exp_47_ram[363] = 196;
    exp_47_ram[364] = 7;
    exp_47_ram[365] = 7;
    exp_47_ram[366] = 7;
    exp_47_ram[367] = 159;
    exp_47_ram[368] = 5;
    exp_47_ram[369] = 7;
    exp_47_ram[370] = 196;
    exp_47_ram[371] = 7;
    exp_47_ram[372] = 193;
    exp_47_ram[373] = 129;
    exp_47_ram[374] = 1;
    exp_47_ram[375] = 0;
    exp_47_ram[376] = 1;
    exp_47_ram[377] = 17;
    exp_47_ram[378] = 129;
    exp_47_ram[379] = 1;
    exp_47_ram[380] = 164;
    exp_47_ram[381] = 180;
    exp_47_ram[382] = 196;
    exp_47_ram[383] = 212;
    exp_47_ram[384] = 228;
    exp_47_ram[385] = 244;
    exp_47_ram[386] = 4;
    exp_47_ram[387] = 20;
    exp_47_ram[388] = 68;
    exp_47_ram[389] = 244;
    exp_47_ram[390] = 4;
    exp_47_ram[391] = 39;
    exp_47_ram[392] = 7;
    exp_47_ram[393] = 4;
    exp_47_ram[394] = 23;
    exp_47_ram[395] = 7;
    exp_47_ram[396] = 132;
    exp_47_ram[397] = 244;
    exp_47_ram[398] = 64;
    exp_47_ram[399] = 68;
    exp_47_ram[400] = 23;
    exp_47_ram[401] = 228;
    exp_47_ram[402] = 196;
    exp_47_ram[403] = 4;
    exp_47_ram[404] = 7;
    exp_47_ram[405] = 132;
    exp_47_ram[406] = 0;
    exp_47_ram[407] = 7;
    exp_47_ram[408] = 196;
    exp_47_ram[409] = 23;
    exp_47_ram[410] = 244;
    exp_47_ram[411] = 196;
    exp_47_ram[412] = 68;
    exp_47_ram[413] = 247;
    exp_47_ram[414] = 0;
    exp_47_ram[415] = 132;
    exp_47_ram[416] = 247;
    exp_47_ram[417] = 244;
    exp_47_ram[418] = 196;
    exp_47_ram[419] = 132;
    exp_47_ram[420] = 247;
    exp_47_ram[421] = 7;
    exp_47_ram[422] = 68;
    exp_47_ram[423] = 23;
    exp_47_ram[424] = 228;
    exp_47_ram[425] = 196;
    exp_47_ram[426] = 4;
    exp_47_ram[427] = 7;
    exp_47_ram[428] = 132;
    exp_47_ram[429] = 7;
    exp_47_ram[430] = 132;
    exp_47_ram[431] = 7;
    exp_47_ram[432] = 4;
    exp_47_ram[433] = 39;
    exp_47_ram[434] = 7;
    exp_47_ram[435] = 128;
    exp_47_ram[436] = 68;
    exp_47_ram[437] = 23;
    exp_47_ram[438] = 228;
    exp_47_ram[439] = 196;
    exp_47_ram[440] = 4;
    exp_47_ram[441] = 7;
    exp_47_ram[442] = 132;
    exp_47_ram[443] = 0;
    exp_47_ram[444] = 7;
    exp_47_ram[445] = 68;
    exp_47_ram[446] = 132;
    exp_47_ram[447] = 247;
    exp_47_ram[448] = 68;
    exp_47_ram[449] = 231;
    exp_47_ram[450] = 68;
    exp_47_ram[451] = 7;
    exp_47_ram[452] = 193;
    exp_47_ram[453] = 129;
    exp_47_ram[454] = 1;
    exp_47_ram[455] = 0;
    exp_47_ram[456] = 1;
    exp_47_ram[457] = 17;
    exp_47_ram[458] = 129;
    exp_47_ram[459] = 1;
    exp_47_ram[460] = 164;
    exp_47_ram[461] = 180;
    exp_47_ram[462] = 196;
    exp_47_ram[463] = 212;
    exp_47_ram[464] = 228;
    exp_47_ram[465] = 244;
    exp_47_ram[466] = 8;
    exp_47_ram[467] = 20;
    exp_47_ram[468] = 244;
    exp_47_ram[469] = 132;
    exp_47_ram[470] = 39;
    exp_47_ram[471] = 7;
    exp_47_ram[472] = 68;
    exp_47_ram[473] = 7;
    exp_47_ram[474] = 132;
    exp_47_ram[475] = 23;
    exp_47_ram[476] = 7;
    exp_47_ram[477] = 116;
    exp_47_ram[478] = 7;
    exp_47_ram[479] = 132;
    exp_47_ram[480] = 199;
    exp_47_ram[481] = 7;
    exp_47_ram[482] = 68;
    exp_47_ram[483] = 247;
    exp_47_ram[484] = 244;
    exp_47_ram[485] = 0;
    exp_47_ram[486] = 132;
    exp_47_ram[487] = 23;
    exp_47_ram[488] = 228;
    exp_47_ram[489] = 196;
    exp_47_ram[490] = 247;
    exp_47_ram[491] = 0;
    exp_47_ram[492] = 231;
    exp_47_ram[493] = 132;
    exp_47_ram[494] = 4;
    exp_47_ram[495] = 247;
    exp_47_ram[496] = 132;
    exp_47_ram[497] = 240;
    exp_47_ram[498] = 231;
    exp_47_ram[499] = 0;
    exp_47_ram[500] = 132;
    exp_47_ram[501] = 23;
    exp_47_ram[502] = 228;
    exp_47_ram[503] = 196;
    exp_47_ram[504] = 247;
    exp_47_ram[505] = 0;
    exp_47_ram[506] = 231;
    exp_47_ram[507] = 132;
    exp_47_ram[508] = 23;
    exp_47_ram[509] = 7;
    exp_47_ram[510] = 132;
    exp_47_ram[511] = 68;
    exp_47_ram[512] = 247;
    exp_47_ram[513] = 132;
    exp_47_ram[514] = 240;
    exp_47_ram[515] = 231;
    exp_47_ram[516] = 132;
    exp_47_ram[517] = 7;
    exp_47_ram[518] = 7;
    exp_47_ram[519] = 132;
    exp_47_ram[520] = 7;
    exp_47_ram[521] = 7;
    exp_47_ram[522] = 132;
    exp_47_ram[523] = 7;
    exp_47_ram[524] = 132;
    exp_47_ram[525] = 4;
    exp_47_ram[526] = 247;
    exp_47_ram[527] = 132;
    exp_47_ram[528] = 68;
    exp_47_ram[529] = 247;
    exp_47_ram[530] = 132;
    exp_47_ram[531] = 247;
    exp_47_ram[532] = 244;
    exp_47_ram[533] = 132;
    exp_47_ram[534] = 7;
    exp_47_ram[535] = 4;
    exp_47_ram[536] = 0;
    exp_47_ram[537] = 247;
    exp_47_ram[538] = 132;
    exp_47_ram[539] = 247;
    exp_47_ram[540] = 244;
    exp_47_ram[541] = 4;
    exp_47_ram[542] = 0;
    exp_47_ram[543] = 247;
    exp_47_ram[544] = 132;
    exp_47_ram[545] = 7;
    exp_47_ram[546] = 7;
    exp_47_ram[547] = 132;
    exp_47_ram[548] = 240;
    exp_47_ram[549] = 231;
    exp_47_ram[550] = 132;
    exp_47_ram[551] = 23;
    exp_47_ram[552] = 228;
    exp_47_ram[553] = 196;
    exp_47_ram[554] = 247;
    exp_47_ram[555] = 128;
    exp_47_ram[556] = 231;
    exp_47_ram[557] = 192;
    exp_47_ram[558] = 4;
    exp_47_ram[559] = 0;
    exp_47_ram[560] = 247;
    exp_47_ram[561] = 132;
    exp_47_ram[562] = 7;
    exp_47_ram[563] = 7;
    exp_47_ram[564] = 132;
    exp_47_ram[565] = 240;
    exp_47_ram[566] = 231;
    exp_47_ram[567] = 132;
    exp_47_ram[568] = 23;
    exp_47_ram[569] = 228;
    exp_47_ram[570] = 196;
    exp_47_ram[571] = 247;
    exp_47_ram[572] = 128;
    exp_47_ram[573] = 231;
    exp_47_ram[574] = 128;
    exp_47_ram[575] = 4;
    exp_47_ram[576] = 32;
    exp_47_ram[577] = 247;
    exp_47_ram[578] = 132;
    exp_47_ram[579] = 240;
    exp_47_ram[580] = 231;
    exp_47_ram[581] = 132;
    exp_47_ram[582] = 23;
    exp_47_ram[583] = 228;
    exp_47_ram[584] = 196;
    exp_47_ram[585] = 247;
    exp_47_ram[586] = 32;
    exp_47_ram[587] = 231;
    exp_47_ram[588] = 132;
    exp_47_ram[589] = 240;
    exp_47_ram[590] = 231;
    exp_47_ram[591] = 132;
    exp_47_ram[592] = 23;
    exp_47_ram[593] = 228;
    exp_47_ram[594] = 196;
    exp_47_ram[595] = 247;
    exp_47_ram[596] = 0;
    exp_47_ram[597] = 231;
    exp_47_ram[598] = 132;
    exp_47_ram[599] = 240;
    exp_47_ram[600] = 231;
    exp_47_ram[601] = 116;
    exp_47_ram[602] = 7;
    exp_47_ram[603] = 132;
    exp_47_ram[604] = 23;
    exp_47_ram[605] = 228;
    exp_47_ram[606] = 196;
    exp_47_ram[607] = 247;
    exp_47_ram[608] = 208;
    exp_47_ram[609] = 231;
    exp_47_ram[610] = 128;
    exp_47_ram[611] = 132;
    exp_47_ram[612] = 71;
    exp_47_ram[613] = 7;
    exp_47_ram[614] = 132;
    exp_47_ram[615] = 23;
    exp_47_ram[616] = 228;
    exp_47_ram[617] = 196;
    exp_47_ram[618] = 247;
    exp_47_ram[619] = 176;
    exp_47_ram[620] = 231;
    exp_47_ram[621] = 192;
    exp_47_ram[622] = 132;
    exp_47_ram[623] = 135;
    exp_47_ram[624] = 7;
    exp_47_ram[625] = 132;
    exp_47_ram[626] = 23;
    exp_47_ram[627] = 228;
    exp_47_ram[628] = 196;
    exp_47_ram[629] = 247;
    exp_47_ram[630] = 0;
    exp_47_ram[631] = 231;
    exp_47_ram[632] = 132;
    exp_47_ram[633] = 68;
    exp_47_ram[634] = 132;
    exp_47_ram[635] = 196;
    exp_47_ram[636] = 4;
    exp_47_ram[637] = 68;
    exp_47_ram[638] = 132;
    exp_47_ram[639] = 196;
    exp_47_ram[640] = 31;
    exp_47_ram[641] = 5;
    exp_47_ram[642] = 7;
    exp_47_ram[643] = 193;
    exp_47_ram[644] = 129;
    exp_47_ram[645] = 1;
    exp_47_ram[646] = 0;
    exp_47_ram[647] = 1;
    exp_47_ram[648] = 17;
    exp_47_ram[649] = 129;
    exp_47_ram[650] = 1;
    exp_47_ram[651] = 164;
    exp_47_ram[652] = 180;
    exp_47_ram[653] = 196;
    exp_47_ram[654] = 212;
    exp_47_ram[655] = 228;
    exp_47_ram[656] = 4;
    exp_47_ram[657] = 20;
    exp_47_ram[658] = 244;
    exp_47_ram[659] = 4;
    exp_47_ram[660] = 196;
    exp_47_ram[661] = 7;
    exp_47_ram[662] = 68;
    exp_47_ram[663] = 247;
    exp_47_ram[664] = 244;
    exp_47_ram[665] = 68;
    exp_47_ram[666] = 7;
    exp_47_ram[667] = 7;
    exp_47_ram[668] = 196;
    exp_47_ram[669] = 7;
    exp_47_ram[670] = 196;
    exp_47_ram[671] = 68;
    exp_47_ram[672] = 247;
    exp_47_ram[673] = 244;
    exp_47_ram[674] = 180;
    exp_47_ram[675] = 144;
    exp_47_ram[676] = 231;
    exp_47_ram[677] = 180;
    exp_47_ram[678] = 7;
    exp_47_ram[679] = 247;
    exp_47_ram[680] = 0;
    exp_47_ram[681] = 68;
    exp_47_ram[682] = 7;
    exp_47_ram[683] = 7;
    exp_47_ram[684] = 16;
    exp_47_ram[685] = 128;
    exp_47_ram[686] = 16;
    exp_47_ram[687] = 180;
    exp_47_ram[688] = 231;
    exp_47_ram[689] = 247;
    exp_47_ram[690] = 103;
    exp_47_ram[691] = 247;
    exp_47_ram[692] = 196;
    exp_47_ram[693] = 23;
    exp_47_ram[694] = 212;
    exp_47_ram[695] = 4;
    exp_47_ram[696] = 230;
    exp_47_ram[697] = 247;
    exp_47_ram[698] = 196;
    exp_47_ram[699] = 68;
    exp_47_ram[700] = 247;
    exp_47_ram[701] = 244;
    exp_47_ram[702] = 196;
    exp_47_ram[703] = 7;
    exp_47_ram[704] = 196;
    exp_47_ram[705] = 240;
    exp_47_ram[706] = 231;
    exp_47_ram[707] = 180;
    exp_47_ram[708] = 132;
    exp_47_ram[709] = 68;
    exp_47_ram[710] = 241;
    exp_47_ram[711] = 4;
    exp_47_ram[712] = 241;
    exp_47_ram[713] = 4;
    exp_47_ram[714] = 241;
    exp_47_ram[715] = 68;
    exp_47_ram[716] = 6;
    exp_47_ram[717] = 196;
    exp_47_ram[718] = 4;
    exp_47_ram[719] = 68;
    exp_47_ram[720] = 132;
    exp_47_ram[721] = 196;
    exp_47_ram[722] = 159;
    exp_47_ram[723] = 5;
    exp_47_ram[724] = 7;
    exp_47_ram[725] = 193;
    exp_47_ram[726] = 129;
    exp_47_ram[727] = 1;
    exp_47_ram[728] = 0;
    exp_47_ram[729] = 1;
    exp_47_ram[730] = 17;
    exp_47_ram[731] = 129;
    exp_47_ram[732] = 1;
    exp_47_ram[733] = 164;
    exp_47_ram[734] = 180;
    exp_47_ram[735] = 196;
    exp_47_ram[736] = 212;
    exp_47_ram[737] = 228;
    exp_47_ram[738] = 4;
    exp_47_ram[739] = 132;
    exp_47_ram[740] = 7;
    exp_47_ram[741] = 64;
    exp_47_ram[742] = 244;
    exp_47_ram[743] = 208;
    exp_47_ram[744] = 4;
    exp_47_ram[745] = 7;
    exp_47_ram[746] = 80;
    exp_47_ram[747] = 247;
    exp_47_ram[748] = 4;
    exp_47_ram[749] = 7;
    exp_47_ram[750] = 196;
    exp_47_ram[751] = 23;
    exp_47_ram[752] = 228;
    exp_47_ram[753] = 196;
    exp_47_ram[754] = 68;
    exp_47_ram[755] = 7;
    exp_47_ram[756] = 132;
    exp_47_ram[757] = 7;
    exp_47_ram[758] = 4;
    exp_47_ram[759] = 23;
    exp_47_ram[760] = 244;
    exp_47_ram[761] = 80;
    exp_47_ram[762] = 4;
    exp_47_ram[763] = 23;
    exp_47_ram[764] = 244;
    exp_47_ram[765] = 4;
    exp_47_ram[766] = 4;
    exp_47_ram[767] = 7;
    exp_47_ram[768] = 7;
    exp_47_ram[769] = 0;
    exp_47_ram[770] = 247;
    exp_47_ram[771] = 39;
    exp_47_ram[772] = 0;
    exp_47_ram[773] = 7;
    exp_47_ram[774] = 247;
    exp_47_ram[775] = 7;
    exp_47_ram[776] = 7;
    exp_47_ram[777] = 196;
    exp_47_ram[778] = 23;
    exp_47_ram[779] = 244;
    exp_47_ram[780] = 4;
    exp_47_ram[781] = 23;
    exp_47_ram[782] = 244;
    exp_47_ram[783] = 16;
    exp_47_ram[784] = 244;
    exp_47_ram[785] = 192;
    exp_47_ram[786] = 196;
    exp_47_ram[787] = 39;
    exp_47_ram[788] = 244;
    exp_47_ram[789] = 4;
    exp_47_ram[790] = 23;
    exp_47_ram[791] = 244;
    exp_47_ram[792] = 16;
    exp_47_ram[793] = 244;
    exp_47_ram[794] = 128;
    exp_47_ram[795] = 196;
    exp_47_ram[796] = 71;
    exp_47_ram[797] = 244;
    exp_47_ram[798] = 4;
    exp_47_ram[799] = 23;
    exp_47_ram[800] = 244;
    exp_47_ram[801] = 16;
    exp_47_ram[802] = 244;
    exp_47_ram[803] = 64;
    exp_47_ram[804] = 196;
    exp_47_ram[805] = 135;
    exp_47_ram[806] = 244;
    exp_47_ram[807] = 4;
    exp_47_ram[808] = 23;
    exp_47_ram[809] = 244;
    exp_47_ram[810] = 16;
    exp_47_ram[811] = 244;
    exp_47_ram[812] = 0;
    exp_47_ram[813] = 196;
    exp_47_ram[814] = 7;
    exp_47_ram[815] = 244;
    exp_47_ram[816] = 4;
    exp_47_ram[817] = 23;
    exp_47_ram[818] = 244;
    exp_47_ram[819] = 16;
    exp_47_ram[820] = 244;
    exp_47_ram[821] = 192;
    exp_47_ram[822] = 4;
    exp_47_ram[823] = 0;
    exp_47_ram[824] = 4;
    exp_47_ram[825] = 7;
    exp_47_ram[826] = 4;
    exp_47_ram[827] = 4;
    exp_47_ram[828] = 7;
    exp_47_ram[829] = 7;
    exp_47_ram[830] = 223;
    exp_47_ram[831] = 5;
    exp_47_ram[832] = 7;
    exp_47_ram[833] = 4;
    exp_47_ram[834] = 7;
    exp_47_ram[835] = 159;
    exp_47_ram[836] = 164;
    exp_47_ram[837] = 0;
    exp_47_ram[838] = 4;
    exp_47_ram[839] = 7;
    exp_47_ram[840] = 160;
    exp_47_ram[841] = 247;
    exp_47_ram[842] = 196;
    exp_47_ram[843] = 71;
    exp_47_ram[844] = 228;
    exp_47_ram[845] = 7;
    exp_47_ram[846] = 244;
    exp_47_ram[847] = 132;
    exp_47_ram[848] = 7;
    exp_47_ram[849] = 196;
    exp_47_ram[850] = 39;
    exp_47_ram[851] = 244;
    exp_47_ram[852] = 132;
    exp_47_ram[853] = 240;
    exp_47_ram[854] = 244;
    exp_47_ram[855] = 192;
    exp_47_ram[856] = 132;
    exp_47_ram[857] = 244;
    exp_47_ram[858] = 4;
    exp_47_ram[859] = 23;
    exp_47_ram[860] = 244;
    exp_47_ram[861] = 4;
    exp_47_ram[862] = 4;
    exp_47_ram[863] = 7;
    exp_47_ram[864] = 224;
    exp_47_ram[865] = 247;
    exp_47_ram[866] = 196;
    exp_47_ram[867] = 7;
    exp_47_ram[868] = 244;
    exp_47_ram[869] = 4;
    exp_47_ram[870] = 23;
    exp_47_ram[871] = 244;
    exp_47_ram[872] = 4;
    exp_47_ram[873] = 7;
    exp_47_ram[874] = 7;
    exp_47_ram[875] = 143;
    exp_47_ram[876] = 5;
    exp_47_ram[877] = 7;
    exp_47_ram[878] = 4;
    exp_47_ram[879] = 7;
    exp_47_ram[880] = 79;
    exp_47_ram[881] = 164;
    exp_47_ram[882] = 64;
    exp_47_ram[883] = 4;
    exp_47_ram[884] = 7;
    exp_47_ram[885] = 160;
    exp_47_ram[886] = 247;
    exp_47_ram[887] = 196;
    exp_47_ram[888] = 71;
    exp_47_ram[889] = 228;
    exp_47_ram[890] = 7;
    exp_47_ram[891] = 244;
    exp_47_ram[892] = 68;
    exp_47_ram[893] = 7;
    exp_47_ram[894] = 0;
    exp_47_ram[895] = 244;
    exp_47_ram[896] = 4;
    exp_47_ram[897] = 23;
    exp_47_ram[898] = 244;
    exp_47_ram[899] = 4;
    exp_47_ram[900] = 7;
    exp_47_ram[901] = 135;
    exp_47_ram[902] = 32;
    exp_47_ram[903] = 247;
    exp_47_ram[904] = 39;
    exp_47_ram[905] = 0;
    exp_47_ram[906] = 71;
    exp_47_ram[907] = 247;
    exp_47_ram[908] = 7;
    exp_47_ram[909] = 7;
    exp_47_ram[910] = 196;
    exp_47_ram[911] = 7;
    exp_47_ram[912] = 244;
    exp_47_ram[913] = 4;
    exp_47_ram[914] = 23;
    exp_47_ram[915] = 244;
    exp_47_ram[916] = 4;
    exp_47_ram[917] = 7;
    exp_47_ram[918] = 192;
    exp_47_ram[919] = 247;
    exp_47_ram[920] = 196;
    exp_47_ram[921] = 7;
    exp_47_ram[922] = 244;
    exp_47_ram[923] = 4;
    exp_47_ram[924] = 23;
    exp_47_ram[925] = 244;
    exp_47_ram[926] = 64;
    exp_47_ram[927] = 196;
    exp_47_ram[928] = 7;
    exp_47_ram[929] = 244;
    exp_47_ram[930] = 4;
    exp_47_ram[931] = 23;
    exp_47_ram[932] = 244;
    exp_47_ram[933] = 4;
    exp_47_ram[934] = 7;
    exp_47_ram[935] = 128;
    exp_47_ram[936] = 247;
    exp_47_ram[937] = 196;
    exp_47_ram[938] = 7;
    exp_47_ram[939] = 244;
    exp_47_ram[940] = 4;
    exp_47_ram[941] = 23;
    exp_47_ram[942] = 244;
    exp_47_ram[943] = 128;
    exp_47_ram[944] = 196;
    exp_47_ram[945] = 7;
    exp_47_ram[946] = 244;
    exp_47_ram[947] = 4;
    exp_47_ram[948] = 23;
    exp_47_ram[949] = 244;
    exp_47_ram[950] = 0;
    exp_47_ram[951] = 196;
    exp_47_ram[952] = 7;
    exp_47_ram[953] = 244;
    exp_47_ram[954] = 4;
    exp_47_ram[955] = 23;
    exp_47_ram[956] = 244;
    exp_47_ram[957] = 64;
    exp_47_ram[958] = 196;
    exp_47_ram[959] = 7;
    exp_47_ram[960] = 244;
    exp_47_ram[961] = 4;
    exp_47_ram[962] = 23;
    exp_47_ram[963] = 244;
    exp_47_ram[964] = 128;
    exp_47_ram[965] = 0;
    exp_47_ram[966] = 0;
    exp_47_ram[967] = 0;
    exp_47_ram[968] = 128;
    exp_47_ram[969] = 0;
    exp_47_ram[970] = 4;
    exp_47_ram[971] = 7;
    exp_47_ram[972] = 183;
    exp_47_ram[973] = 48;
    exp_47_ram[974] = 247;
    exp_47_ram[975] = 39;
    exp_47_ram[976] = 0;
    exp_47_ram[977] = 7;
    exp_47_ram[978] = 247;
    exp_47_ram[979] = 7;
    exp_47_ram[980] = 7;
    exp_47_ram[981] = 4;
    exp_47_ram[982] = 7;
    exp_47_ram[983] = 128;
    exp_47_ram[984] = 247;
    exp_47_ram[985] = 4;
    exp_47_ram[986] = 7;
    exp_47_ram[987] = 128;
    exp_47_ram[988] = 247;
    exp_47_ram[989] = 0;
    exp_47_ram[990] = 244;
    exp_47_ram[991] = 0;
    exp_47_ram[992] = 4;
    exp_47_ram[993] = 7;
    exp_47_ram[994] = 240;
    exp_47_ram[995] = 247;
    exp_47_ram[996] = 128;
    exp_47_ram[997] = 244;
    exp_47_ram[998] = 64;
    exp_47_ram[999] = 4;
    exp_47_ram[1000] = 7;
    exp_47_ram[1001] = 32;
    exp_47_ram[1002] = 247;
    exp_47_ram[1003] = 32;
    exp_47_ram[1004] = 244;
    exp_47_ram[1005] = 128;
    exp_47_ram[1006] = 160;
    exp_47_ram[1007] = 244;
    exp_47_ram[1008] = 196;
    exp_47_ram[1009] = 247;
    exp_47_ram[1010] = 244;
    exp_47_ram[1011] = 4;
    exp_47_ram[1012] = 7;
    exp_47_ram[1013] = 128;
    exp_47_ram[1014] = 247;
    exp_47_ram[1015] = 196;
    exp_47_ram[1016] = 7;
    exp_47_ram[1017] = 244;
    exp_47_ram[1018] = 4;
    exp_47_ram[1019] = 7;
    exp_47_ram[1020] = 144;
    exp_47_ram[1021] = 247;
    exp_47_ram[1022] = 4;
    exp_47_ram[1023] = 7;
    exp_47_ram[1024] = 64;
    exp_47_ram[1025] = 247;
    exp_47_ram[1026] = 196;
    exp_47_ram[1027] = 55;
    exp_47_ram[1028] = 244;
    exp_47_ram[1029] = 196;
    exp_47_ram[1030] = 7;
    exp_47_ram[1031] = 7;
    exp_47_ram[1032] = 196;
    exp_47_ram[1033] = 231;
    exp_47_ram[1034] = 244;
    exp_47_ram[1035] = 4;
    exp_47_ram[1036] = 7;
    exp_47_ram[1037] = 144;
    exp_47_ram[1038] = 247;
    exp_47_ram[1039] = 4;
    exp_47_ram[1040] = 7;
    exp_47_ram[1041] = 64;
    exp_47_ram[1042] = 247;
    exp_47_ram[1043] = 196;
    exp_47_ram[1044] = 7;
    exp_47_ram[1045] = 7;
    exp_47_ram[1046] = 196;
    exp_47_ram[1047] = 7;
    exp_47_ram[1048] = 7;
    exp_47_ram[1049] = 196;
    exp_47_ram[1050] = 71;
    exp_47_ram[1051] = 228;
    exp_47_ram[1052] = 7;
    exp_47_ram[1053] = 244;
    exp_47_ram[1054] = 132;
    exp_47_ram[1055] = 247;
    exp_47_ram[1056] = 132;
    exp_47_ram[1057] = 247;
    exp_47_ram[1058] = 231;
    exp_47_ram[1059] = 7;
    exp_47_ram[1060] = 132;
    exp_47_ram[1061] = 247;
    exp_47_ram[1062] = 247;
    exp_47_ram[1063] = 196;
    exp_47_ram[1064] = 241;
    exp_47_ram[1065] = 132;
    exp_47_ram[1066] = 241;
    exp_47_ram[1067] = 68;
    exp_47_ram[1068] = 132;
    exp_47_ram[1069] = 7;
    exp_47_ram[1070] = 6;
    exp_47_ram[1071] = 68;
    exp_47_ram[1072] = 196;
    exp_47_ram[1073] = 132;
    exp_47_ram[1074] = 196;
    exp_47_ram[1075] = 31;
    exp_47_ram[1076] = 164;
    exp_47_ram[1077] = 192;
    exp_47_ram[1078] = 196;
    exp_47_ram[1079] = 7;
    exp_47_ram[1080] = 7;
    exp_47_ram[1081] = 196;
    exp_47_ram[1082] = 71;
    exp_47_ram[1083] = 228;
    exp_47_ram[1084] = 7;
    exp_47_ram[1085] = 247;
    exp_47_ram[1086] = 192;
    exp_47_ram[1087] = 196;
    exp_47_ram[1088] = 7;
    exp_47_ram[1089] = 7;
    exp_47_ram[1090] = 196;
    exp_47_ram[1091] = 71;
    exp_47_ram[1092] = 228;
    exp_47_ram[1093] = 7;
    exp_47_ram[1094] = 7;
    exp_47_ram[1095] = 7;
    exp_47_ram[1096] = 64;
    exp_47_ram[1097] = 196;
    exp_47_ram[1098] = 71;
    exp_47_ram[1099] = 228;
    exp_47_ram[1100] = 7;
    exp_47_ram[1101] = 244;
    exp_47_ram[1102] = 196;
    exp_47_ram[1103] = 247;
    exp_47_ram[1104] = 196;
    exp_47_ram[1105] = 247;
    exp_47_ram[1106] = 231;
    exp_47_ram[1107] = 7;
    exp_47_ram[1108] = 196;
    exp_47_ram[1109] = 247;
    exp_47_ram[1110] = 247;
    exp_47_ram[1111] = 196;
    exp_47_ram[1112] = 241;
    exp_47_ram[1113] = 132;
    exp_47_ram[1114] = 241;
    exp_47_ram[1115] = 68;
    exp_47_ram[1116] = 132;
    exp_47_ram[1117] = 7;
    exp_47_ram[1118] = 6;
    exp_47_ram[1119] = 68;
    exp_47_ram[1120] = 196;
    exp_47_ram[1121] = 132;
    exp_47_ram[1122] = 196;
    exp_47_ram[1123] = 31;
    exp_47_ram[1124] = 164;
    exp_47_ram[1125] = 192;
    exp_47_ram[1126] = 196;
    exp_47_ram[1127] = 7;
    exp_47_ram[1128] = 7;
    exp_47_ram[1129] = 196;
    exp_47_ram[1130] = 7;
    exp_47_ram[1131] = 7;
    exp_47_ram[1132] = 196;
    exp_47_ram[1133] = 71;
    exp_47_ram[1134] = 228;
    exp_47_ram[1135] = 7;
    exp_47_ram[1136] = 196;
    exp_47_ram[1137] = 241;
    exp_47_ram[1138] = 132;
    exp_47_ram[1139] = 241;
    exp_47_ram[1140] = 68;
    exp_47_ram[1141] = 132;
    exp_47_ram[1142] = 0;
    exp_47_ram[1143] = 68;
    exp_47_ram[1144] = 196;
    exp_47_ram[1145] = 132;
    exp_47_ram[1146] = 196;
    exp_47_ram[1147] = 31;
    exp_47_ram[1148] = 164;
    exp_47_ram[1149] = 192;
    exp_47_ram[1150] = 196;
    exp_47_ram[1151] = 7;
    exp_47_ram[1152] = 7;
    exp_47_ram[1153] = 196;
    exp_47_ram[1154] = 71;
    exp_47_ram[1155] = 228;
    exp_47_ram[1156] = 7;
    exp_47_ram[1157] = 247;
    exp_47_ram[1158] = 192;
    exp_47_ram[1159] = 196;
    exp_47_ram[1160] = 7;
    exp_47_ram[1161] = 7;
    exp_47_ram[1162] = 196;
    exp_47_ram[1163] = 71;
    exp_47_ram[1164] = 228;
    exp_47_ram[1165] = 7;
    exp_47_ram[1166] = 7;
    exp_47_ram[1167] = 7;
    exp_47_ram[1168] = 64;
    exp_47_ram[1169] = 196;
    exp_47_ram[1170] = 71;
    exp_47_ram[1171] = 228;
    exp_47_ram[1172] = 7;
    exp_47_ram[1173] = 244;
    exp_47_ram[1174] = 196;
    exp_47_ram[1175] = 241;
    exp_47_ram[1176] = 132;
    exp_47_ram[1177] = 241;
    exp_47_ram[1178] = 68;
    exp_47_ram[1179] = 132;
    exp_47_ram[1180] = 0;
    exp_47_ram[1181] = 4;
    exp_47_ram[1182] = 68;
    exp_47_ram[1183] = 196;
    exp_47_ram[1184] = 132;
    exp_47_ram[1185] = 196;
    exp_47_ram[1186] = 79;
    exp_47_ram[1187] = 164;
    exp_47_ram[1188] = 4;
    exp_47_ram[1189] = 23;
    exp_47_ram[1190] = 244;
    exp_47_ram[1191] = 192;
    exp_47_ram[1192] = 16;
    exp_47_ram[1193] = 244;
    exp_47_ram[1194] = 196;
    exp_47_ram[1195] = 39;
    exp_47_ram[1196] = 7;
    exp_47_ram[1197] = 128;
    exp_47_ram[1198] = 196;
    exp_47_ram[1199] = 23;
    exp_47_ram[1200] = 228;
    exp_47_ram[1201] = 196;
    exp_47_ram[1202] = 68;
    exp_47_ram[1203] = 7;
    exp_47_ram[1204] = 132;
    exp_47_ram[1205] = 0;
    exp_47_ram[1206] = 7;
    exp_47_ram[1207] = 68;
    exp_47_ram[1208] = 23;
    exp_47_ram[1209] = 228;
    exp_47_ram[1210] = 132;
    exp_47_ram[1211] = 231;
    exp_47_ram[1212] = 196;
    exp_47_ram[1213] = 71;
    exp_47_ram[1214] = 228;
    exp_47_ram[1215] = 7;
    exp_47_ram[1216] = 247;
    exp_47_ram[1217] = 196;
    exp_47_ram[1218] = 23;
    exp_47_ram[1219] = 228;
    exp_47_ram[1220] = 196;
    exp_47_ram[1221] = 68;
    exp_47_ram[1222] = 7;
    exp_47_ram[1223] = 132;
    exp_47_ram[1224] = 7;
    exp_47_ram[1225] = 196;
    exp_47_ram[1226] = 39;
    exp_47_ram[1227] = 7;
    exp_47_ram[1228] = 128;
    exp_47_ram[1229] = 196;
    exp_47_ram[1230] = 23;
    exp_47_ram[1231] = 228;
    exp_47_ram[1232] = 196;
    exp_47_ram[1233] = 68;
    exp_47_ram[1234] = 7;
    exp_47_ram[1235] = 132;
    exp_47_ram[1236] = 0;
    exp_47_ram[1237] = 7;
    exp_47_ram[1238] = 68;
    exp_47_ram[1239] = 23;
    exp_47_ram[1240] = 228;
    exp_47_ram[1241] = 132;
    exp_47_ram[1242] = 231;
    exp_47_ram[1243] = 4;
    exp_47_ram[1244] = 23;
    exp_47_ram[1245] = 244;
    exp_47_ram[1246] = 0;
    exp_47_ram[1247] = 196;
    exp_47_ram[1248] = 71;
    exp_47_ram[1249] = 228;
    exp_47_ram[1250] = 7;
    exp_47_ram[1251] = 244;
    exp_47_ram[1252] = 68;
    exp_47_ram[1253] = 7;
    exp_47_ram[1254] = 68;
    exp_47_ram[1255] = 128;
    exp_47_ram[1256] = 240;
    exp_47_ram[1257] = 7;
    exp_47_ram[1258] = 4;
    exp_47_ram[1259] = 79;
    exp_47_ram[1260] = 164;
    exp_47_ram[1261] = 196;
    exp_47_ram[1262] = 7;
    exp_47_ram[1263] = 7;
    exp_47_ram[1264] = 196;
    exp_47_ram[1265] = 68;
    exp_47_ram[1266] = 247;
    exp_47_ram[1267] = 7;
    exp_47_ram[1268] = 244;
    exp_47_ram[1269] = 196;
    exp_47_ram[1270] = 39;
    exp_47_ram[1271] = 7;
    exp_47_ram[1272] = 128;
    exp_47_ram[1273] = 196;
    exp_47_ram[1274] = 23;
    exp_47_ram[1275] = 228;
    exp_47_ram[1276] = 196;
    exp_47_ram[1277] = 68;
    exp_47_ram[1278] = 7;
    exp_47_ram[1279] = 132;
    exp_47_ram[1280] = 0;
    exp_47_ram[1281] = 7;
    exp_47_ram[1282] = 196;
    exp_47_ram[1283] = 23;
    exp_47_ram[1284] = 228;
    exp_47_ram[1285] = 132;
    exp_47_ram[1286] = 231;
    exp_47_ram[1287] = 64;
    exp_47_ram[1288] = 4;
    exp_47_ram[1289] = 23;
    exp_47_ram[1290] = 228;
    exp_47_ram[1291] = 7;
    exp_47_ram[1292] = 196;
    exp_47_ram[1293] = 23;
    exp_47_ram[1294] = 228;
    exp_47_ram[1295] = 196;
    exp_47_ram[1296] = 68;
    exp_47_ram[1297] = 7;
    exp_47_ram[1298] = 132;
    exp_47_ram[1299] = 7;
    exp_47_ram[1300] = 4;
    exp_47_ram[1301] = 7;
    exp_47_ram[1302] = 7;
    exp_47_ram[1303] = 196;
    exp_47_ram[1304] = 7;
    exp_47_ram[1305] = 7;
    exp_47_ram[1306] = 68;
    exp_47_ram[1307] = 247;
    exp_47_ram[1308] = 228;
    exp_47_ram[1309] = 7;
    exp_47_ram[1310] = 196;
    exp_47_ram[1311] = 39;
    exp_47_ram[1312] = 7;
    exp_47_ram[1313] = 128;
    exp_47_ram[1314] = 196;
    exp_47_ram[1315] = 23;
    exp_47_ram[1316] = 228;
    exp_47_ram[1317] = 196;
    exp_47_ram[1318] = 68;
    exp_47_ram[1319] = 7;
    exp_47_ram[1320] = 132;
    exp_47_ram[1321] = 0;
    exp_47_ram[1322] = 7;
    exp_47_ram[1323] = 196;
    exp_47_ram[1324] = 23;
    exp_47_ram[1325] = 228;
    exp_47_ram[1326] = 132;
    exp_47_ram[1327] = 231;
    exp_47_ram[1328] = 4;
    exp_47_ram[1329] = 23;
    exp_47_ram[1330] = 244;
    exp_47_ram[1331] = 192;
    exp_47_ram[1332] = 128;
    exp_47_ram[1333] = 244;
    exp_47_ram[1334] = 196;
    exp_47_ram[1335] = 23;
    exp_47_ram[1336] = 244;
    exp_47_ram[1337] = 196;
    exp_47_ram[1338] = 71;
    exp_47_ram[1339] = 228;
    exp_47_ram[1340] = 7;
    exp_47_ram[1341] = 7;
    exp_47_ram[1342] = 196;
    exp_47_ram[1343] = 241;
    exp_47_ram[1344] = 132;
    exp_47_ram[1345] = 241;
    exp_47_ram[1346] = 68;
    exp_47_ram[1347] = 0;
    exp_47_ram[1348] = 0;
    exp_47_ram[1349] = 68;
    exp_47_ram[1350] = 196;
    exp_47_ram[1351] = 132;
    exp_47_ram[1352] = 196;
    exp_47_ram[1353] = 143;
    exp_47_ram[1354] = 164;
    exp_47_ram[1355] = 4;
    exp_47_ram[1356] = 23;
    exp_47_ram[1357] = 244;
    exp_47_ram[1358] = 0;
    exp_47_ram[1359] = 196;
    exp_47_ram[1360] = 23;
    exp_47_ram[1361] = 228;
    exp_47_ram[1362] = 196;
    exp_47_ram[1363] = 68;
    exp_47_ram[1364] = 7;
    exp_47_ram[1365] = 132;
    exp_47_ram[1366] = 80;
    exp_47_ram[1367] = 7;
    exp_47_ram[1368] = 4;
    exp_47_ram[1369] = 23;
    exp_47_ram[1370] = 244;
    exp_47_ram[1371] = 192;
    exp_47_ram[1372] = 4;
    exp_47_ram[1373] = 7;
    exp_47_ram[1374] = 196;
    exp_47_ram[1375] = 23;
    exp_47_ram[1376] = 228;
    exp_47_ram[1377] = 196;
    exp_47_ram[1378] = 68;
    exp_47_ram[1379] = 7;
    exp_47_ram[1380] = 132;
    exp_47_ram[1381] = 7;
    exp_47_ram[1382] = 4;
    exp_47_ram[1383] = 23;
    exp_47_ram[1384] = 244;
    exp_47_ram[1385] = 0;
    exp_47_ram[1386] = 4;
    exp_47_ram[1387] = 7;
    exp_47_ram[1388] = 7;
    exp_47_ram[1389] = 196;
    exp_47_ram[1390] = 68;
    exp_47_ram[1391] = 247;
    exp_47_ram[1392] = 68;
    exp_47_ram[1393] = 247;
    exp_47_ram[1394] = 128;
    exp_47_ram[1395] = 196;
    exp_47_ram[1396] = 196;
    exp_47_ram[1397] = 68;
    exp_47_ram[1398] = 7;
    exp_47_ram[1399] = 132;
    exp_47_ram[1400] = 0;
    exp_47_ram[1401] = 7;
    exp_47_ram[1402] = 196;
    exp_47_ram[1403] = 7;
    exp_47_ram[1404] = 193;
    exp_47_ram[1405] = 129;
    exp_47_ram[1406] = 1;
    exp_47_ram[1407] = 0;
    exp_47_ram[1408] = 1;
    exp_47_ram[1409] = 17;
    exp_47_ram[1410] = 129;
    exp_47_ram[1411] = 1;
    exp_47_ram[1412] = 164;
    exp_47_ram[1413] = 180;
    exp_47_ram[1414] = 196;
    exp_47_ram[1415] = 212;
    exp_47_ram[1416] = 228;
    exp_47_ram[1417] = 244;
    exp_47_ram[1418] = 4;
    exp_47_ram[1419] = 20;
    exp_47_ram[1420] = 4;
    exp_47_ram[1421] = 244;
    exp_47_ram[1422] = 132;
    exp_47_ram[1423] = 71;
    exp_47_ram[1424] = 244;
    exp_47_ram[1425] = 132;
    exp_47_ram[1426] = 68;
    exp_47_ram[1427] = 196;
    exp_47_ram[1428] = 240;
    exp_47_ram[1429] = 7;
    exp_47_ram[1430] = 64;
    exp_47_ram[1431] = 143;
    exp_47_ram[1432] = 164;
    exp_47_ram[1433] = 196;
    exp_47_ram[1434] = 7;
    exp_47_ram[1435] = 193;
    exp_47_ram[1436] = 129;
    exp_47_ram[1437] = 1;
    exp_47_ram[1438] = 0;
    exp_47_ram[1439] = 1;
    exp_47_ram[1440] = 17;
    exp_47_ram[1441] = 129;
    exp_47_ram[1442] = 1;
    exp_47_ram[1443] = 5;
    exp_47_ram[1444] = 244;
    exp_47_ram[1445] = 244;
    exp_47_ram[1446] = 0;
    exp_47_ram[1447] = 199;
    exp_47_ram[1448] = 7;
    exp_47_ram[1449] = 7;
    exp_47_ram[1450] = 159;
    exp_47_ram[1451] = 0;
    exp_47_ram[1452] = 193;
    exp_47_ram[1453] = 129;
    exp_47_ram[1454] = 1;
    exp_47_ram[1455] = 0;
    exp_47_ram[1456] = 1;
    exp_47_ram[1457] = 17;
    exp_47_ram[1458] = 129;
    exp_47_ram[1459] = 1;
    exp_47_ram[1460] = 192;
    exp_47_ram[1461] = 159;
    exp_47_ram[1462] = 0;
    exp_47_ram[1463] = 64;
    exp_47_ram[1464] = 7;
    exp_47_ram[1465] = 7;
    exp_47_ram[1466] = 192;
    exp_47_ram[1467] = 95;
    exp_47_ram[1468] = 128;
    exp_47_ram[1469] = 192;
    exp_47_ram[1470] = 7;
    exp_47_ram[1471] = 7;
    exp_47_ram[1472] = 192;
    exp_47_ram[1473] = 223;
    exp_47_ram[1474] = 0;
    exp_47_ram[1475] = 64;
    exp_47_ram[1476] = 7;
    exp_47_ram[1477] = 7;
    exp_47_ram[1478] = 192;
    exp_47_ram[1479] = 95;
    exp_47_ram[1480] = 128;
    exp_47_ram[1481] = 192;
    exp_47_ram[1482] = 7;
    exp_47_ram[1483] = 7;
    exp_47_ram[1484] = 192;
    exp_47_ram[1485] = 223;
    exp_47_ram[1486] = 0;
    exp_47_ram[1487] = 64;
    exp_47_ram[1488] = 7;
    exp_47_ram[1489] = 7;
    exp_47_ram[1490] = 192;
    exp_47_ram[1491] = 95;
    exp_47_ram[1492] = 128;
    exp_47_ram[1493] = 192;
    exp_47_ram[1494] = 7;
    exp_47_ram[1495] = 7;
    exp_47_ram[1496] = 192;
    exp_47_ram[1497] = 223;
    exp_47_ram[1498] = 0;
    exp_47_ram[1499] = 0;
    exp_47_ram[1500] = 192;
    exp_47_ram[1501] = 223;
    exp_47_ram[1502] = 0;
    exp_47_ram[1503] = 64;
    exp_47_ram[1504] = 7;
    exp_47_ram[1505] = 7;
    exp_47_ram[1506] = 192;
    exp_47_ram[1507] = 95;
    exp_47_ram[1508] = 128;
    exp_47_ram[1509] = 192;
    exp_47_ram[1510] = 7;
    exp_47_ram[1511] = 7;
    exp_47_ram[1512] = 192;
    exp_47_ram[1513] = 223;
    exp_47_ram[1514] = 0;
    exp_47_ram[1515] = 64;
    exp_47_ram[1516] = 7;
    exp_47_ram[1517] = 7;
    exp_47_ram[1518] = 192;
    exp_47_ram[1519] = 95;
    exp_47_ram[1520] = 128;
    exp_47_ram[1521] = 192;
    exp_47_ram[1522] = 7;
    exp_47_ram[1523] = 7;
    exp_47_ram[1524] = 192;
    exp_47_ram[1525] = 223;
    exp_47_ram[1526] = 0;
    exp_47_ram[1527] = 64;
    exp_47_ram[1528] = 7;
    exp_47_ram[1529] = 7;
    exp_47_ram[1530] = 192;
    exp_47_ram[1531] = 95;
    exp_47_ram[1532] = 128;
    exp_47_ram[1533] = 192;
    exp_47_ram[1534] = 7;
    exp_47_ram[1535] = 7;
    exp_47_ram[1536] = 192;
    exp_47_ram[1537] = 223;
    exp_47_ram[1538] = 0;
    exp_47_ram[1539] = 64;
    exp_47_ram[1540] = 7;
    exp_47_ram[1541] = 7;
    exp_47_ram[1542] = 0;
    exp_47_ram[1543] = 95;
    exp_47_ram[1544] = 128;
    exp_47_ram[1545] = 192;
    exp_47_ram[1546] = 7;
    exp_47_ram[1547] = 7;
    exp_47_ram[1548] = 0;
    exp_47_ram[1549] = 223;
    exp_47_ram[1550] = 0;
    exp_47_ram[1551] = 64;
    exp_47_ram[1552] = 7;
    exp_47_ram[1553] = 7;
    exp_47_ram[1554] = 0;
    exp_47_ram[1555] = 95;
    exp_47_ram[1556] = 128;
    exp_47_ram[1557] = 192;
    exp_47_ram[1558] = 7;
    exp_47_ram[1559] = 7;
    exp_47_ram[1560] = 0;
    exp_47_ram[1561] = 223;
    exp_47_ram[1562] = 0;
    exp_47_ram[1563] = 64;
    exp_47_ram[1564] = 7;
    exp_47_ram[1565] = 7;
    exp_47_ram[1566] = 0;
    exp_47_ram[1567] = 95;
    exp_47_ram[1568] = 128;
    exp_47_ram[1569] = 192;
    exp_47_ram[1570] = 7;
    exp_47_ram[1571] = 7;
    exp_47_ram[1572] = 0;
    exp_47_ram[1573] = 223;
    exp_47_ram[1574] = 0;
    exp_47_ram[1575] = 0;
    exp_47_ram[1576] = 0;
    exp_47_ram[1577] = 223;
    exp_47_ram[1578] = 0;
    exp_47_ram[1579] = 64;
    exp_47_ram[1580] = 7;
    exp_47_ram[1581] = 7;
    exp_47_ram[1582] = 0;
    exp_47_ram[1583] = 95;
    exp_47_ram[1584] = 128;
    exp_47_ram[1585] = 192;
    exp_47_ram[1586] = 7;
    exp_47_ram[1587] = 7;
    exp_47_ram[1588] = 0;
    exp_47_ram[1589] = 223;
    exp_47_ram[1590] = 0;
    exp_47_ram[1591] = 64;
    exp_47_ram[1592] = 7;
    exp_47_ram[1593] = 7;
    exp_47_ram[1594] = 0;
    exp_47_ram[1595] = 95;
    exp_47_ram[1596] = 128;
    exp_47_ram[1597] = 192;
    exp_47_ram[1598] = 7;
    exp_47_ram[1599] = 7;
    exp_47_ram[1600] = 0;
    exp_47_ram[1601] = 223;
    exp_47_ram[1602] = 0;
    exp_47_ram[1603] = 64;
    exp_47_ram[1604] = 7;
    exp_47_ram[1605] = 7;
    exp_47_ram[1606] = 0;
    exp_47_ram[1607] = 95;
    exp_47_ram[1608] = 128;
    exp_47_ram[1609] = 192;
    exp_47_ram[1610] = 7;
    exp_47_ram[1611] = 7;
    exp_47_ram[1612] = 0;
    exp_47_ram[1613] = 223;
    exp_47_ram[1614] = 0;
    exp_47_ram[1615] = 64;
    exp_47_ram[1616] = 7;
    exp_47_ram[1617] = 7;
    exp_47_ram[1618] = 192;
    exp_47_ram[1619] = 95;
    exp_47_ram[1620] = 128;
    exp_47_ram[1621] = 192;
    exp_47_ram[1622] = 7;
    exp_47_ram[1623] = 7;
    exp_47_ram[1624] = 192;
    exp_47_ram[1625] = 223;
    exp_47_ram[1626] = 0;
    exp_47_ram[1627] = 64;
    exp_47_ram[1628] = 7;
    exp_47_ram[1629] = 7;
    exp_47_ram[1630] = 192;
    exp_47_ram[1631] = 95;
    exp_47_ram[1632] = 128;
    exp_47_ram[1633] = 192;
    exp_47_ram[1634] = 7;
    exp_47_ram[1635] = 7;
    exp_47_ram[1636] = 192;
    exp_47_ram[1637] = 223;
    exp_47_ram[1638] = 0;
    exp_47_ram[1639] = 64;
    exp_47_ram[1640] = 7;
    exp_47_ram[1641] = 7;
    exp_47_ram[1642] = 192;
    exp_47_ram[1643] = 95;
    exp_47_ram[1644] = 128;
    exp_47_ram[1645] = 192;
    exp_47_ram[1646] = 7;
    exp_47_ram[1647] = 7;
    exp_47_ram[1648] = 192;
    exp_47_ram[1649] = 223;
    exp_47_ram[1650] = 0;
    exp_47_ram[1651] = 0;
    exp_47_ram[1652] = 192;
    exp_47_ram[1653] = 223;
    exp_47_ram[1654] = 0;
    exp_47_ram[1655] = 64;
    exp_47_ram[1656] = 7;
    exp_47_ram[1657] = 7;
    exp_47_ram[1658] = 192;
    exp_47_ram[1659] = 95;
    exp_47_ram[1660] = 128;
    exp_47_ram[1661] = 192;
    exp_47_ram[1662] = 7;
    exp_47_ram[1663] = 7;
    exp_47_ram[1664] = 192;
    exp_47_ram[1665] = 223;
    exp_47_ram[1666] = 0;
    exp_47_ram[1667] = 64;
    exp_47_ram[1668] = 7;
    exp_47_ram[1669] = 7;
    exp_47_ram[1670] = 192;
    exp_47_ram[1671] = 95;
    exp_47_ram[1672] = 128;
    exp_47_ram[1673] = 192;
    exp_47_ram[1674] = 7;
    exp_47_ram[1675] = 7;
    exp_47_ram[1676] = 192;
    exp_47_ram[1677] = 223;
    exp_47_ram[1678] = 0;
    exp_47_ram[1679] = 64;
    exp_47_ram[1680] = 7;
    exp_47_ram[1681] = 7;
    exp_47_ram[1682] = 192;
    exp_47_ram[1683] = 95;
    exp_47_ram[1684] = 128;
    exp_47_ram[1685] = 192;
    exp_47_ram[1686] = 7;
    exp_47_ram[1687] = 7;
    exp_47_ram[1688] = 192;
    exp_47_ram[1689] = 223;
    exp_47_ram[1690] = 0;
    exp_47_ram[1691] = 64;
    exp_47_ram[1692] = 7;
    exp_47_ram[1693] = 7;
    exp_47_ram[1694] = 0;
    exp_47_ram[1695] = 95;
    exp_47_ram[1696] = 128;
    exp_47_ram[1697] = 192;
    exp_47_ram[1698] = 7;
    exp_47_ram[1699] = 7;
    exp_47_ram[1700] = 0;
    exp_47_ram[1701] = 223;
    exp_47_ram[1702] = 0;
    exp_47_ram[1703] = 64;
    exp_47_ram[1704] = 7;
    exp_47_ram[1705] = 7;
    exp_47_ram[1706] = 0;
    exp_47_ram[1707] = 95;
    exp_47_ram[1708] = 128;
    exp_47_ram[1709] = 192;
    exp_47_ram[1710] = 7;
    exp_47_ram[1711] = 7;
    exp_47_ram[1712] = 0;
    exp_47_ram[1713] = 223;
    exp_47_ram[1714] = 0;
    exp_47_ram[1715] = 64;
    exp_47_ram[1716] = 7;
    exp_47_ram[1717] = 7;
    exp_47_ram[1718] = 0;
    exp_47_ram[1719] = 95;
    exp_47_ram[1720] = 128;
    exp_47_ram[1721] = 192;
    exp_47_ram[1722] = 7;
    exp_47_ram[1723] = 7;
    exp_47_ram[1724] = 0;
    exp_47_ram[1725] = 223;
    exp_47_ram[1726] = 0;
    exp_47_ram[1727] = 0;
    exp_47_ram[1728] = 0;
    exp_47_ram[1729] = 223;
    exp_47_ram[1730] = 0;
    exp_47_ram[1731] = 64;
    exp_47_ram[1732] = 7;
    exp_47_ram[1733] = 7;
    exp_47_ram[1734] = 0;
    exp_47_ram[1735] = 95;
    exp_47_ram[1736] = 128;
    exp_47_ram[1737] = 192;
    exp_47_ram[1738] = 7;
    exp_47_ram[1739] = 7;
    exp_47_ram[1740] = 0;
    exp_47_ram[1741] = 223;
    exp_47_ram[1742] = 0;
    exp_47_ram[1743] = 64;
    exp_47_ram[1744] = 7;
    exp_47_ram[1745] = 7;
    exp_47_ram[1746] = 0;
    exp_47_ram[1747] = 95;
    exp_47_ram[1748] = 128;
    exp_47_ram[1749] = 192;
    exp_47_ram[1750] = 7;
    exp_47_ram[1751] = 7;
    exp_47_ram[1752] = 0;
    exp_47_ram[1753] = 223;
    exp_47_ram[1754] = 0;
    exp_47_ram[1755] = 64;
    exp_47_ram[1756] = 7;
    exp_47_ram[1757] = 7;
    exp_47_ram[1758] = 0;
    exp_47_ram[1759] = 95;
    exp_47_ram[1760] = 128;
    exp_47_ram[1761] = 192;
    exp_47_ram[1762] = 7;
    exp_47_ram[1763] = 7;
    exp_47_ram[1764] = 0;
    exp_47_ram[1765] = 223;
    exp_47_ram[1766] = 0;
    exp_47_ram[1767] = 64;
    exp_47_ram[1768] = 7;
    exp_47_ram[1769] = 7;
    exp_47_ram[1770] = 0;
    exp_47_ram[1771] = 95;
    exp_47_ram[1772] = 128;
    exp_47_ram[1773] = 192;
    exp_47_ram[1774] = 7;
    exp_47_ram[1775] = 7;
    exp_47_ram[1776] = 0;
    exp_47_ram[1777] = 223;
    exp_47_ram[1778] = 0;
    exp_47_ram[1779] = 64;
    exp_47_ram[1780] = 7;
    exp_47_ram[1781] = 7;
    exp_47_ram[1782] = 0;
    exp_47_ram[1783] = 95;
    exp_47_ram[1784] = 128;
    exp_47_ram[1785] = 192;
    exp_47_ram[1786] = 7;
    exp_47_ram[1787] = 7;
    exp_47_ram[1788] = 0;
    exp_47_ram[1789] = 223;
    exp_47_ram[1790] = 0;
    exp_47_ram[1791] = 64;
    exp_47_ram[1792] = 7;
    exp_47_ram[1793] = 7;
    exp_47_ram[1794] = 192;
    exp_47_ram[1795] = 95;
    exp_47_ram[1796] = 0;
    exp_47_ram[1797] = 64;
    exp_47_ram[1798] = 7;
    exp_47_ram[1799] = 7;
    exp_47_ram[1800] = 64;
    exp_47_ram[1801] = 223;
    exp_47_ram[1802] = 0;
    exp_47_ram[1803] = 64;
    exp_47_ram[1804] = 7;
    exp_47_ram[1805] = 7;
    exp_47_ram[1806] = 128;
    exp_47_ram[1807] = 95;
    exp_47_ram[1808] = 0;
    exp_47_ram[1809] = 64;
    exp_47_ram[1810] = 7;
    exp_47_ram[1811] = 7;
    exp_47_ram[1812] = 192;
    exp_47_ram[1813] = 223;
    exp_47_ram[1814] = 128;
    exp_47_ram[1815] = 192;
    exp_47_ram[1816] = 7;
    exp_47_ram[1817] = 7;
    exp_47_ram[1818] = 192;
    exp_47_ram[1819] = 95;
    exp_47_ram[1820] = 128;
    exp_47_ram[1821] = 192;
    exp_47_ram[1822] = 7;
    exp_47_ram[1823] = 7;
    exp_47_ram[1824] = 64;
    exp_47_ram[1825] = 223;
    exp_47_ram[1826] = 128;
    exp_47_ram[1827] = 192;
    exp_47_ram[1828] = 7;
    exp_47_ram[1829] = 7;
    exp_47_ram[1830] = 128;
    exp_47_ram[1831] = 95;
    exp_47_ram[1832] = 128;
    exp_47_ram[1833] = 192;
    exp_47_ram[1834] = 7;
    exp_47_ram[1835] = 7;
    exp_47_ram[1836] = 192;
    exp_47_ram[1837] = 223;
    exp_47_ram[1838] = 0;
    exp_47_ram[1839] = 64;
    exp_47_ram[1840] = 7;
    exp_47_ram[1841] = 7;
    exp_47_ram[1842] = 192;
    exp_47_ram[1843] = 95;
    exp_47_ram[1844] = 0;
    exp_47_ram[1845] = 64;
    exp_47_ram[1846] = 7;
    exp_47_ram[1847] = 7;
    exp_47_ram[1848] = 64;
    exp_47_ram[1849] = 223;
    exp_47_ram[1850] = 0;
    exp_47_ram[1851] = 64;
    exp_47_ram[1852] = 7;
    exp_47_ram[1853] = 7;
    exp_47_ram[1854] = 128;
    exp_47_ram[1855] = 95;
    exp_47_ram[1856] = 0;
    exp_47_ram[1857] = 64;
    exp_47_ram[1858] = 7;
    exp_47_ram[1859] = 7;
    exp_47_ram[1860] = 192;
    exp_47_ram[1861] = 223;
    exp_47_ram[1862] = 128;
    exp_47_ram[1863] = 192;
    exp_47_ram[1864] = 7;
    exp_47_ram[1865] = 7;
    exp_47_ram[1866] = 192;
    exp_47_ram[1867] = 95;
    exp_47_ram[1868] = 128;
    exp_47_ram[1869] = 192;
    exp_47_ram[1870] = 7;
    exp_47_ram[1871] = 7;
    exp_47_ram[1872] = 64;
    exp_47_ram[1873] = 223;
    exp_47_ram[1874] = 128;
    exp_47_ram[1875] = 192;
    exp_47_ram[1876] = 7;
    exp_47_ram[1877] = 7;
    exp_47_ram[1878] = 128;
    exp_47_ram[1879] = 95;
    exp_47_ram[1880] = 128;
    exp_47_ram[1881] = 192;
    exp_47_ram[1882] = 7;
    exp_47_ram[1883] = 7;
    exp_47_ram[1884] = 192;
    exp_47_ram[1885] = 223;
    exp_47_ram[1886] = 192;
    exp_47_ram[1887] = 15;
    exp_47_ram[1888] = 0;
    exp_47_ram[1889] = 193;
    exp_47_ram[1890] = 129;
    exp_47_ram[1891] = 1;
    exp_47_ram[1892] = 0;
    exp_47_ram[1893] = 1;
    exp_47_ram[1894] = 17;
    exp_47_ram[1895] = 129;
    exp_47_ram[1896] = 1;
    exp_47_ram[1897] = 223;
    exp_47_ram[1898] = 0;
    exp_47_ram[1899] = 193;
    exp_47_ram[1900] = 129;
    exp_47_ram[1901] = 1;
    exp_47_ram[1902] = 0;
    exp_47_ram[1903] = 0;
    exp_47_ram[1904] = 0;
    exp_47_ram[1905] = 0;
    exp_47_ram[1906] = 0;
    exp_47_ram[1907] = 0;
    exp_47_ram[1908] = 0;
    exp_47_ram[1909] = 0;
    exp_47_ram[1910] = 0;
    exp_47_ram[1911] = 0;
    exp_47_ram[1912] = 0;
    exp_47_ram[1913] = 0;
    exp_47_ram[1914] = 0;
    exp_47_ram[1915] = 0;
    exp_47_ram[1916] = 0;
    exp_47_ram[1917] = 0;
    exp_47_ram[1918] = 0;
    exp_47_ram[1919] = 0;
    exp_47_ram[1920] = 0;
    exp_47_ram[1921] = 0;
    exp_47_ram[1922] = 0;
    exp_47_ram[1923] = 0;
    exp_47_ram[1924] = 0;
    exp_47_ram[1925] = 0;
    exp_47_ram[1926] = 0;
    exp_47_ram[1927] = 0;
    exp_47_ram[1928] = 0;
    exp_47_ram[1929] = 0;
    exp_47_ram[1930] = 0;
    exp_47_ram[1931] = 0;
    exp_47_ram[1932] = 0;
    exp_47_ram[1933] = 0;
    exp_47_ram[1934] = 0;
    exp_47_ram[1935] = 0;
    exp_47_ram[1936] = 0;
    exp_47_ram[1937] = 0;
    exp_47_ram[1938] = 0;
    exp_47_ram[1939] = 0;
    exp_47_ram[1940] = 0;
    exp_47_ram[1941] = 0;
    exp_47_ram[1942] = 0;
    exp_47_ram[1943] = 0;
    exp_47_ram[1944] = 0;
    exp_47_ram[1945] = 0;
    exp_47_ram[1946] = 0;
    exp_47_ram[1947] = 0;
    exp_47_ram[1948] = 0;
    exp_47_ram[1949] = 0;
    exp_47_ram[1950] = 0;
    exp_47_ram[1951] = 0;
    exp_47_ram[1952] = 0;
    exp_47_ram[1953] = 0;
    exp_47_ram[1954] = 0;
    exp_47_ram[1955] = 0;
    exp_47_ram[1956] = 0;
    exp_47_ram[1957] = 0;
    exp_47_ram[1958] = 0;
    exp_47_ram[1959] = 0;
    exp_47_ram[1960] = 0;
    exp_47_ram[1961] = 0;
    exp_47_ram[1962] = 0;
    exp_47_ram[1963] = 0;
    exp_47_ram[1964] = 0;
    exp_47_ram[1965] = 0;
    exp_47_ram[1966] = 0;
    exp_47_ram[1967] = 0;
    exp_47_ram[1968] = 0;
    exp_47_ram[1969] = 0;
    exp_47_ram[1970] = 0;
    exp_47_ram[1971] = 0;
    exp_47_ram[1972] = 0;
    exp_47_ram[1973] = 0;
    exp_47_ram[1974] = 0;
    exp_47_ram[1975] = 0;
    exp_47_ram[1976] = 0;
    exp_47_ram[1977] = 0;
    exp_47_ram[1978] = 0;
    exp_47_ram[1979] = 0;
    exp_47_ram[1980] = 0;
    exp_47_ram[1981] = 0;
    exp_47_ram[1982] = 0;
    exp_47_ram[1983] = 0;
    exp_47_ram[1984] = 0;
    exp_47_ram[1985] = 0;
    exp_47_ram[1986] = 0;
    exp_47_ram[1987] = 0;
    exp_47_ram[1988] = 0;
    exp_47_ram[1989] = 0;
    exp_47_ram[1990] = 0;
    exp_47_ram[1991] = 0;
    exp_47_ram[1992] = 0;
    exp_47_ram[1993] = 0;
    exp_47_ram[1994] = 0;
    exp_47_ram[1995] = 0;
    exp_47_ram[1996] = 0;
    exp_47_ram[1997] = 0;
    exp_47_ram[1998] = 0;
    exp_47_ram[1999] = 0;
    exp_47_ram[2000] = 0;
    exp_47_ram[2001] = 0;
    exp_47_ram[2002] = 0;
    exp_47_ram[2003] = 0;
    exp_47_ram[2004] = 0;
    exp_47_ram[2005] = 0;
    exp_47_ram[2006] = 0;
    exp_47_ram[2007] = 0;
    exp_47_ram[2008] = 0;
    exp_47_ram[2009] = 0;
    exp_47_ram[2010] = 0;
    exp_47_ram[2011] = 0;
    exp_47_ram[2012] = 0;
    exp_47_ram[2013] = 0;
    exp_47_ram[2014] = 0;
    exp_47_ram[2015] = 0;
    exp_47_ram[2016] = 0;
    exp_47_ram[2017] = 0;
    exp_47_ram[2018] = 0;
    exp_47_ram[2019] = 0;
    exp_47_ram[2020] = 0;
    exp_47_ram[2021] = 0;
    exp_47_ram[2022] = 0;
    exp_47_ram[2023] = 0;
    exp_47_ram[2024] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 81;
    exp_40_ram[32] = 1;
    exp_40_ram[33] = 16;
    exp_40_ram[34] = 0;
    exp_40_ram[35] = 0;
    exp_40_ram[36] = 116;
    exp_40_ram[37] = 116;
    exp_40_ram[38] = 0;
    exp_40_ram[39] = 108;
    exp_40_ram[40] = 101;
    exp_40_ram[41] = 0;
    exp_40_ram[42] = 32;
    exp_40_ram[43] = 108;
    exp_40_ram[44] = 32;
    exp_40_ram[45] = 108;
    exp_40_ram[46] = 101;
    exp_40_ram[47] = 32;
    exp_40_ram[48] = 108;
    exp_40_ram[49] = 32;
    exp_40_ram[50] = 108;
    exp_40_ram[51] = 97;
    exp_40_ram[52] = 0;
    exp_40_ram[53] = 116;
    exp_40_ram[54] = 97;
    exp_40_ram[55] = 46;
    exp_40_ram[56] = 108;
    exp_40_ram[57] = 122;
    exp_40_ram[58] = 101;
    exp_40_ram[59] = 112;
    exp_40_ram[60] = 0;
    exp_40_ram[61] = 116;
    exp_40_ram[62] = 112;
    exp_40_ram[63] = 0;
    exp_40_ram[64] = 116;
    exp_40_ram[65] = 109;
    exp_40_ram[66] = 46;
    exp_40_ram[67] = 101;
    exp_40_ram[68] = 114;
    exp_40_ram[69] = 0;
    exp_40_ram[70] = 32;
    exp_40_ram[71] = 108;
    exp_40_ram[72] = 116;
    exp_40_ram[73] = 114;
    exp_40_ram[74] = 0;
    exp_40_ram[75] = 32;
    exp_40_ram[76] = 108;
    exp_40_ram[77] = 116;
    exp_40_ram[78] = 112;
    exp_40_ram[79] = 46;
    exp_40_ram[80] = 115;
    exp_40_ram[81] = 0;
    exp_40_ram[82] = 115;
    exp_40_ram[83] = 115;
    exp_40_ram[84] = 0;
    exp_40_ram[85] = 115;
    exp_40_ram[86] = 115;
    exp_40_ram[87] = 0;
    exp_40_ram[88] = 115;
    exp_40_ram[89] = 100;
    exp_40_ram[90] = 0;
    exp_40_ram[91] = 115;
    exp_40_ram[92] = 115;
    exp_40_ram[93] = 0;
    exp_40_ram[94] = 116;
    exp_40_ram[95] = 114;
    exp_40_ram[96] = 46;
    exp_40_ram[97] = 115;
    exp_40_ram[98] = 115;
    exp_40_ram[99] = 0;
    exp_40_ram[100] = 100;
    exp_40_ram[101] = 115;
    exp_40_ram[102] = 107;
    exp_40_ram[103] = 107;
    exp_40_ram[104] = 97;
    exp_40_ram[105] = 0;
    exp_40_ram[106] = 115;
    exp_40_ram[107] = 115;
    exp_40_ram[108] = 0;
    exp_40_ram[109] = 116;
    exp_40_ram[110] = 104;
    exp_40_ram[111] = 46;
    exp_40_ram[112] = 116;
    exp_40_ram[113] = 110;
    exp_40_ram[114] = 0;
    exp_40_ram[115] = 115;
    exp_40_ram[116] = 102;
    exp_40_ram[117] = 115;
    exp_40_ram[118] = 49;
    exp_40_ram[119] = 102;
    exp_40_ram[120] = 115;
    exp_40_ram[121] = 97;
    exp_40_ram[122] = 102;
    exp_40_ram[123] = 115;
    exp_40_ram[124] = 50;
    exp_40_ram[125] = 51;
    exp_40_ram[126] = 0;
    exp_40_ram[127] = 116;
    exp_40_ram[128] = 114;
    exp_40_ram[129] = 0;
    exp_40_ram[130] = 50;
    exp_40_ram[131] = 0;
    exp_40_ram[132] = 51;
    exp_40_ram[133] = 52;
    exp_40_ram[134] = 101;
    exp_40_ram[135] = 116;
    exp_40_ram[136] = 0;
    exp_40_ram[137] = 50;
    exp_40_ram[138] = 0;
    exp_40_ram[139] = 98;
    exp_40_ram[140] = 0;
    exp_40_ram[141] = 99;
    exp_40_ram[142] = 0;
    exp_40_ram[143] = 100;
    exp_40_ram[144] = 0;
    exp_40_ram[145] = 116;
    exp_40_ram[146] = 110;
    exp_40_ram[147] = 0;
    exp_40_ram[148] = 105;
    exp_40_ram[149] = 46;
    exp_40_ram[150] = 104;
    exp_40_ram[151] = 101;
    exp_40_ram[152] = 55;
    exp_40_ram[153] = 58;
    exp_40_ram[154] = 48;
    exp_40_ram[155] = 48;
    exp_40_ram[156] = 0;
    exp_40_ram[157] = 104;
    exp_40_ram[158] = 101;
    exp_40_ram[159] = 55;
    exp_40_ram[160] = 58;
    exp_40_ram[161] = 48;
    exp_40_ram[162] = 48;
    exp_40_ram[163] = 0;
    exp_40_ram[164] = 32;
    exp_40_ram[165] = 108;
    exp_40_ram[166] = 32;
    exp_40_ram[167] = 108;
    exp_40_ram[168] = 32;
    exp_40_ram[169] = 108;
    exp_40_ram[170] = 104;
    exp_40_ram[171] = 101;
    exp_40_ram[172] = 55;
    exp_40_ram[173] = 58;
    exp_40_ram[174] = 48;
    exp_40_ram[175] = 48;
    exp_40_ram[176] = 0;
    exp_40_ram[177] = 48;
    exp_40_ram[178] = 105;
    exp_40_ram[179] = 49;
    exp_40_ram[180] = 105;
    exp_40_ram[181] = 50;
    exp_40_ram[182] = 105;
    exp_40_ram[183] = 101;
    exp_40_ram[184] = 112;
    exp_40_ram[185] = 116;
    exp_40_ram[186] = 46;
    exp_40_ram[187] = 102;
    exp_40_ram[188] = 50;
    exp_40_ram[189] = 48;
    exp_40_ram[190] = 0;
    exp_40_ram[191] = 101;
    exp_40_ram[192] = 105;
    exp_40_ram[193] = 32;
    exp_40_ram[194] = 37;
    exp_40_ram[195] = 52;
    exp_40_ram[196] = 0;
    exp_40_ram[197] = 69;
    exp_40_ram[198] = 103;
    exp_40_ram[199] = 71;
    exp_40_ram[200] = 237;
    exp_40_ram[201] = 198;
    exp_40_ram[202] = 104;
    exp_40_ram[203] = 248;
    exp_40_ram[204] = 67;
    exp_40_ram[205] = 54;
    exp_40_ram[206] = 169;
    exp_40_ram[207] = 98;
    exp_40_ram[208] = 20;
    exp_40_ram[209] = 122;
    exp_40_ram[210] = 153;
    exp_40_ram[211] = 153;
    exp_40_ram[212] = 0;
    exp_40_ram[213] = 0;
    exp_40_ram[214] = 0;
    exp_40_ram[215] = 0;
    exp_40_ram[216] = 0;
    exp_40_ram[217] = 0;
    exp_40_ram[218] = 0;
    exp_40_ram[219] = 64;
    exp_40_ram[220] = 0;
    exp_40_ram[221] = 136;
    exp_40_ram[222] = 0;
    exp_40_ram[223] = 106;
    exp_40_ram[224] = 0;
    exp_40_ram[225] = 132;
    exp_40_ram[226] = 0;
    exp_40_ram[227] = 18;
    exp_40_ram[228] = 0;
    exp_40_ram[229] = 215;
    exp_40_ram[230] = 0;
    exp_40_ram[231] = 205;
    exp_40_ram[232] = 0;
    exp_40_ram[233] = 0;
    exp_40_ram[234] = 0;
    exp_40_ram[235] = 0;
    exp_40_ram[236] = 0;
    exp_40_ram[237] = 0;
    exp_40_ram[238] = 0;
    exp_40_ram[239] = 0;
    exp_40_ram[240] = 160;
    exp_40_ram[241] = 128;
    exp_40_ram[242] = 7;
    exp_40_ram[243] = 5;
    exp_40_ram[244] = 135;
    exp_40_ram[245] = 71;
    exp_40_ram[246] = 20;
    exp_40_ram[247] = 128;
    exp_40_ram[248] = 5;
    exp_40_ram[249] = 160;
    exp_40_ram[250] = 240;
    exp_40_ram[251] = 1;
    exp_40_ram[252] = 39;
    exp_40_ram[253] = 36;
    exp_40_ram[254] = 164;
    exp_40_ram[255] = 38;
    exp_40_ram[256] = 5;
    exp_40_ram[257] = 240;
    exp_40_ram[258] = 7;
    exp_40_ram[259] = 32;
    exp_40_ram[260] = 32;
    exp_40_ram[261] = 36;
    exp_40_ram[262] = 5;
    exp_40_ram[263] = 1;
    exp_40_ram[264] = 128;
    exp_40_ram[265] = 1;
    exp_40_ram[266] = 46;
    exp_40_ram[267] = 4;
    exp_40_ram[268] = 7;
    exp_40_ram[269] = 36;
    exp_40_ram[270] = 34;
    exp_40_ram[271] = 32;
    exp_40_ram[272] = 7;
    exp_40_ram[273] = 0;
    exp_40_ram[274] = 36;
    exp_40_ram[275] = 1;
    exp_40_ram[276] = 128;
    exp_40_ram[277] = 1;
    exp_40_ram[278] = 46;
    exp_40_ram[279] = 44;
    exp_40_ram[280] = 4;
    exp_40_ram[281] = 7;
    exp_40_ram[282] = 36;
    exp_40_ram[283] = 34;
    exp_40_ram[284] = 32;
    exp_40_ram[285] = 7;
    exp_40_ram[286] = 71;
    exp_40_ram[287] = 136;
    exp_40_ram[288] = 71;
    exp_40_ram[289] = 133;
    exp_40_ram[290] = 16;
    exp_40_ram[291] = 0;
    exp_40_ram[292] = 32;
    exp_40_ram[293] = 36;
    exp_40_ram[294] = 1;
    exp_40_ram[295] = 128;
    exp_40_ram[296] = 1;
    exp_40_ram[297] = 38;
    exp_40_ram[298] = 4;
    exp_40_ram[299] = 46;
    exp_40_ram[300] = 44;
    exp_40_ram[301] = 39;
    exp_40_ram[302] = 38;
    exp_40_ram[303] = 0;
    exp_40_ram[304] = 39;
    exp_40_ram[305] = 135;
    exp_40_ram[306] = 38;
    exp_40_ram[307] = 39;
    exp_40_ram[308] = 199;
    exp_40_ram[309] = 138;
    exp_40_ram[310] = 39;
    exp_40_ram[311] = 135;
    exp_40_ram[312] = 44;
    exp_40_ram[313] = 158;
    exp_40_ram[314] = 39;
    exp_40_ram[315] = 39;
    exp_40_ram[316] = 7;
    exp_40_ram[317] = 133;
    exp_40_ram[318] = 36;
    exp_40_ram[319] = 1;
    exp_40_ram[320] = 128;
    exp_40_ram[321] = 1;
    exp_40_ram[322] = 46;
    exp_40_ram[323] = 4;
    exp_40_ram[324] = 7;
    exp_40_ram[325] = 7;
    exp_40_ram[326] = 71;
    exp_40_ram[327] = 7;
    exp_40_ram[328] = 252;
    exp_40_ram[329] = 71;
    exp_40_ram[330] = 7;
    exp_40_ram[331] = 230;
    exp_40_ram[332] = 7;
    exp_40_ram[333] = 0;
    exp_40_ram[334] = 7;
    exp_40_ram[335] = 247;
    exp_40_ram[336] = 247;
    exp_40_ram[337] = 133;
    exp_40_ram[338] = 36;
    exp_40_ram[339] = 1;
    exp_40_ram[340] = 128;
    exp_40_ram[341] = 1;
    exp_40_ram[342] = 38;
    exp_40_ram[343] = 36;
    exp_40_ram[344] = 4;
    exp_40_ram[345] = 46;
    exp_40_ram[346] = 38;
    exp_40_ram[347] = 0;
    exp_40_ram[348] = 39;
    exp_40_ram[349] = 7;
    exp_40_ram[350] = 151;
    exp_40_ram[351] = 135;
    exp_40_ram[352] = 151;
    exp_40_ram[353] = 134;
    exp_40_ram[354] = 39;
    exp_40_ram[355] = 167;
    exp_40_ram[356] = 134;
    exp_40_ram[357] = 39;
    exp_40_ram[358] = 32;
    exp_40_ram[359] = 199;
    exp_40_ram[360] = 7;
    exp_40_ram[361] = 135;
    exp_40_ram[362] = 38;
    exp_40_ram[363] = 39;
    exp_40_ram[364] = 167;
    exp_40_ram[365] = 199;
    exp_40_ram[366] = 133;
    exp_40_ram[367] = 240;
    exp_40_ram[368] = 7;
    exp_40_ram[369] = 150;
    exp_40_ram[370] = 39;
    exp_40_ram[371] = 133;
    exp_40_ram[372] = 32;
    exp_40_ram[373] = 36;
    exp_40_ram[374] = 1;
    exp_40_ram[375] = 128;
    exp_40_ram[376] = 1;
    exp_40_ram[377] = 46;
    exp_40_ram[378] = 44;
    exp_40_ram[379] = 4;
    exp_40_ram[380] = 46;
    exp_40_ram[381] = 44;
    exp_40_ram[382] = 42;
    exp_40_ram[383] = 40;
    exp_40_ram[384] = 38;
    exp_40_ram[385] = 36;
    exp_40_ram[386] = 34;
    exp_40_ram[387] = 32;
    exp_40_ram[388] = 39;
    exp_40_ram[389] = 36;
    exp_40_ram[390] = 39;
    exp_40_ram[391] = 247;
    exp_40_ram[392] = 156;
    exp_40_ram[393] = 39;
    exp_40_ram[394] = 247;
    exp_40_ram[395] = 150;
    exp_40_ram[396] = 39;
    exp_40_ram[397] = 38;
    exp_40_ram[398] = 0;
    exp_40_ram[399] = 39;
    exp_40_ram[400] = 135;
    exp_40_ram[401] = 42;
    exp_40_ram[402] = 39;
    exp_40_ram[403] = 38;
    exp_40_ram[404] = 134;
    exp_40_ram[405] = 37;
    exp_40_ram[406] = 5;
    exp_40_ram[407] = 0;
    exp_40_ram[408] = 39;
    exp_40_ram[409] = 135;
    exp_40_ram[410] = 38;
    exp_40_ram[411] = 39;
    exp_40_ram[412] = 39;
    exp_40_ram[413] = 100;
    exp_40_ram[414] = 0;
    exp_40_ram[415] = 39;
    exp_40_ram[416] = 135;
    exp_40_ram[417] = 36;
    exp_40_ram[418] = 39;
    exp_40_ram[419] = 39;
    exp_40_ram[420] = 7;
    exp_40_ram[421] = 197;
    exp_40_ram[422] = 39;
    exp_40_ram[423] = 135;
    exp_40_ram[424] = 42;
    exp_40_ram[425] = 39;
    exp_40_ram[426] = 38;
    exp_40_ram[427] = 134;
    exp_40_ram[428] = 37;
    exp_40_ram[429] = 0;
    exp_40_ram[430] = 39;
    exp_40_ram[431] = 144;
    exp_40_ram[432] = 39;
    exp_40_ram[433] = 247;
    exp_40_ram[434] = 128;
    exp_40_ram[435] = 0;
    exp_40_ram[436] = 39;
    exp_40_ram[437] = 135;
    exp_40_ram[438] = 42;
    exp_40_ram[439] = 39;
    exp_40_ram[440] = 38;
    exp_40_ram[441] = 134;
    exp_40_ram[442] = 37;
    exp_40_ram[443] = 5;
    exp_40_ram[444] = 0;
    exp_40_ram[445] = 39;
    exp_40_ram[446] = 39;
    exp_40_ram[447] = 7;
    exp_40_ram[448] = 39;
    exp_40_ram[449] = 230;
    exp_40_ram[450] = 39;
    exp_40_ram[451] = 133;
    exp_40_ram[452] = 32;
    exp_40_ram[453] = 36;
    exp_40_ram[454] = 1;
    exp_40_ram[455] = 128;
    exp_40_ram[456] = 1;
    exp_40_ram[457] = 38;
    exp_40_ram[458] = 36;
    exp_40_ram[459] = 4;
    exp_40_ram[460] = 38;
    exp_40_ram[461] = 36;
    exp_40_ram[462] = 34;
    exp_40_ram[463] = 32;
    exp_40_ram[464] = 46;
    exp_40_ram[465] = 44;
    exp_40_ram[466] = 7;
    exp_40_ram[467] = 40;
    exp_40_ram[468] = 11;
    exp_40_ram[469] = 39;
    exp_40_ram[470] = 247;
    exp_40_ram[471] = 154;
    exp_40_ram[472] = 39;
    exp_40_ram[473] = 136;
    exp_40_ram[474] = 39;
    exp_40_ram[475] = 247;
    exp_40_ram[476] = 130;
    exp_40_ram[477] = 71;
    exp_40_ram[478] = 152;
    exp_40_ram[479] = 39;
    exp_40_ram[480] = 247;
    exp_40_ram[481] = 136;
    exp_40_ram[482] = 39;
    exp_40_ram[483] = 135;
    exp_40_ram[484] = 34;
    exp_40_ram[485] = 0;
    exp_40_ram[486] = 39;
    exp_40_ram[487] = 135;
    exp_40_ram[488] = 44;
    exp_40_ram[489] = 39;
    exp_40_ram[490] = 7;
    exp_40_ram[491] = 7;
    exp_40_ram[492] = 128;
    exp_40_ram[493] = 39;
    exp_40_ram[494] = 39;
    exp_40_ram[495] = 120;
    exp_40_ram[496] = 39;
    exp_40_ram[497] = 7;
    exp_40_ram[498] = 248;
    exp_40_ram[499] = 0;
    exp_40_ram[500] = 39;
    exp_40_ram[501] = 135;
    exp_40_ram[502] = 44;
    exp_40_ram[503] = 39;
    exp_40_ram[504] = 7;
    exp_40_ram[505] = 7;
    exp_40_ram[506] = 128;
    exp_40_ram[507] = 39;
    exp_40_ram[508] = 247;
    exp_40_ram[509] = 142;
    exp_40_ram[510] = 39;
    exp_40_ram[511] = 39;
    exp_40_ram[512] = 120;
    exp_40_ram[513] = 39;
    exp_40_ram[514] = 7;
    exp_40_ram[515] = 242;
    exp_40_ram[516] = 39;
    exp_40_ram[517] = 247;
    exp_40_ram[518] = 128;
    exp_40_ram[519] = 39;
    exp_40_ram[520] = 247;
    exp_40_ram[521] = 152;
    exp_40_ram[522] = 39;
    exp_40_ram[523] = 132;
    exp_40_ram[524] = 39;
    exp_40_ram[525] = 39;
    exp_40_ram[526] = 8;
    exp_40_ram[527] = 39;
    exp_40_ram[528] = 39;
    exp_40_ram[529] = 24;
    exp_40_ram[530] = 39;
    exp_40_ram[531] = 135;
    exp_40_ram[532] = 44;
    exp_40_ram[533] = 39;
    exp_40_ram[534] = 142;
    exp_40_ram[535] = 39;
    exp_40_ram[536] = 7;
    exp_40_ram[537] = 24;
    exp_40_ram[538] = 39;
    exp_40_ram[539] = 135;
    exp_40_ram[540] = 44;
    exp_40_ram[541] = 39;
    exp_40_ram[542] = 7;
    exp_40_ram[543] = 30;
    exp_40_ram[544] = 39;
    exp_40_ram[545] = 247;
    exp_40_ram[546] = 152;
    exp_40_ram[547] = 39;
    exp_40_ram[548] = 7;
    exp_40_ram[549] = 226;
    exp_40_ram[550] = 39;
    exp_40_ram[551] = 135;
    exp_40_ram[552] = 44;
    exp_40_ram[553] = 39;
    exp_40_ram[554] = 7;
    exp_40_ram[555] = 7;
    exp_40_ram[556] = 128;
    exp_40_ram[557] = 0;
    exp_40_ram[558] = 39;
    exp_40_ram[559] = 7;
    exp_40_ram[560] = 30;
    exp_40_ram[561] = 39;
    exp_40_ram[562] = 247;
    exp_40_ram[563] = 136;
    exp_40_ram[564] = 39;
    exp_40_ram[565] = 7;
    exp_40_ram[566] = 226;
    exp_40_ram[567] = 39;
    exp_40_ram[568] = 135;
    exp_40_ram[569] = 44;
    exp_40_ram[570] = 39;
    exp_40_ram[571] = 7;
    exp_40_ram[572] = 7;
    exp_40_ram[573] = 128;
    exp_40_ram[574] = 0;
    exp_40_ram[575] = 39;
    exp_40_ram[576] = 7;
    exp_40_ram[577] = 22;
    exp_40_ram[578] = 39;
    exp_40_ram[579] = 7;
    exp_40_ram[580] = 224;
    exp_40_ram[581] = 39;
    exp_40_ram[582] = 135;
    exp_40_ram[583] = 44;
    exp_40_ram[584] = 39;
    exp_40_ram[585] = 7;
    exp_40_ram[586] = 7;
    exp_40_ram[587] = 128;
    exp_40_ram[588] = 39;
    exp_40_ram[589] = 7;
    exp_40_ram[590] = 224;
    exp_40_ram[591] = 39;
    exp_40_ram[592] = 135;
    exp_40_ram[593] = 44;
    exp_40_ram[594] = 39;
    exp_40_ram[595] = 7;
    exp_40_ram[596] = 7;
    exp_40_ram[597] = 128;
    exp_40_ram[598] = 39;
    exp_40_ram[599] = 7;
    exp_40_ram[600] = 224;
    exp_40_ram[601] = 71;
    exp_40_ram[602] = 130;
    exp_40_ram[603] = 39;
    exp_40_ram[604] = 135;
    exp_40_ram[605] = 44;
    exp_40_ram[606] = 39;
    exp_40_ram[607] = 7;
    exp_40_ram[608] = 7;
    exp_40_ram[609] = 128;
    exp_40_ram[610] = 0;
    exp_40_ram[611] = 39;
    exp_40_ram[612] = 247;
    exp_40_ram[613] = 130;
    exp_40_ram[614] = 39;
    exp_40_ram[615] = 135;
    exp_40_ram[616] = 44;
    exp_40_ram[617] = 39;
    exp_40_ram[618] = 7;
    exp_40_ram[619] = 7;
    exp_40_ram[620] = 128;
    exp_40_ram[621] = 0;
    exp_40_ram[622] = 39;
    exp_40_ram[623] = 247;
    exp_40_ram[624] = 128;
    exp_40_ram[625] = 39;
    exp_40_ram[626] = 135;
    exp_40_ram[627] = 44;
    exp_40_ram[628] = 39;
    exp_40_ram[629] = 7;
    exp_40_ram[630] = 7;
    exp_40_ram[631] = 128;
    exp_40_ram[632] = 40;
    exp_40_ram[633] = 40;
    exp_40_ram[634] = 39;
    exp_40_ram[635] = 39;
    exp_40_ram[636] = 38;
    exp_40_ram[637] = 38;
    exp_40_ram[638] = 37;
    exp_40_ram[639] = 37;
    exp_40_ram[640] = 240;
    exp_40_ram[641] = 7;
    exp_40_ram[642] = 133;
    exp_40_ram[643] = 32;
    exp_40_ram[644] = 36;
    exp_40_ram[645] = 1;
    exp_40_ram[646] = 128;
    exp_40_ram[647] = 1;
    exp_40_ram[648] = 38;
    exp_40_ram[649] = 36;
    exp_40_ram[650] = 4;
    exp_40_ram[651] = 46;
    exp_40_ram[652] = 44;
    exp_40_ram[653] = 42;
    exp_40_ram[654] = 40;
    exp_40_ram[655] = 38;
    exp_40_ram[656] = 34;
    exp_40_ram[657] = 32;
    exp_40_ram[658] = 5;
    exp_40_ram[659] = 38;
    exp_40_ram[660] = 39;
    exp_40_ram[661] = 152;
    exp_40_ram[662] = 39;
    exp_40_ram[663] = 247;
    exp_40_ram[664] = 34;
    exp_40_ram[665] = 39;
    exp_40_ram[666] = 247;
    exp_40_ram[667] = 134;
    exp_40_ram[668] = 39;
    exp_40_ram[669] = 140;
    exp_40_ram[670] = 39;
    exp_40_ram[671] = 39;
    exp_40_ram[672] = 119;
    exp_40_ram[673] = 5;
    exp_40_ram[674] = 71;
    exp_40_ram[675] = 7;
    exp_40_ram[676] = 234;
    exp_40_ram[677] = 71;
    exp_40_ram[678] = 135;
    exp_40_ram[679] = 247;
    exp_40_ram[680] = 0;
    exp_40_ram[681] = 39;
    exp_40_ram[682] = 247;
    exp_40_ram[683] = 134;
    exp_40_ram[684] = 7;
    exp_40_ram[685] = 0;
    exp_40_ram[686] = 7;
    exp_40_ram[687] = 71;
    exp_40_ram[688] = 135;
    exp_40_ram[689] = 247;
    exp_40_ram[690] = 135;
    exp_40_ram[691] = 247;
    exp_40_ram[692] = 39;
    exp_40_ram[693] = 6;
    exp_40_ram[694] = 38;
    exp_40_ram[695] = 6;
    exp_40_ram[696] = 135;
    exp_40_ram[697] = 12;
    exp_40_ram[698] = 39;
    exp_40_ram[699] = 39;
    exp_40_ram[700] = 87;
    exp_40_ram[701] = 38;
    exp_40_ram[702] = 39;
    exp_40_ram[703] = 136;
    exp_40_ram[704] = 39;
    exp_40_ram[705] = 7;
    exp_40_ram[706] = 248;
    exp_40_ram[707] = 70;
    exp_40_ram[708] = 7;
    exp_40_ram[709] = 39;
    exp_40_ram[710] = 36;
    exp_40_ram[711] = 39;
    exp_40_ram[712] = 34;
    exp_40_ram[713] = 39;
    exp_40_ram[714] = 32;
    exp_40_ram[715] = 40;
    exp_40_ram[716] = 136;
    exp_40_ram[717] = 39;
    exp_40_ram[718] = 38;
    exp_40_ram[719] = 38;
    exp_40_ram[720] = 37;
    exp_40_ram[721] = 37;
    exp_40_ram[722] = 240;
    exp_40_ram[723] = 7;
    exp_40_ram[724] = 133;
    exp_40_ram[725] = 32;
    exp_40_ram[726] = 36;
    exp_40_ram[727] = 1;
    exp_40_ram[728] = 128;
    exp_40_ram[729] = 1;
    exp_40_ram[730] = 46;
    exp_40_ram[731] = 44;
    exp_40_ram[732] = 4;
    exp_40_ram[733] = 38;
    exp_40_ram[734] = 36;
    exp_40_ram[735] = 34;
    exp_40_ram[736] = 32;
    exp_40_ram[737] = 46;
    exp_40_ram[738] = 46;
    exp_40_ram[739] = 39;
    exp_40_ram[740] = 156;
    exp_40_ram[741] = 7;
    exp_40_ram[742] = 38;
    exp_40_ram[743] = 0;
    exp_40_ram[744] = 39;
    exp_40_ram[745] = 199;
    exp_40_ram[746] = 7;
    exp_40_ram[747] = 14;
    exp_40_ram[748] = 39;
    exp_40_ram[749] = 197;
    exp_40_ram[750] = 39;
    exp_40_ram[751] = 135;
    exp_40_ram[752] = 46;
    exp_40_ram[753] = 39;
    exp_40_ram[754] = 38;
    exp_40_ram[755] = 134;
    exp_40_ram[756] = 37;
    exp_40_ram[757] = 0;
    exp_40_ram[758] = 39;
    exp_40_ram[759] = 135;
    exp_40_ram[760] = 32;
    exp_40_ram[761] = 0;
    exp_40_ram[762] = 39;
    exp_40_ram[763] = 135;
    exp_40_ram[764] = 32;
    exp_40_ram[765] = 38;
    exp_40_ram[766] = 39;
    exp_40_ram[767] = 199;
    exp_40_ram[768] = 135;
    exp_40_ram[769] = 7;
    exp_40_ram[770] = 104;
    exp_40_ram[771] = 151;
    exp_40_ram[772] = 39;
    exp_40_ram[773] = 135;
    exp_40_ram[774] = 7;
    exp_40_ram[775] = 167;
    exp_40_ram[776] = 128;
    exp_40_ram[777] = 39;
    exp_40_ram[778] = 231;
    exp_40_ram[779] = 38;
    exp_40_ram[780] = 39;
    exp_40_ram[781] = 135;
    exp_40_ram[782] = 32;
    exp_40_ram[783] = 7;
    exp_40_ram[784] = 32;
    exp_40_ram[785] = 0;
    exp_40_ram[786] = 39;
    exp_40_ram[787] = 231;
    exp_40_ram[788] = 38;
    exp_40_ram[789] = 39;
    exp_40_ram[790] = 135;
    exp_40_ram[791] = 32;
    exp_40_ram[792] = 7;
    exp_40_ram[793] = 32;
    exp_40_ram[794] = 0;
    exp_40_ram[795] = 39;
    exp_40_ram[796] = 231;
    exp_40_ram[797] = 38;
    exp_40_ram[798] = 39;
    exp_40_ram[799] = 135;
    exp_40_ram[800] = 32;
    exp_40_ram[801] = 7;
    exp_40_ram[802] = 32;
    exp_40_ram[803] = 0;
    exp_40_ram[804] = 39;
    exp_40_ram[805] = 231;
    exp_40_ram[806] = 38;
    exp_40_ram[807] = 39;
    exp_40_ram[808] = 135;
    exp_40_ram[809] = 32;
    exp_40_ram[810] = 7;
    exp_40_ram[811] = 32;
    exp_40_ram[812] = 0;
    exp_40_ram[813] = 39;
    exp_40_ram[814] = 231;
    exp_40_ram[815] = 38;
    exp_40_ram[816] = 39;
    exp_40_ram[817] = 135;
    exp_40_ram[818] = 32;
    exp_40_ram[819] = 7;
    exp_40_ram[820] = 32;
    exp_40_ram[821] = 0;
    exp_40_ram[822] = 32;
    exp_40_ram[823] = 0;
    exp_40_ram[824] = 39;
    exp_40_ram[825] = 154;
    exp_40_ram[826] = 36;
    exp_40_ram[827] = 39;
    exp_40_ram[828] = 199;
    exp_40_ram[829] = 133;
    exp_40_ram[830] = 240;
    exp_40_ram[831] = 7;
    exp_40_ram[832] = 140;
    exp_40_ram[833] = 7;
    exp_40_ram[834] = 133;
    exp_40_ram[835] = 240;
    exp_40_ram[836] = 36;
    exp_40_ram[837] = 0;
    exp_40_ram[838] = 39;
    exp_40_ram[839] = 199;
    exp_40_ram[840] = 7;
    exp_40_ram[841] = 24;
    exp_40_ram[842] = 39;
    exp_40_ram[843] = 135;
    exp_40_ram[844] = 46;
    exp_40_ram[845] = 167;
    exp_40_ram[846] = 36;
    exp_40_ram[847] = 39;
    exp_40_ram[848] = 208;
    exp_40_ram[849] = 39;
    exp_40_ram[850] = 231;
    exp_40_ram[851] = 38;
    exp_40_ram[852] = 39;
    exp_40_ram[853] = 7;
    exp_40_ram[854] = 36;
    exp_40_ram[855] = 0;
    exp_40_ram[856] = 39;
    exp_40_ram[857] = 36;
    exp_40_ram[858] = 39;
    exp_40_ram[859] = 135;
    exp_40_ram[860] = 32;
    exp_40_ram[861] = 34;
    exp_40_ram[862] = 39;
    exp_40_ram[863] = 199;
    exp_40_ram[864] = 7;
    exp_40_ram[865] = 20;
    exp_40_ram[866] = 39;
    exp_40_ram[867] = 231;
    exp_40_ram[868] = 38;
    exp_40_ram[869] = 39;
    exp_40_ram[870] = 135;
    exp_40_ram[871] = 32;
    exp_40_ram[872] = 39;
    exp_40_ram[873] = 199;
    exp_40_ram[874] = 133;
    exp_40_ram[875] = 240;
    exp_40_ram[876] = 7;
    exp_40_ram[877] = 140;
    exp_40_ram[878] = 7;
    exp_40_ram[879] = 133;
    exp_40_ram[880] = 240;
    exp_40_ram[881] = 34;
    exp_40_ram[882] = 0;
    exp_40_ram[883] = 39;
    exp_40_ram[884] = 199;
    exp_40_ram[885] = 7;
    exp_40_ram[886] = 26;
    exp_40_ram[887] = 39;
    exp_40_ram[888] = 135;
    exp_40_ram[889] = 46;
    exp_40_ram[890] = 167;
    exp_40_ram[891] = 34;
    exp_40_ram[892] = 39;
    exp_40_ram[893] = 212;
    exp_40_ram[894] = 7;
    exp_40_ram[895] = 34;
    exp_40_ram[896] = 39;
    exp_40_ram[897] = 135;
    exp_40_ram[898] = 32;
    exp_40_ram[899] = 39;
    exp_40_ram[900] = 199;
    exp_40_ram[901] = 135;
    exp_40_ram[902] = 7;
    exp_40_ram[903] = 108;
    exp_40_ram[904] = 151;
    exp_40_ram[905] = 39;
    exp_40_ram[906] = 135;
    exp_40_ram[907] = 7;
    exp_40_ram[908] = 167;
    exp_40_ram[909] = 128;
    exp_40_ram[910] = 39;
    exp_40_ram[911] = 231;
    exp_40_ram[912] = 38;
    exp_40_ram[913] = 39;
    exp_40_ram[914] = 135;
    exp_40_ram[915] = 32;
    exp_40_ram[916] = 39;
    exp_40_ram[917] = 199;
    exp_40_ram[918] = 7;
    exp_40_ram[919] = 16;
    exp_40_ram[920] = 39;
    exp_40_ram[921] = 231;
    exp_40_ram[922] = 38;
    exp_40_ram[923] = 39;
    exp_40_ram[924] = 135;
    exp_40_ram[925] = 32;
    exp_40_ram[926] = 0;
    exp_40_ram[927] = 39;
    exp_40_ram[928] = 231;
    exp_40_ram[929] = 38;
    exp_40_ram[930] = 39;
    exp_40_ram[931] = 135;
    exp_40_ram[932] = 32;
    exp_40_ram[933] = 39;
    exp_40_ram[934] = 199;
    exp_40_ram[935] = 7;
    exp_40_ram[936] = 18;
    exp_40_ram[937] = 39;
    exp_40_ram[938] = 231;
    exp_40_ram[939] = 38;
    exp_40_ram[940] = 39;
    exp_40_ram[941] = 135;
    exp_40_ram[942] = 32;
    exp_40_ram[943] = 0;
    exp_40_ram[944] = 39;
    exp_40_ram[945] = 231;
    exp_40_ram[946] = 38;
    exp_40_ram[947] = 39;
    exp_40_ram[948] = 135;
    exp_40_ram[949] = 32;
    exp_40_ram[950] = 0;
    exp_40_ram[951] = 39;
    exp_40_ram[952] = 231;
    exp_40_ram[953] = 38;
    exp_40_ram[954] = 39;
    exp_40_ram[955] = 135;
    exp_40_ram[956] = 32;
    exp_40_ram[957] = 0;
    exp_40_ram[958] = 39;
    exp_40_ram[959] = 231;
    exp_40_ram[960] = 38;
    exp_40_ram[961] = 39;
    exp_40_ram[962] = 135;
    exp_40_ram[963] = 32;
    exp_40_ram[964] = 0;
    exp_40_ram[965] = 0;
    exp_40_ram[966] = 0;
    exp_40_ram[967] = 0;
    exp_40_ram[968] = 0;
    exp_40_ram[969] = 0;
    exp_40_ram[970] = 39;
    exp_40_ram[971] = 199;
    exp_40_ram[972] = 135;
    exp_40_ram[973] = 7;
    exp_40_ram[974] = 108;
    exp_40_ram[975] = 151;
    exp_40_ram[976] = 39;
    exp_40_ram[977] = 135;
    exp_40_ram[978] = 7;
    exp_40_ram[979] = 167;
    exp_40_ram[980] = 128;
    exp_40_ram[981] = 39;
    exp_40_ram[982] = 199;
    exp_40_ram[983] = 7;
    exp_40_ram[984] = 10;
    exp_40_ram[985] = 39;
    exp_40_ram[986] = 199;
    exp_40_ram[987] = 7;
    exp_40_ram[988] = 24;
    exp_40_ram[989] = 7;
    exp_40_ram[990] = 44;
    exp_40_ram[991] = 0;
    exp_40_ram[992] = 39;
    exp_40_ram[993] = 199;
    exp_40_ram[994] = 7;
    exp_40_ram[995] = 24;
    exp_40_ram[996] = 7;
    exp_40_ram[997] = 44;
    exp_40_ram[998] = 0;
    exp_40_ram[999] = 39;
    exp_40_ram[1000] = 199;
    exp_40_ram[1001] = 7;
    exp_40_ram[1002] = 24;
    exp_40_ram[1003] = 7;
    exp_40_ram[1004] = 44;
    exp_40_ram[1005] = 0;
    exp_40_ram[1006] = 7;
    exp_40_ram[1007] = 44;
    exp_40_ram[1008] = 39;
    exp_40_ram[1009] = 247;
    exp_40_ram[1010] = 38;
    exp_40_ram[1011] = 39;
    exp_40_ram[1012] = 199;
    exp_40_ram[1013] = 7;
    exp_40_ram[1014] = 24;
    exp_40_ram[1015] = 39;
    exp_40_ram[1016] = 231;
    exp_40_ram[1017] = 38;
    exp_40_ram[1018] = 39;
    exp_40_ram[1019] = 199;
    exp_40_ram[1020] = 7;
    exp_40_ram[1021] = 0;
    exp_40_ram[1022] = 39;
    exp_40_ram[1023] = 199;
    exp_40_ram[1024] = 7;
    exp_40_ram[1025] = 8;
    exp_40_ram[1026] = 39;
    exp_40_ram[1027] = 247;
    exp_40_ram[1028] = 38;
    exp_40_ram[1029] = 39;
    exp_40_ram[1030] = 247;
    exp_40_ram[1031] = 136;
    exp_40_ram[1032] = 39;
    exp_40_ram[1033] = 247;
    exp_40_ram[1034] = 38;
    exp_40_ram[1035] = 39;
    exp_40_ram[1036] = 199;
    exp_40_ram[1037] = 7;
    exp_40_ram[1038] = 10;
    exp_40_ram[1039] = 39;
    exp_40_ram[1040] = 199;
    exp_40_ram[1041] = 7;
    exp_40_ram[1042] = 24;
    exp_40_ram[1043] = 39;
    exp_40_ram[1044] = 247;
    exp_40_ram[1045] = 158;
    exp_40_ram[1046] = 39;
    exp_40_ram[1047] = 247;
    exp_40_ram[1048] = 140;
    exp_40_ram[1049] = 39;
    exp_40_ram[1050] = 135;
    exp_40_ram[1051] = 46;
    exp_40_ram[1052] = 167;
    exp_40_ram[1053] = 44;
    exp_40_ram[1054] = 39;
    exp_40_ram[1055] = 215;
    exp_40_ram[1056] = 39;
    exp_40_ram[1057] = 71;
    exp_40_ram[1058] = 135;
    exp_40_ram[1059] = 134;
    exp_40_ram[1060] = 39;
    exp_40_ram[1061] = 215;
    exp_40_ram[1062] = 247;
    exp_40_ram[1063] = 39;
    exp_40_ram[1064] = 34;
    exp_40_ram[1065] = 39;
    exp_40_ram[1066] = 32;
    exp_40_ram[1067] = 40;
    exp_40_ram[1068] = 40;
    exp_40_ram[1069] = 7;
    exp_40_ram[1070] = 135;
    exp_40_ram[1071] = 38;
    exp_40_ram[1072] = 38;
    exp_40_ram[1073] = 37;
    exp_40_ram[1074] = 37;
    exp_40_ram[1075] = 240;
    exp_40_ram[1076] = 46;
    exp_40_ram[1077] = 0;
    exp_40_ram[1078] = 39;
    exp_40_ram[1079] = 247;
    exp_40_ram[1080] = 142;
    exp_40_ram[1081] = 39;
    exp_40_ram[1082] = 135;
    exp_40_ram[1083] = 46;
    exp_40_ram[1084] = 167;
    exp_40_ram[1085] = 247;
    exp_40_ram[1086] = 0;
    exp_40_ram[1087] = 39;
    exp_40_ram[1088] = 247;
    exp_40_ram[1089] = 128;
    exp_40_ram[1090] = 39;
    exp_40_ram[1091] = 135;
    exp_40_ram[1092] = 46;
    exp_40_ram[1093] = 167;
    exp_40_ram[1094] = 151;
    exp_40_ram[1095] = 215;
    exp_40_ram[1096] = 0;
    exp_40_ram[1097] = 39;
    exp_40_ram[1098] = 135;
    exp_40_ram[1099] = 46;
    exp_40_ram[1100] = 167;
    exp_40_ram[1101] = 46;
    exp_40_ram[1102] = 39;
    exp_40_ram[1103] = 215;
    exp_40_ram[1104] = 39;
    exp_40_ram[1105] = 71;
    exp_40_ram[1106] = 135;
    exp_40_ram[1107] = 134;
    exp_40_ram[1108] = 39;
    exp_40_ram[1109] = 215;
    exp_40_ram[1110] = 247;
    exp_40_ram[1111] = 39;
    exp_40_ram[1112] = 34;
    exp_40_ram[1113] = 39;
    exp_40_ram[1114] = 32;
    exp_40_ram[1115] = 40;
    exp_40_ram[1116] = 40;
    exp_40_ram[1117] = 7;
    exp_40_ram[1118] = 135;
    exp_40_ram[1119] = 38;
    exp_40_ram[1120] = 38;
    exp_40_ram[1121] = 37;
    exp_40_ram[1122] = 37;
    exp_40_ram[1123] = 240;
    exp_40_ram[1124] = 46;
    exp_40_ram[1125] = 0;
    exp_40_ram[1126] = 39;
    exp_40_ram[1127] = 247;
    exp_40_ram[1128] = 152;
    exp_40_ram[1129] = 39;
    exp_40_ram[1130] = 247;
    exp_40_ram[1131] = 134;
    exp_40_ram[1132] = 39;
    exp_40_ram[1133] = 135;
    exp_40_ram[1134] = 46;
    exp_40_ram[1135] = 167;
    exp_40_ram[1136] = 39;
    exp_40_ram[1137] = 34;
    exp_40_ram[1138] = 39;
    exp_40_ram[1139] = 32;
    exp_40_ram[1140] = 40;
    exp_40_ram[1141] = 40;
    exp_40_ram[1142] = 7;
    exp_40_ram[1143] = 38;
    exp_40_ram[1144] = 38;
    exp_40_ram[1145] = 37;
    exp_40_ram[1146] = 37;
    exp_40_ram[1147] = 240;
    exp_40_ram[1148] = 46;
    exp_40_ram[1149] = 0;
    exp_40_ram[1150] = 39;
    exp_40_ram[1151] = 247;
    exp_40_ram[1152] = 142;
    exp_40_ram[1153] = 39;
    exp_40_ram[1154] = 135;
    exp_40_ram[1155] = 46;
    exp_40_ram[1156] = 167;
    exp_40_ram[1157] = 247;
    exp_40_ram[1158] = 0;
    exp_40_ram[1159] = 39;
    exp_40_ram[1160] = 247;
    exp_40_ram[1161] = 128;
    exp_40_ram[1162] = 39;
    exp_40_ram[1163] = 135;
    exp_40_ram[1164] = 46;
    exp_40_ram[1165] = 167;
    exp_40_ram[1166] = 151;
    exp_40_ram[1167] = 215;
    exp_40_ram[1168] = 0;
    exp_40_ram[1169] = 39;
    exp_40_ram[1170] = 135;
    exp_40_ram[1171] = 46;
    exp_40_ram[1172] = 167;
    exp_40_ram[1173] = 32;
    exp_40_ram[1174] = 39;
    exp_40_ram[1175] = 34;
    exp_40_ram[1176] = 39;
    exp_40_ram[1177] = 32;
    exp_40_ram[1178] = 40;
    exp_40_ram[1179] = 40;
    exp_40_ram[1180] = 7;
    exp_40_ram[1181] = 39;
    exp_40_ram[1182] = 38;
    exp_40_ram[1183] = 38;
    exp_40_ram[1184] = 37;
    exp_40_ram[1185] = 37;
    exp_40_ram[1186] = 240;
    exp_40_ram[1187] = 46;
    exp_40_ram[1188] = 39;
    exp_40_ram[1189] = 135;
    exp_40_ram[1190] = 32;
    exp_40_ram[1191] = 0;
    exp_40_ram[1192] = 7;
    exp_40_ram[1193] = 42;
    exp_40_ram[1194] = 39;
    exp_40_ram[1195] = 247;
    exp_40_ram[1196] = 144;
    exp_40_ram[1197] = 0;
    exp_40_ram[1198] = 39;
    exp_40_ram[1199] = 135;
    exp_40_ram[1200] = 46;
    exp_40_ram[1201] = 39;
    exp_40_ram[1202] = 38;
    exp_40_ram[1203] = 134;
    exp_40_ram[1204] = 37;
    exp_40_ram[1205] = 5;
    exp_40_ram[1206] = 0;
    exp_40_ram[1207] = 39;
    exp_40_ram[1208] = 135;
    exp_40_ram[1209] = 42;
    exp_40_ram[1210] = 39;
    exp_40_ram[1211] = 230;
    exp_40_ram[1212] = 39;
    exp_40_ram[1213] = 135;
    exp_40_ram[1214] = 46;
    exp_40_ram[1215] = 167;
    exp_40_ram[1216] = 245;
    exp_40_ram[1217] = 39;
    exp_40_ram[1218] = 135;
    exp_40_ram[1219] = 46;
    exp_40_ram[1220] = 39;
    exp_40_ram[1221] = 38;
    exp_40_ram[1222] = 134;
    exp_40_ram[1223] = 37;
    exp_40_ram[1224] = 0;
    exp_40_ram[1225] = 39;
    exp_40_ram[1226] = 247;
    exp_40_ram[1227] = 128;
    exp_40_ram[1228] = 0;
    exp_40_ram[1229] = 39;
    exp_40_ram[1230] = 135;
    exp_40_ram[1231] = 46;
    exp_40_ram[1232] = 39;
    exp_40_ram[1233] = 38;
    exp_40_ram[1234] = 134;
    exp_40_ram[1235] = 37;
    exp_40_ram[1236] = 5;
    exp_40_ram[1237] = 0;
    exp_40_ram[1238] = 39;
    exp_40_ram[1239] = 135;
    exp_40_ram[1240] = 42;
    exp_40_ram[1241] = 39;
    exp_40_ram[1242] = 230;
    exp_40_ram[1243] = 39;
    exp_40_ram[1244] = 135;
    exp_40_ram[1245] = 32;
    exp_40_ram[1246] = 0;
    exp_40_ram[1247] = 39;
    exp_40_ram[1248] = 135;
    exp_40_ram[1249] = 46;
    exp_40_ram[1250] = 167;
    exp_40_ram[1251] = 40;
    exp_40_ram[1252] = 39;
    exp_40_ram[1253] = 134;
    exp_40_ram[1254] = 39;
    exp_40_ram[1255] = 0;
    exp_40_ram[1256] = 7;
    exp_40_ram[1257] = 133;
    exp_40_ram[1258] = 37;
    exp_40_ram[1259] = 240;
    exp_40_ram[1260] = 38;
    exp_40_ram[1261] = 39;
    exp_40_ram[1262] = 247;
    exp_40_ram[1263] = 140;
    exp_40_ram[1264] = 39;
    exp_40_ram[1265] = 39;
    exp_40_ram[1266] = 116;
    exp_40_ram[1267] = 7;
    exp_40_ram[1268] = 38;
    exp_40_ram[1269] = 39;
    exp_40_ram[1270] = 247;
    exp_40_ram[1271] = 154;
    exp_40_ram[1272] = 0;
    exp_40_ram[1273] = 39;
    exp_40_ram[1274] = 135;
    exp_40_ram[1275] = 46;
    exp_40_ram[1276] = 39;
    exp_40_ram[1277] = 38;
    exp_40_ram[1278] = 134;
    exp_40_ram[1279] = 37;
    exp_40_ram[1280] = 5;
    exp_40_ram[1281] = 0;
    exp_40_ram[1282] = 39;
    exp_40_ram[1283] = 135;
    exp_40_ram[1284] = 38;
    exp_40_ram[1285] = 39;
    exp_40_ram[1286] = 230;
    exp_40_ram[1287] = 0;
    exp_40_ram[1288] = 39;
    exp_40_ram[1289] = 135;
    exp_40_ram[1290] = 40;
    exp_40_ram[1291] = 197;
    exp_40_ram[1292] = 39;
    exp_40_ram[1293] = 135;
    exp_40_ram[1294] = 46;
    exp_40_ram[1295] = 39;
    exp_40_ram[1296] = 38;
    exp_40_ram[1297] = 134;
    exp_40_ram[1298] = 37;
    exp_40_ram[1299] = 0;
    exp_40_ram[1300] = 39;
    exp_40_ram[1301] = 199;
    exp_40_ram[1302] = 128;
    exp_40_ram[1303] = 39;
    exp_40_ram[1304] = 247;
    exp_40_ram[1305] = 142;
    exp_40_ram[1306] = 39;
    exp_40_ram[1307] = 135;
    exp_40_ram[1308] = 34;
    exp_40_ram[1309] = 150;
    exp_40_ram[1310] = 39;
    exp_40_ram[1311] = 247;
    exp_40_ram[1312] = 128;
    exp_40_ram[1313] = 0;
    exp_40_ram[1314] = 39;
    exp_40_ram[1315] = 135;
    exp_40_ram[1316] = 46;
    exp_40_ram[1317] = 39;
    exp_40_ram[1318] = 38;
    exp_40_ram[1319] = 134;
    exp_40_ram[1320] = 37;
    exp_40_ram[1321] = 5;
    exp_40_ram[1322] = 0;
    exp_40_ram[1323] = 39;
    exp_40_ram[1324] = 135;
    exp_40_ram[1325] = 38;
    exp_40_ram[1326] = 39;
    exp_40_ram[1327] = 230;
    exp_40_ram[1328] = 39;
    exp_40_ram[1329] = 135;
    exp_40_ram[1330] = 32;
    exp_40_ram[1331] = 0;
    exp_40_ram[1332] = 7;
    exp_40_ram[1333] = 36;
    exp_40_ram[1334] = 39;
    exp_40_ram[1335] = 231;
    exp_40_ram[1336] = 38;
    exp_40_ram[1337] = 39;
    exp_40_ram[1338] = 135;
    exp_40_ram[1339] = 46;
    exp_40_ram[1340] = 167;
    exp_40_ram[1341] = 135;
    exp_40_ram[1342] = 39;
    exp_40_ram[1343] = 34;
    exp_40_ram[1344] = 39;
    exp_40_ram[1345] = 32;
    exp_40_ram[1346] = 40;
    exp_40_ram[1347] = 8;
    exp_40_ram[1348] = 7;
    exp_40_ram[1349] = 38;
    exp_40_ram[1350] = 38;
    exp_40_ram[1351] = 37;
    exp_40_ram[1352] = 37;
    exp_40_ram[1353] = 240;
    exp_40_ram[1354] = 46;
    exp_40_ram[1355] = 39;
    exp_40_ram[1356] = 135;
    exp_40_ram[1357] = 32;
    exp_40_ram[1358] = 0;
    exp_40_ram[1359] = 39;
    exp_40_ram[1360] = 135;
    exp_40_ram[1361] = 46;
    exp_40_ram[1362] = 39;
    exp_40_ram[1363] = 38;
    exp_40_ram[1364] = 134;
    exp_40_ram[1365] = 37;
    exp_40_ram[1366] = 5;
    exp_40_ram[1367] = 0;
    exp_40_ram[1368] = 39;
    exp_40_ram[1369] = 135;
    exp_40_ram[1370] = 32;
    exp_40_ram[1371] = 0;
    exp_40_ram[1372] = 39;
    exp_40_ram[1373] = 197;
    exp_40_ram[1374] = 39;
    exp_40_ram[1375] = 135;
    exp_40_ram[1376] = 46;
    exp_40_ram[1377] = 39;
    exp_40_ram[1378] = 38;
    exp_40_ram[1379] = 134;
    exp_40_ram[1380] = 37;
    exp_40_ram[1381] = 0;
    exp_40_ram[1382] = 39;
    exp_40_ram[1383] = 135;
    exp_40_ram[1384] = 32;
    exp_40_ram[1385] = 0;
    exp_40_ram[1386] = 39;
    exp_40_ram[1387] = 199;
    exp_40_ram[1388] = 152;
    exp_40_ram[1389] = 39;
    exp_40_ram[1390] = 39;
    exp_40_ram[1391] = 104;
    exp_40_ram[1392] = 39;
    exp_40_ram[1393] = 135;
    exp_40_ram[1394] = 0;
    exp_40_ram[1395] = 39;
    exp_40_ram[1396] = 39;
    exp_40_ram[1397] = 38;
    exp_40_ram[1398] = 134;
    exp_40_ram[1399] = 37;
    exp_40_ram[1400] = 5;
    exp_40_ram[1401] = 0;
    exp_40_ram[1402] = 39;
    exp_40_ram[1403] = 133;
    exp_40_ram[1404] = 32;
    exp_40_ram[1405] = 36;
    exp_40_ram[1406] = 1;
    exp_40_ram[1407] = 128;
    exp_40_ram[1408] = 1;
    exp_40_ram[1409] = 38;
    exp_40_ram[1410] = 36;
    exp_40_ram[1411] = 4;
    exp_40_ram[1412] = 46;
    exp_40_ram[1413] = 34;
    exp_40_ram[1414] = 36;
    exp_40_ram[1415] = 38;
    exp_40_ram[1416] = 40;
    exp_40_ram[1417] = 42;
    exp_40_ram[1418] = 44;
    exp_40_ram[1419] = 46;
    exp_40_ram[1420] = 7;
    exp_40_ram[1421] = 44;
    exp_40_ram[1422] = 39;
    exp_40_ram[1423] = 135;
    exp_40_ram[1424] = 36;
    exp_40_ram[1425] = 39;
    exp_40_ram[1426] = 7;
    exp_40_ram[1427] = 38;
    exp_40_ram[1428] = 6;
    exp_40_ram[1429] = 133;
    exp_40_ram[1430] = 5;
    exp_40_ram[1431] = 240;
    exp_40_ram[1432] = 38;
    exp_40_ram[1433] = 39;
    exp_40_ram[1434] = 133;
    exp_40_ram[1435] = 32;
    exp_40_ram[1436] = 36;
    exp_40_ram[1437] = 1;
    exp_40_ram[1438] = 128;
    exp_40_ram[1439] = 1;
    exp_40_ram[1440] = 46;
    exp_40_ram[1441] = 44;
    exp_40_ram[1442] = 4;
    exp_40_ram[1443] = 7;
    exp_40_ram[1444] = 7;
    exp_40_ram[1445] = 71;
    exp_40_ram[1446] = 39;
    exp_40_ram[1447] = 167;
    exp_40_ram[1448] = 133;
    exp_40_ram[1449] = 5;
    exp_40_ram[1450] = 224;
    exp_40_ram[1451] = 0;
    exp_40_ram[1452] = 32;
    exp_40_ram[1453] = 36;
    exp_40_ram[1454] = 1;
    exp_40_ram[1455] = 128;
    exp_40_ram[1456] = 1;
    exp_40_ram[1457] = 38;
    exp_40_ram[1458] = 36;
    exp_40_ram[1459] = 4;
    exp_40_ram[1460] = 5;
    exp_40_ram[1461] = 224;
    exp_40_ram[1462] = 39;
    exp_40_ram[1463] = 39;
    exp_40_ram[1464] = 6;
    exp_40_ram[1465] = 134;
    exp_40_ram[1466] = 5;
    exp_40_ram[1467] = 240;
    exp_40_ram[1468] = 39;
    exp_40_ram[1469] = 39;
    exp_40_ram[1470] = 6;
    exp_40_ram[1471] = 134;
    exp_40_ram[1472] = 5;
    exp_40_ram[1473] = 240;
    exp_40_ram[1474] = 39;
    exp_40_ram[1475] = 39;
    exp_40_ram[1476] = 6;
    exp_40_ram[1477] = 134;
    exp_40_ram[1478] = 5;
    exp_40_ram[1479] = 240;
    exp_40_ram[1480] = 39;
    exp_40_ram[1481] = 39;
    exp_40_ram[1482] = 6;
    exp_40_ram[1483] = 134;
    exp_40_ram[1484] = 5;
    exp_40_ram[1485] = 240;
    exp_40_ram[1486] = 39;
    exp_40_ram[1487] = 39;
    exp_40_ram[1488] = 6;
    exp_40_ram[1489] = 134;
    exp_40_ram[1490] = 5;
    exp_40_ram[1491] = 240;
    exp_40_ram[1492] = 39;
    exp_40_ram[1493] = 39;
    exp_40_ram[1494] = 6;
    exp_40_ram[1495] = 134;
    exp_40_ram[1496] = 5;
    exp_40_ram[1497] = 240;
    exp_40_ram[1498] = 6;
    exp_40_ram[1499] = 6;
    exp_40_ram[1500] = 5;
    exp_40_ram[1501] = 240;
    exp_40_ram[1502] = 39;
    exp_40_ram[1503] = 39;
    exp_40_ram[1504] = 6;
    exp_40_ram[1505] = 134;
    exp_40_ram[1506] = 5;
    exp_40_ram[1507] = 240;
    exp_40_ram[1508] = 39;
    exp_40_ram[1509] = 39;
    exp_40_ram[1510] = 6;
    exp_40_ram[1511] = 134;
    exp_40_ram[1512] = 5;
    exp_40_ram[1513] = 240;
    exp_40_ram[1514] = 39;
    exp_40_ram[1515] = 39;
    exp_40_ram[1516] = 6;
    exp_40_ram[1517] = 134;
    exp_40_ram[1518] = 5;
    exp_40_ram[1519] = 240;
    exp_40_ram[1520] = 39;
    exp_40_ram[1521] = 39;
    exp_40_ram[1522] = 6;
    exp_40_ram[1523] = 134;
    exp_40_ram[1524] = 5;
    exp_40_ram[1525] = 240;
    exp_40_ram[1526] = 39;
    exp_40_ram[1527] = 39;
    exp_40_ram[1528] = 6;
    exp_40_ram[1529] = 134;
    exp_40_ram[1530] = 5;
    exp_40_ram[1531] = 240;
    exp_40_ram[1532] = 39;
    exp_40_ram[1533] = 39;
    exp_40_ram[1534] = 6;
    exp_40_ram[1535] = 134;
    exp_40_ram[1536] = 5;
    exp_40_ram[1537] = 240;
    exp_40_ram[1538] = 39;
    exp_40_ram[1539] = 39;
    exp_40_ram[1540] = 6;
    exp_40_ram[1541] = 134;
    exp_40_ram[1542] = 5;
    exp_40_ram[1543] = 240;
    exp_40_ram[1544] = 39;
    exp_40_ram[1545] = 39;
    exp_40_ram[1546] = 6;
    exp_40_ram[1547] = 134;
    exp_40_ram[1548] = 5;
    exp_40_ram[1549] = 240;
    exp_40_ram[1550] = 39;
    exp_40_ram[1551] = 39;
    exp_40_ram[1552] = 6;
    exp_40_ram[1553] = 134;
    exp_40_ram[1554] = 5;
    exp_40_ram[1555] = 240;
    exp_40_ram[1556] = 39;
    exp_40_ram[1557] = 39;
    exp_40_ram[1558] = 6;
    exp_40_ram[1559] = 134;
    exp_40_ram[1560] = 5;
    exp_40_ram[1561] = 240;
    exp_40_ram[1562] = 39;
    exp_40_ram[1563] = 39;
    exp_40_ram[1564] = 6;
    exp_40_ram[1565] = 134;
    exp_40_ram[1566] = 5;
    exp_40_ram[1567] = 240;
    exp_40_ram[1568] = 39;
    exp_40_ram[1569] = 39;
    exp_40_ram[1570] = 6;
    exp_40_ram[1571] = 134;
    exp_40_ram[1572] = 5;
    exp_40_ram[1573] = 240;
    exp_40_ram[1574] = 6;
    exp_40_ram[1575] = 6;
    exp_40_ram[1576] = 5;
    exp_40_ram[1577] = 240;
    exp_40_ram[1578] = 39;
    exp_40_ram[1579] = 39;
    exp_40_ram[1580] = 6;
    exp_40_ram[1581] = 134;
    exp_40_ram[1582] = 5;
    exp_40_ram[1583] = 240;
    exp_40_ram[1584] = 39;
    exp_40_ram[1585] = 39;
    exp_40_ram[1586] = 6;
    exp_40_ram[1587] = 134;
    exp_40_ram[1588] = 5;
    exp_40_ram[1589] = 240;
    exp_40_ram[1590] = 39;
    exp_40_ram[1591] = 39;
    exp_40_ram[1592] = 6;
    exp_40_ram[1593] = 134;
    exp_40_ram[1594] = 5;
    exp_40_ram[1595] = 240;
    exp_40_ram[1596] = 39;
    exp_40_ram[1597] = 39;
    exp_40_ram[1598] = 6;
    exp_40_ram[1599] = 134;
    exp_40_ram[1600] = 5;
    exp_40_ram[1601] = 240;
    exp_40_ram[1602] = 39;
    exp_40_ram[1603] = 39;
    exp_40_ram[1604] = 6;
    exp_40_ram[1605] = 134;
    exp_40_ram[1606] = 5;
    exp_40_ram[1607] = 240;
    exp_40_ram[1608] = 39;
    exp_40_ram[1609] = 39;
    exp_40_ram[1610] = 6;
    exp_40_ram[1611] = 134;
    exp_40_ram[1612] = 5;
    exp_40_ram[1613] = 240;
    exp_40_ram[1614] = 39;
    exp_40_ram[1615] = 39;
    exp_40_ram[1616] = 6;
    exp_40_ram[1617] = 134;
    exp_40_ram[1618] = 5;
    exp_40_ram[1619] = 240;
    exp_40_ram[1620] = 39;
    exp_40_ram[1621] = 39;
    exp_40_ram[1622] = 6;
    exp_40_ram[1623] = 134;
    exp_40_ram[1624] = 5;
    exp_40_ram[1625] = 240;
    exp_40_ram[1626] = 39;
    exp_40_ram[1627] = 39;
    exp_40_ram[1628] = 6;
    exp_40_ram[1629] = 134;
    exp_40_ram[1630] = 5;
    exp_40_ram[1631] = 240;
    exp_40_ram[1632] = 39;
    exp_40_ram[1633] = 39;
    exp_40_ram[1634] = 6;
    exp_40_ram[1635] = 134;
    exp_40_ram[1636] = 5;
    exp_40_ram[1637] = 240;
    exp_40_ram[1638] = 39;
    exp_40_ram[1639] = 39;
    exp_40_ram[1640] = 6;
    exp_40_ram[1641] = 134;
    exp_40_ram[1642] = 5;
    exp_40_ram[1643] = 240;
    exp_40_ram[1644] = 39;
    exp_40_ram[1645] = 39;
    exp_40_ram[1646] = 6;
    exp_40_ram[1647] = 134;
    exp_40_ram[1648] = 5;
    exp_40_ram[1649] = 240;
    exp_40_ram[1650] = 6;
    exp_40_ram[1651] = 6;
    exp_40_ram[1652] = 5;
    exp_40_ram[1653] = 240;
    exp_40_ram[1654] = 39;
    exp_40_ram[1655] = 39;
    exp_40_ram[1656] = 6;
    exp_40_ram[1657] = 134;
    exp_40_ram[1658] = 5;
    exp_40_ram[1659] = 240;
    exp_40_ram[1660] = 39;
    exp_40_ram[1661] = 39;
    exp_40_ram[1662] = 6;
    exp_40_ram[1663] = 134;
    exp_40_ram[1664] = 5;
    exp_40_ram[1665] = 240;
    exp_40_ram[1666] = 39;
    exp_40_ram[1667] = 39;
    exp_40_ram[1668] = 6;
    exp_40_ram[1669] = 134;
    exp_40_ram[1670] = 5;
    exp_40_ram[1671] = 240;
    exp_40_ram[1672] = 39;
    exp_40_ram[1673] = 39;
    exp_40_ram[1674] = 6;
    exp_40_ram[1675] = 134;
    exp_40_ram[1676] = 5;
    exp_40_ram[1677] = 240;
    exp_40_ram[1678] = 39;
    exp_40_ram[1679] = 39;
    exp_40_ram[1680] = 6;
    exp_40_ram[1681] = 134;
    exp_40_ram[1682] = 5;
    exp_40_ram[1683] = 240;
    exp_40_ram[1684] = 39;
    exp_40_ram[1685] = 39;
    exp_40_ram[1686] = 6;
    exp_40_ram[1687] = 134;
    exp_40_ram[1688] = 5;
    exp_40_ram[1689] = 240;
    exp_40_ram[1690] = 39;
    exp_40_ram[1691] = 39;
    exp_40_ram[1692] = 6;
    exp_40_ram[1693] = 134;
    exp_40_ram[1694] = 5;
    exp_40_ram[1695] = 240;
    exp_40_ram[1696] = 39;
    exp_40_ram[1697] = 39;
    exp_40_ram[1698] = 6;
    exp_40_ram[1699] = 134;
    exp_40_ram[1700] = 5;
    exp_40_ram[1701] = 240;
    exp_40_ram[1702] = 39;
    exp_40_ram[1703] = 39;
    exp_40_ram[1704] = 6;
    exp_40_ram[1705] = 134;
    exp_40_ram[1706] = 5;
    exp_40_ram[1707] = 240;
    exp_40_ram[1708] = 39;
    exp_40_ram[1709] = 39;
    exp_40_ram[1710] = 6;
    exp_40_ram[1711] = 134;
    exp_40_ram[1712] = 5;
    exp_40_ram[1713] = 240;
    exp_40_ram[1714] = 39;
    exp_40_ram[1715] = 39;
    exp_40_ram[1716] = 6;
    exp_40_ram[1717] = 134;
    exp_40_ram[1718] = 5;
    exp_40_ram[1719] = 240;
    exp_40_ram[1720] = 39;
    exp_40_ram[1721] = 39;
    exp_40_ram[1722] = 6;
    exp_40_ram[1723] = 134;
    exp_40_ram[1724] = 5;
    exp_40_ram[1725] = 240;
    exp_40_ram[1726] = 6;
    exp_40_ram[1727] = 6;
    exp_40_ram[1728] = 5;
    exp_40_ram[1729] = 240;
    exp_40_ram[1730] = 39;
    exp_40_ram[1731] = 39;
    exp_40_ram[1732] = 6;
    exp_40_ram[1733] = 134;
    exp_40_ram[1734] = 5;
    exp_40_ram[1735] = 240;
    exp_40_ram[1736] = 39;
    exp_40_ram[1737] = 39;
    exp_40_ram[1738] = 6;
    exp_40_ram[1739] = 134;
    exp_40_ram[1740] = 5;
    exp_40_ram[1741] = 240;
    exp_40_ram[1742] = 39;
    exp_40_ram[1743] = 39;
    exp_40_ram[1744] = 6;
    exp_40_ram[1745] = 134;
    exp_40_ram[1746] = 5;
    exp_40_ram[1747] = 240;
    exp_40_ram[1748] = 39;
    exp_40_ram[1749] = 39;
    exp_40_ram[1750] = 6;
    exp_40_ram[1751] = 134;
    exp_40_ram[1752] = 5;
    exp_40_ram[1753] = 240;
    exp_40_ram[1754] = 39;
    exp_40_ram[1755] = 39;
    exp_40_ram[1756] = 6;
    exp_40_ram[1757] = 134;
    exp_40_ram[1758] = 5;
    exp_40_ram[1759] = 240;
    exp_40_ram[1760] = 39;
    exp_40_ram[1761] = 39;
    exp_40_ram[1762] = 6;
    exp_40_ram[1763] = 134;
    exp_40_ram[1764] = 5;
    exp_40_ram[1765] = 240;
    exp_40_ram[1766] = 39;
    exp_40_ram[1767] = 39;
    exp_40_ram[1768] = 6;
    exp_40_ram[1769] = 134;
    exp_40_ram[1770] = 5;
    exp_40_ram[1771] = 240;
    exp_40_ram[1772] = 39;
    exp_40_ram[1773] = 39;
    exp_40_ram[1774] = 6;
    exp_40_ram[1775] = 134;
    exp_40_ram[1776] = 5;
    exp_40_ram[1777] = 240;
    exp_40_ram[1778] = 39;
    exp_40_ram[1779] = 39;
    exp_40_ram[1780] = 6;
    exp_40_ram[1781] = 134;
    exp_40_ram[1782] = 5;
    exp_40_ram[1783] = 240;
    exp_40_ram[1784] = 39;
    exp_40_ram[1785] = 39;
    exp_40_ram[1786] = 6;
    exp_40_ram[1787] = 134;
    exp_40_ram[1788] = 5;
    exp_40_ram[1789] = 240;
    exp_40_ram[1790] = 39;
    exp_40_ram[1791] = 39;
    exp_40_ram[1792] = 6;
    exp_40_ram[1793] = 134;
    exp_40_ram[1794] = 5;
    exp_40_ram[1795] = 240;
    exp_40_ram[1796] = 39;
    exp_40_ram[1797] = 39;
    exp_40_ram[1798] = 6;
    exp_40_ram[1799] = 134;
    exp_40_ram[1800] = 5;
    exp_40_ram[1801] = 240;
    exp_40_ram[1802] = 39;
    exp_40_ram[1803] = 39;
    exp_40_ram[1804] = 6;
    exp_40_ram[1805] = 134;
    exp_40_ram[1806] = 5;
    exp_40_ram[1807] = 240;
    exp_40_ram[1808] = 39;
    exp_40_ram[1809] = 39;
    exp_40_ram[1810] = 6;
    exp_40_ram[1811] = 134;
    exp_40_ram[1812] = 5;
    exp_40_ram[1813] = 240;
    exp_40_ram[1814] = 39;
    exp_40_ram[1815] = 39;
    exp_40_ram[1816] = 6;
    exp_40_ram[1817] = 134;
    exp_40_ram[1818] = 5;
    exp_40_ram[1819] = 240;
    exp_40_ram[1820] = 39;
    exp_40_ram[1821] = 39;
    exp_40_ram[1822] = 6;
    exp_40_ram[1823] = 134;
    exp_40_ram[1824] = 5;
    exp_40_ram[1825] = 240;
    exp_40_ram[1826] = 39;
    exp_40_ram[1827] = 39;
    exp_40_ram[1828] = 6;
    exp_40_ram[1829] = 134;
    exp_40_ram[1830] = 5;
    exp_40_ram[1831] = 240;
    exp_40_ram[1832] = 39;
    exp_40_ram[1833] = 39;
    exp_40_ram[1834] = 6;
    exp_40_ram[1835] = 134;
    exp_40_ram[1836] = 5;
    exp_40_ram[1837] = 240;
    exp_40_ram[1838] = 39;
    exp_40_ram[1839] = 39;
    exp_40_ram[1840] = 6;
    exp_40_ram[1841] = 134;
    exp_40_ram[1842] = 5;
    exp_40_ram[1843] = 240;
    exp_40_ram[1844] = 39;
    exp_40_ram[1845] = 39;
    exp_40_ram[1846] = 6;
    exp_40_ram[1847] = 134;
    exp_40_ram[1848] = 5;
    exp_40_ram[1849] = 240;
    exp_40_ram[1850] = 39;
    exp_40_ram[1851] = 39;
    exp_40_ram[1852] = 6;
    exp_40_ram[1853] = 134;
    exp_40_ram[1854] = 5;
    exp_40_ram[1855] = 240;
    exp_40_ram[1856] = 39;
    exp_40_ram[1857] = 39;
    exp_40_ram[1858] = 6;
    exp_40_ram[1859] = 134;
    exp_40_ram[1860] = 5;
    exp_40_ram[1861] = 240;
    exp_40_ram[1862] = 39;
    exp_40_ram[1863] = 39;
    exp_40_ram[1864] = 6;
    exp_40_ram[1865] = 134;
    exp_40_ram[1866] = 5;
    exp_40_ram[1867] = 240;
    exp_40_ram[1868] = 39;
    exp_40_ram[1869] = 39;
    exp_40_ram[1870] = 6;
    exp_40_ram[1871] = 134;
    exp_40_ram[1872] = 5;
    exp_40_ram[1873] = 240;
    exp_40_ram[1874] = 39;
    exp_40_ram[1875] = 39;
    exp_40_ram[1876] = 6;
    exp_40_ram[1877] = 134;
    exp_40_ram[1878] = 5;
    exp_40_ram[1879] = 240;
    exp_40_ram[1880] = 39;
    exp_40_ram[1881] = 39;
    exp_40_ram[1882] = 6;
    exp_40_ram[1883] = 134;
    exp_40_ram[1884] = 5;
    exp_40_ram[1885] = 240;
    exp_40_ram[1886] = 5;
    exp_40_ram[1887] = 224;
    exp_40_ram[1888] = 0;
    exp_40_ram[1889] = 32;
    exp_40_ram[1890] = 36;
    exp_40_ram[1891] = 1;
    exp_40_ram[1892] = 128;
    exp_40_ram[1893] = 1;
    exp_40_ram[1894] = 38;
    exp_40_ram[1895] = 36;
    exp_40_ram[1896] = 4;
    exp_40_ram[1897] = 240;
    exp_40_ram[1898] = 0;
    exp_40_ram[1899] = 32;
    exp_40_ram[1900] = 36;
    exp_40_ram[1901] = 1;
    exp_40_ram[1902] = 128;
    exp_40_ram[1903] = 0;
    exp_40_ram[1904] = 12;
    exp_40_ram[1905] = 12;
    exp_40_ram[1906] = 12;
    exp_40_ram[1907] = 12;
    exp_40_ram[1908] = 12;
    exp_40_ram[1909] = 12;
    exp_40_ram[1910] = 12;
    exp_40_ram[1911] = 12;
    exp_40_ram[1912] = 12;
    exp_40_ram[1913] = 12;
    exp_40_ram[1914] = 12;
    exp_40_ram[1915] = 12;
    exp_40_ram[1916] = 12;
    exp_40_ram[1917] = 12;
    exp_40_ram[1918] = 12;
    exp_40_ram[1919] = 12;
    exp_40_ram[1920] = 12;
    exp_40_ram[1921] = 14;
    exp_40_ram[1922] = 15;
    exp_40_ram[1923] = 14;
    exp_40_ram[1924] = 15;
    exp_40_ram[1925] = 14;
    exp_40_ram[1926] = 15;
    exp_40_ram[1927] = 15;
    exp_40_ram[1928] = 15;
    exp_40_ram[1929] = 15;
    exp_40_ram[1930] = 15;
    exp_40_ram[1931] = 15;
    exp_40_ram[1932] = 15;
    exp_40_ram[1933] = 14;
    exp_40_ram[1934] = 15;
    exp_40_ram[1935] = 15;
    exp_40_ram[1936] = 15;
    exp_40_ram[1937] = 15;
    exp_40_ram[1938] = 15;
    exp_40_ram[1939] = 14;
    exp_40_ram[1940] = 21;
    exp_40_ram[1941] = 21;
    exp_40_ram[1942] = 21;
    exp_40_ram[1943] = 21;
    exp_40_ram[1944] = 21;
    exp_40_ram[1945] = 21;
    exp_40_ram[1946] = 21;
    exp_40_ram[1947] = 21;
    exp_40_ram[1948] = 21;
    exp_40_ram[1949] = 21;
    exp_40_ram[1950] = 21;
    exp_40_ram[1951] = 21;
    exp_40_ram[1952] = 21;
    exp_40_ram[1953] = 21;
    exp_40_ram[1954] = 21;
    exp_40_ram[1955] = 21;
    exp_40_ram[1956] = 21;
    exp_40_ram[1957] = 21;
    exp_40_ram[1958] = 21;
    exp_40_ram[1959] = 21;
    exp_40_ram[1960] = 21;
    exp_40_ram[1961] = 21;
    exp_40_ram[1962] = 21;
    exp_40_ram[1963] = 21;
    exp_40_ram[1964] = 21;
    exp_40_ram[1965] = 21;
    exp_40_ram[1966] = 21;
    exp_40_ram[1967] = 21;
    exp_40_ram[1968] = 21;
    exp_40_ram[1969] = 21;
    exp_40_ram[1970] = 21;
    exp_40_ram[1971] = 21;
    exp_40_ram[1972] = 21;
    exp_40_ram[1973] = 21;
    exp_40_ram[1974] = 21;
    exp_40_ram[1975] = 21;
    exp_40_ram[1976] = 21;
    exp_40_ram[1977] = 21;
    exp_40_ram[1978] = 21;
    exp_40_ram[1979] = 21;
    exp_40_ram[1980] = 21;
    exp_40_ram[1981] = 21;
    exp_40_ram[1982] = 21;
    exp_40_ram[1983] = 21;
    exp_40_ram[1984] = 21;
    exp_40_ram[1985] = 21;
    exp_40_ram[1986] = 21;
    exp_40_ram[1987] = 21;
    exp_40_ram[1988] = 21;
    exp_40_ram[1989] = 21;
    exp_40_ram[1990] = 21;
    exp_40_ram[1991] = 15;
    exp_40_ram[1992] = 21;
    exp_40_ram[1993] = 21;
    exp_40_ram[1994] = 21;
    exp_40_ram[1995] = 21;
    exp_40_ram[1996] = 21;
    exp_40_ram[1997] = 21;
    exp_40_ram[1998] = 21;
    exp_40_ram[1999] = 21;
    exp_40_ram[2000] = 21;
    exp_40_ram[2001] = 15;
    exp_40_ram[2002] = 18;
    exp_40_ram[2003] = 15;
    exp_40_ram[2004] = 21;
    exp_40_ram[2005] = 21;
    exp_40_ram[2006] = 21;
    exp_40_ram[2007] = 21;
    exp_40_ram[2008] = 15;
    exp_40_ram[2009] = 21;
    exp_40_ram[2010] = 21;
    exp_40_ram[2011] = 21;
    exp_40_ram[2012] = 21;
    exp_40_ram[2013] = 21;
    exp_40_ram[2014] = 15;
    exp_40_ram[2015] = 20;
    exp_40_ram[2016] = 21;
    exp_40_ram[2017] = 21;
    exp_40_ram[2018] = 19;
    exp_40_ram[2019] = 21;
    exp_40_ram[2020] = 15;
    exp_40_ram[2021] = 21;
    exp_40_ram[2022] = 21;
    exp_40_ram[2023] = 15;
    exp_40_ram[2024] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 55;
    exp_33_ram[32] = 19;
    exp_33_ram[33] = 239;
    exp_33_ram[34] = 111;
    exp_33_ram[35] = 0;
    exp_33_ram[36] = 115;
    exp_33_ram[37] = 97;
    exp_33_ram[38] = 46;
    exp_33_ram[39] = 108;
    exp_33_ram[40] = 72;
    exp_33_ram[41] = 111;
    exp_33_ram[42] = 49;
    exp_33_ram[43] = 105;
    exp_33_ram[44] = 50;
    exp_33_ram[45] = 105;
    exp_33_ram[46] = 72;
    exp_33_ram[47] = 51;
    exp_33_ram[48] = 105;
    exp_33_ram[49] = 52;
    exp_33_ram[50] = 105;
    exp_33_ram[51] = 112;
    exp_33_ram[52] = 0;
    exp_33_ram[53] = 115;
    exp_33_ram[54] = 99;
    exp_33_ram[55] = 46;
    exp_33_ram[56] = 108;
    exp_33_ram[57] = 121;
    exp_33_ram[58] = 109;
    exp_33_ram[59] = 109;
    exp_33_ram[60] = 46;
    exp_33_ram[61] = 115;
    exp_33_ram[62] = 109;
    exp_33_ram[63] = 46;
    exp_33_ram[64] = 115;
    exp_33_ram[65] = 99;
    exp_33_ram[66] = 46;
    exp_33_ram[67] = 109;
    exp_33_ram[68] = 104;
    exp_33_ram[69] = 46;
    exp_33_ram[70] = 53;
    exp_33_ram[71] = 105;
    exp_33_ram[72] = 115;
    exp_33_ram[73] = 104;
    exp_33_ram[74] = 46;
    exp_33_ram[75] = 54;
    exp_33_ram[76] = 105;
    exp_33_ram[77] = 115;
    exp_33_ram[78] = 115;
    exp_33_ram[79] = 46;
    exp_33_ram[80] = 97;
    exp_33_ram[81] = 49;
    exp_33_ram[82] = 97;
    exp_33_ram[83] = 97;
    exp_33_ram[84] = 50;
    exp_33_ram[85] = 97;
    exp_33_ram[86] = 97;
    exp_33_ram[87] = 51;
    exp_33_ram[88] = 97;
    exp_33_ram[89] = 115;
    exp_33_ram[90] = 0;
    exp_33_ram[91] = 97;
    exp_33_ram[92] = 97;
    exp_33_ram[93] = 0;
    exp_33_ram[94] = 115;
    exp_33_ram[95] = 98;
    exp_33_ram[96] = 46;
    exp_33_ram[97] = 97;
    exp_33_ram[98] = 97;
    exp_33_ram[99] = 0;
    exp_33_ram[100] = 97;
    exp_33_ram[101] = 97;
    exp_33_ram[102] = 108;
    exp_33_ram[103] = 108;
    exp_33_ram[104] = 52;
    exp_33_ram[105] = 102;
    exp_33_ram[106] = 97;
    exp_33_ram[107] = 97;
    exp_33_ram[108] = 0;
    exp_33_ram[109] = 115;
    exp_33_ram[110] = 99;
    exp_33_ram[111] = 46;
    exp_33_ram[112] = 115;
    exp_33_ram[113] = 112;
    exp_33_ram[114] = 46;
    exp_33_ram[115] = 97;
    exp_33_ram[116] = 52;
    exp_33_ram[117] = 97;
    exp_33_ram[118] = 102;
    exp_33_ram[119] = 100;
    exp_33_ram[120] = 97;
    exp_33_ram[121] = 49;
    exp_33_ram[122] = 100;
    exp_33_ram[123] = 97;
    exp_33_ram[124] = 102;
    exp_33_ram[125] = 115;
    exp_33_ram[126] = 0;
    exp_33_ram[127] = 115;
    exp_33_ram[128] = 116;
    exp_33_ram[129] = 46;
    exp_33_ram[130] = 49;
    exp_33_ram[131] = 0;
    exp_33_ram[132] = 50;
    exp_33_ram[133] = 51;
    exp_33_ram[134] = 109;
    exp_33_ram[135] = 101;
    exp_33_ram[136] = 46;
    exp_33_ram[137] = 97;
    exp_33_ram[138] = 0;
    exp_33_ram[139] = 98;
    exp_33_ram[140] = 0;
    exp_33_ram[141] = 99;
    exp_33_ram[142] = 0;
    exp_33_ram[143] = 100;
    exp_33_ram[144] = 0;
    exp_33_ram[145] = 115;
    exp_33_ram[146] = 101;
    exp_33_ram[147] = 46;
    exp_33_ram[148] = 116;
    exp_33_ram[149] = 46;
    exp_33_ram[150] = 84;
    exp_33_ram[151] = 83;
    exp_33_ram[152] = 49;
    exp_33_ram[153] = 48;
    exp_33_ram[154] = 58;
    exp_33_ram[155] = 50;
    exp_33_ram[156] = 10;
    exp_33_ram[157] = 84;
    exp_33_ram[158] = 83;
    exp_33_ram[159] = 49;
    exp_33_ram[160] = 49;
    exp_33_ram[161] = 58;
    exp_33_ram[162] = 50;
    exp_33_ram[163] = 10;
    exp_33_ram[164] = 55;
    exp_33_ram[165] = 105;
    exp_33_ram[166] = 56;
    exp_33_ram[167] = 105;
    exp_33_ram[168] = 57;
    exp_33_ram[169] = 105;
    exp_33_ram[170] = 84;
    exp_33_ram[171] = 83;
    exp_33_ram[172] = 49;
    exp_33_ram[173] = 50;
    exp_33_ram[174] = 58;
    exp_33_ram[175] = 50;
    exp_33_ram[176] = 10;
    exp_33_ram[177] = 49;
    exp_33_ram[178] = 97;
    exp_33_ram[179] = 49;
    exp_33_ram[180] = 97;
    exp_33_ram[181] = 49;
    exp_33_ram[182] = 97;
    exp_33_ram[183] = 116;
    exp_33_ram[184] = 32;
    exp_33_ram[185] = 110;
    exp_33_ram[186] = 46;
    exp_33_ram[187] = 37;
    exp_33_ram[188] = 37;
    exp_33_ram[189] = 49;
    exp_33_ram[190] = 0;
    exp_33_ram[191] = 37;
    exp_33_ram[192] = 119;
    exp_33_ram[193] = 104;
    exp_33_ram[194] = 32;
    exp_33_ram[195] = 46;
    exp_33_ram[196] = 0;
    exp_33_ram[197] = 37;
    exp_33_ram[198] = 37;
    exp_33_ram[199] = 37;
    exp_33_ram[200] = 141;
    exp_33_ram[201] = 247;
    exp_33_ram[202] = 241;
    exp_33_ram[203] = 181;
    exp_33_ram[204] = 45;
    exp_33_ram[205] = 226;
    exp_33_ram[206] = 252;
    exp_33_ram[207] = 77;
    exp_33_ram[208] = 123;
    exp_33_ram[209] = 225;
    exp_33_ram[210] = 154;
    exp_33_ram[211] = 153;
    exp_33_ram[212] = 0;
    exp_33_ram[213] = 0;
    exp_33_ram[214] = 0;
    exp_33_ram[215] = 0;
    exp_33_ram[216] = 0;
    exp_33_ram[217] = 0;
    exp_33_ram[218] = 0;
    exp_33_ram[219] = 0;
    exp_33_ram[220] = 0;
    exp_33_ram[221] = 0;
    exp_33_ram[222] = 0;
    exp_33_ram[223] = 0;
    exp_33_ram[224] = 0;
    exp_33_ram[225] = 128;
    exp_33_ram[226] = 0;
    exp_33_ram[227] = 208;
    exp_33_ram[228] = 0;
    exp_33_ram[229] = 132;
    exp_33_ram[230] = 0;
    exp_33_ram[231] = 101;
    exp_33_ram[232] = 0;
    exp_33_ram[233] = 0;
    exp_33_ram[234] = 0;
    exp_33_ram[235] = 0;
    exp_33_ram[236] = 0;
    exp_33_ram[237] = 0;
    exp_33_ram[238] = 0;
    exp_33_ram[239] = 0;
    exp_33_ram[240] = 35;
    exp_33_ram[241] = 103;
    exp_33_ram[242] = 147;
    exp_33_ram[243] = 19;
    exp_33_ram[244] = 51;
    exp_33_ram[245] = 3;
    exp_33_ram[246] = 99;
    exp_33_ram[247] = 103;
    exp_33_ram[248] = 19;
    exp_33_ram[249] = 35;
    exp_33_ram[250] = 111;
    exp_33_ram[251] = 19;
    exp_33_ram[252] = 183;
    exp_33_ram[253] = 35;
    exp_33_ram[254] = 3;
    exp_33_ram[255] = 35;
    exp_33_ram[256] = 147;
    exp_33_ram[257] = 239;
    exp_33_ram[258] = 147;
    exp_33_ram[259] = 131;
    exp_33_ram[260] = 35;
    exp_33_ram[261] = 3;
    exp_33_ram[262] = 19;
    exp_33_ram[263] = 19;
    exp_33_ram[264] = 103;
    exp_33_ram[265] = 19;
    exp_33_ram[266] = 35;
    exp_33_ram[267] = 19;
    exp_33_ram[268] = 147;
    exp_33_ram[269] = 35;
    exp_33_ram[270] = 35;
    exp_33_ram[271] = 35;
    exp_33_ram[272] = 163;
    exp_33_ram[273] = 19;
    exp_33_ram[274] = 3;
    exp_33_ram[275] = 19;
    exp_33_ram[276] = 103;
    exp_33_ram[277] = 19;
    exp_33_ram[278] = 35;
    exp_33_ram[279] = 35;
    exp_33_ram[280] = 19;
    exp_33_ram[281] = 147;
    exp_33_ram[282] = 35;
    exp_33_ram[283] = 35;
    exp_33_ram[284] = 35;
    exp_33_ram[285] = 163;
    exp_33_ram[286] = 131;
    exp_33_ram[287] = 99;
    exp_33_ram[288] = 131;
    exp_33_ram[289] = 19;
    exp_33_ram[290] = 239;
    exp_33_ram[291] = 19;
    exp_33_ram[292] = 131;
    exp_33_ram[293] = 3;
    exp_33_ram[294] = 19;
    exp_33_ram[295] = 103;
    exp_33_ram[296] = 19;
    exp_33_ram[297] = 35;
    exp_33_ram[298] = 19;
    exp_33_ram[299] = 35;
    exp_33_ram[300] = 35;
    exp_33_ram[301] = 131;
    exp_33_ram[302] = 35;
    exp_33_ram[303] = 111;
    exp_33_ram[304] = 131;
    exp_33_ram[305] = 147;
    exp_33_ram[306] = 35;
    exp_33_ram[307] = 131;
    exp_33_ram[308] = 131;
    exp_33_ram[309] = 99;
    exp_33_ram[310] = 131;
    exp_33_ram[311] = 19;
    exp_33_ram[312] = 35;
    exp_33_ram[313] = 227;
    exp_33_ram[314] = 3;
    exp_33_ram[315] = 131;
    exp_33_ram[316] = 179;
    exp_33_ram[317] = 19;
    exp_33_ram[318] = 3;
    exp_33_ram[319] = 19;
    exp_33_ram[320] = 103;
    exp_33_ram[321] = 19;
    exp_33_ram[322] = 35;
    exp_33_ram[323] = 19;
    exp_33_ram[324] = 147;
    exp_33_ram[325] = 163;
    exp_33_ram[326] = 3;
    exp_33_ram[327] = 147;
    exp_33_ram[328] = 99;
    exp_33_ram[329] = 3;
    exp_33_ram[330] = 147;
    exp_33_ram[331] = 99;
    exp_33_ram[332] = 147;
    exp_33_ram[333] = 111;
    exp_33_ram[334] = 147;
    exp_33_ram[335] = 147;
    exp_33_ram[336] = 147;
    exp_33_ram[337] = 19;
    exp_33_ram[338] = 3;
    exp_33_ram[339] = 19;
    exp_33_ram[340] = 103;
    exp_33_ram[341] = 19;
    exp_33_ram[342] = 35;
    exp_33_ram[343] = 35;
    exp_33_ram[344] = 19;
    exp_33_ram[345] = 35;
    exp_33_ram[346] = 35;
    exp_33_ram[347] = 111;
    exp_33_ram[348] = 3;
    exp_33_ram[349] = 147;
    exp_33_ram[350] = 147;
    exp_33_ram[351] = 179;
    exp_33_ram[352] = 147;
    exp_33_ram[353] = 19;
    exp_33_ram[354] = 131;
    exp_33_ram[355] = 131;
    exp_33_ram[356] = 147;
    exp_33_ram[357] = 3;
    exp_33_ram[358] = 35;
    exp_33_ram[359] = 131;
    exp_33_ram[360] = 179;
    exp_33_ram[361] = 147;
    exp_33_ram[362] = 35;
    exp_33_ram[363] = 131;
    exp_33_ram[364] = 131;
    exp_33_ram[365] = 131;
    exp_33_ram[366] = 19;
    exp_33_ram[367] = 239;
    exp_33_ram[368] = 147;
    exp_33_ram[369] = 227;
    exp_33_ram[370] = 131;
    exp_33_ram[371] = 19;
    exp_33_ram[372] = 131;
    exp_33_ram[373] = 3;
    exp_33_ram[374] = 19;
    exp_33_ram[375] = 103;
    exp_33_ram[376] = 19;
    exp_33_ram[377] = 35;
    exp_33_ram[378] = 35;
    exp_33_ram[379] = 19;
    exp_33_ram[380] = 35;
    exp_33_ram[381] = 35;
    exp_33_ram[382] = 35;
    exp_33_ram[383] = 35;
    exp_33_ram[384] = 35;
    exp_33_ram[385] = 35;
    exp_33_ram[386] = 35;
    exp_33_ram[387] = 35;
    exp_33_ram[388] = 131;
    exp_33_ram[389] = 35;
    exp_33_ram[390] = 131;
    exp_33_ram[391] = 147;
    exp_33_ram[392] = 99;
    exp_33_ram[393] = 131;
    exp_33_ram[394] = 147;
    exp_33_ram[395] = 99;
    exp_33_ram[396] = 131;
    exp_33_ram[397] = 35;
    exp_33_ram[398] = 111;
    exp_33_ram[399] = 131;
    exp_33_ram[400] = 19;
    exp_33_ram[401] = 35;
    exp_33_ram[402] = 3;
    exp_33_ram[403] = 131;
    exp_33_ram[404] = 19;
    exp_33_ram[405] = 131;
    exp_33_ram[406] = 19;
    exp_33_ram[407] = 231;
    exp_33_ram[408] = 131;
    exp_33_ram[409] = 147;
    exp_33_ram[410] = 35;
    exp_33_ram[411] = 3;
    exp_33_ram[412] = 131;
    exp_33_ram[413] = 227;
    exp_33_ram[414] = 111;
    exp_33_ram[415] = 131;
    exp_33_ram[416] = 147;
    exp_33_ram[417] = 35;
    exp_33_ram[418] = 3;
    exp_33_ram[419] = 131;
    exp_33_ram[420] = 179;
    exp_33_ram[421] = 3;
    exp_33_ram[422] = 131;
    exp_33_ram[423] = 19;
    exp_33_ram[424] = 35;
    exp_33_ram[425] = 3;
    exp_33_ram[426] = 131;
    exp_33_ram[427] = 19;
    exp_33_ram[428] = 131;
    exp_33_ram[429] = 231;
    exp_33_ram[430] = 131;
    exp_33_ram[431] = 227;
    exp_33_ram[432] = 131;
    exp_33_ram[433] = 147;
    exp_33_ram[434] = 99;
    exp_33_ram[435] = 111;
    exp_33_ram[436] = 131;
    exp_33_ram[437] = 19;
    exp_33_ram[438] = 35;
    exp_33_ram[439] = 3;
    exp_33_ram[440] = 131;
    exp_33_ram[441] = 19;
    exp_33_ram[442] = 131;
    exp_33_ram[443] = 19;
    exp_33_ram[444] = 231;
    exp_33_ram[445] = 3;
    exp_33_ram[446] = 131;
    exp_33_ram[447] = 179;
    exp_33_ram[448] = 3;
    exp_33_ram[449] = 227;
    exp_33_ram[450] = 131;
    exp_33_ram[451] = 19;
    exp_33_ram[452] = 131;
    exp_33_ram[453] = 3;
    exp_33_ram[454] = 19;
    exp_33_ram[455] = 103;
    exp_33_ram[456] = 19;
    exp_33_ram[457] = 35;
    exp_33_ram[458] = 35;
    exp_33_ram[459] = 19;
    exp_33_ram[460] = 35;
    exp_33_ram[461] = 35;
    exp_33_ram[462] = 35;
    exp_33_ram[463] = 35;
    exp_33_ram[464] = 35;
    exp_33_ram[465] = 35;
    exp_33_ram[466] = 147;
    exp_33_ram[467] = 35;
    exp_33_ram[468] = 163;
    exp_33_ram[469] = 131;
    exp_33_ram[470] = 147;
    exp_33_ram[471] = 99;
    exp_33_ram[472] = 131;
    exp_33_ram[473] = 99;
    exp_33_ram[474] = 131;
    exp_33_ram[475] = 147;
    exp_33_ram[476] = 99;
    exp_33_ram[477] = 131;
    exp_33_ram[478] = 99;
    exp_33_ram[479] = 131;
    exp_33_ram[480] = 147;
    exp_33_ram[481] = 99;
    exp_33_ram[482] = 131;
    exp_33_ram[483] = 147;
    exp_33_ram[484] = 35;
    exp_33_ram[485] = 111;
    exp_33_ram[486] = 131;
    exp_33_ram[487] = 19;
    exp_33_ram[488] = 35;
    exp_33_ram[489] = 3;
    exp_33_ram[490] = 179;
    exp_33_ram[491] = 19;
    exp_33_ram[492] = 35;
    exp_33_ram[493] = 3;
    exp_33_ram[494] = 131;
    exp_33_ram[495] = 99;
    exp_33_ram[496] = 3;
    exp_33_ram[497] = 147;
    exp_33_ram[498] = 227;
    exp_33_ram[499] = 111;
    exp_33_ram[500] = 131;
    exp_33_ram[501] = 19;
    exp_33_ram[502] = 35;
    exp_33_ram[503] = 3;
    exp_33_ram[504] = 179;
    exp_33_ram[505] = 19;
    exp_33_ram[506] = 35;
    exp_33_ram[507] = 131;
    exp_33_ram[508] = 147;
    exp_33_ram[509] = 99;
    exp_33_ram[510] = 3;
    exp_33_ram[511] = 131;
    exp_33_ram[512] = 99;
    exp_33_ram[513] = 3;
    exp_33_ram[514] = 147;
    exp_33_ram[515] = 227;
    exp_33_ram[516] = 131;
    exp_33_ram[517] = 147;
    exp_33_ram[518] = 99;
    exp_33_ram[519] = 131;
    exp_33_ram[520] = 147;
    exp_33_ram[521] = 99;
    exp_33_ram[522] = 131;
    exp_33_ram[523] = 99;
    exp_33_ram[524] = 3;
    exp_33_ram[525] = 131;
    exp_33_ram[526] = 99;
    exp_33_ram[527] = 3;
    exp_33_ram[528] = 131;
    exp_33_ram[529] = 99;
    exp_33_ram[530] = 131;
    exp_33_ram[531] = 147;
    exp_33_ram[532] = 35;
    exp_33_ram[533] = 131;
    exp_33_ram[534] = 99;
    exp_33_ram[535] = 3;
    exp_33_ram[536] = 147;
    exp_33_ram[537] = 99;
    exp_33_ram[538] = 131;
    exp_33_ram[539] = 147;
    exp_33_ram[540] = 35;
    exp_33_ram[541] = 3;
    exp_33_ram[542] = 147;
    exp_33_ram[543] = 99;
    exp_33_ram[544] = 131;
    exp_33_ram[545] = 147;
    exp_33_ram[546] = 99;
    exp_33_ram[547] = 3;
    exp_33_ram[548] = 147;
    exp_33_ram[549] = 99;
    exp_33_ram[550] = 131;
    exp_33_ram[551] = 19;
    exp_33_ram[552] = 35;
    exp_33_ram[553] = 3;
    exp_33_ram[554] = 179;
    exp_33_ram[555] = 19;
    exp_33_ram[556] = 35;
    exp_33_ram[557] = 111;
    exp_33_ram[558] = 3;
    exp_33_ram[559] = 147;
    exp_33_ram[560] = 99;
    exp_33_ram[561] = 131;
    exp_33_ram[562] = 147;
    exp_33_ram[563] = 99;
    exp_33_ram[564] = 3;
    exp_33_ram[565] = 147;
    exp_33_ram[566] = 99;
    exp_33_ram[567] = 131;
    exp_33_ram[568] = 19;
    exp_33_ram[569] = 35;
    exp_33_ram[570] = 3;
    exp_33_ram[571] = 179;
    exp_33_ram[572] = 19;
    exp_33_ram[573] = 35;
    exp_33_ram[574] = 111;
    exp_33_ram[575] = 3;
    exp_33_ram[576] = 147;
    exp_33_ram[577] = 99;
    exp_33_ram[578] = 3;
    exp_33_ram[579] = 147;
    exp_33_ram[580] = 99;
    exp_33_ram[581] = 131;
    exp_33_ram[582] = 19;
    exp_33_ram[583] = 35;
    exp_33_ram[584] = 3;
    exp_33_ram[585] = 179;
    exp_33_ram[586] = 19;
    exp_33_ram[587] = 35;
    exp_33_ram[588] = 3;
    exp_33_ram[589] = 147;
    exp_33_ram[590] = 99;
    exp_33_ram[591] = 131;
    exp_33_ram[592] = 19;
    exp_33_ram[593] = 35;
    exp_33_ram[594] = 3;
    exp_33_ram[595] = 179;
    exp_33_ram[596] = 19;
    exp_33_ram[597] = 35;
    exp_33_ram[598] = 3;
    exp_33_ram[599] = 147;
    exp_33_ram[600] = 99;
    exp_33_ram[601] = 131;
    exp_33_ram[602] = 99;
    exp_33_ram[603] = 131;
    exp_33_ram[604] = 19;
    exp_33_ram[605] = 35;
    exp_33_ram[606] = 3;
    exp_33_ram[607] = 179;
    exp_33_ram[608] = 19;
    exp_33_ram[609] = 35;
    exp_33_ram[610] = 111;
    exp_33_ram[611] = 131;
    exp_33_ram[612] = 147;
    exp_33_ram[613] = 99;
    exp_33_ram[614] = 131;
    exp_33_ram[615] = 19;
    exp_33_ram[616] = 35;
    exp_33_ram[617] = 3;
    exp_33_ram[618] = 179;
    exp_33_ram[619] = 19;
    exp_33_ram[620] = 35;
    exp_33_ram[621] = 111;
    exp_33_ram[622] = 131;
    exp_33_ram[623] = 147;
    exp_33_ram[624] = 99;
    exp_33_ram[625] = 131;
    exp_33_ram[626] = 19;
    exp_33_ram[627] = 35;
    exp_33_ram[628] = 3;
    exp_33_ram[629] = 179;
    exp_33_ram[630] = 19;
    exp_33_ram[631] = 35;
    exp_33_ram[632] = 131;
    exp_33_ram[633] = 3;
    exp_33_ram[634] = 131;
    exp_33_ram[635] = 3;
    exp_33_ram[636] = 131;
    exp_33_ram[637] = 3;
    exp_33_ram[638] = 131;
    exp_33_ram[639] = 3;
    exp_33_ram[640] = 239;
    exp_33_ram[641] = 147;
    exp_33_ram[642] = 19;
    exp_33_ram[643] = 131;
    exp_33_ram[644] = 3;
    exp_33_ram[645] = 19;
    exp_33_ram[646] = 103;
    exp_33_ram[647] = 19;
    exp_33_ram[648] = 35;
    exp_33_ram[649] = 35;
    exp_33_ram[650] = 19;
    exp_33_ram[651] = 35;
    exp_33_ram[652] = 35;
    exp_33_ram[653] = 35;
    exp_33_ram[654] = 35;
    exp_33_ram[655] = 35;
    exp_33_ram[656] = 35;
    exp_33_ram[657] = 35;
    exp_33_ram[658] = 163;
    exp_33_ram[659] = 35;
    exp_33_ram[660] = 131;
    exp_33_ram[661] = 99;
    exp_33_ram[662] = 131;
    exp_33_ram[663] = 147;
    exp_33_ram[664] = 35;
    exp_33_ram[665] = 131;
    exp_33_ram[666] = 147;
    exp_33_ram[667] = 99;
    exp_33_ram[668] = 131;
    exp_33_ram[669] = 99;
    exp_33_ram[670] = 3;
    exp_33_ram[671] = 131;
    exp_33_ram[672] = 179;
    exp_33_ram[673] = 163;
    exp_33_ram[674] = 3;
    exp_33_ram[675] = 147;
    exp_33_ram[676] = 99;
    exp_33_ram[677] = 131;
    exp_33_ram[678] = 147;
    exp_33_ram[679] = 147;
    exp_33_ram[680] = 111;
    exp_33_ram[681] = 131;
    exp_33_ram[682] = 147;
    exp_33_ram[683] = 99;
    exp_33_ram[684] = 147;
    exp_33_ram[685] = 111;
    exp_33_ram[686] = 147;
    exp_33_ram[687] = 3;
    exp_33_ram[688] = 179;
    exp_33_ram[689] = 147;
    exp_33_ram[690] = 147;
    exp_33_ram[691] = 147;
    exp_33_ram[692] = 3;
    exp_33_ram[693] = 147;
    exp_33_ram[694] = 35;
    exp_33_ram[695] = 147;
    exp_33_ram[696] = 51;
    exp_33_ram[697] = 35;
    exp_33_ram[698] = 3;
    exp_33_ram[699] = 131;
    exp_33_ram[700] = 179;
    exp_33_ram[701] = 35;
    exp_33_ram[702] = 131;
    exp_33_ram[703] = 99;
    exp_33_ram[704] = 3;
    exp_33_ram[705] = 147;
    exp_33_ram[706] = 227;
    exp_33_ram[707] = 131;
    exp_33_ram[708] = 19;
    exp_33_ram[709] = 131;
    exp_33_ram[710] = 35;
    exp_33_ram[711] = 131;
    exp_33_ram[712] = 35;
    exp_33_ram[713] = 131;
    exp_33_ram[714] = 35;
    exp_33_ram[715] = 131;
    exp_33_ram[716] = 19;
    exp_33_ram[717] = 131;
    exp_33_ram[718] = 131;
    exp_33_ram[719] = 3;
    exp_33_ram[720] = 131;
    exp_33_ram[721] = 3;
    exp_33_ram[722] = 239;
    exp_33_ram[723] = 147;
    exp_33_ram[724] = 19;
    exp_33_ram[725] = 131;
    exp_33_ram[726] = 3;
    exp_33_ram[727] = 19;
    exp_33_ram[728] = 103;
    exp_33_ram[729] = 19;
    exp_33_ram[730] = 35;
    exp_33_ram[731] = 35;
    exp_33_ram[732] = 19;
    exp_33_ram[733] = 35;
    exp_33_ram[734] = 35;
    exp_33_ram[735] = 35;
    exp_33_ram[736] = 35;
    exp_33_ram[737] = 35;
    exp_33_ram[738] = 35;
    exp_33_ram[739] = 131;
    exp_33_ram[740] = 227;
    exp_33_ram[741] = 147;
    exp_33_ram[742] = 35;
    exp_33_ram[743] = 111;
    exp_33_ram[744] = 131;
    exp_33_ram[745] = 3;
    exp_33_ram[746] = 147;
    exp_33_ram[747] = 99;
    exp_33_ram[748] = 131;
    exp_33_ram[749] = 3;
    exp_33_ram[750] = 131;
    exp_33_ram[751] = 19;
    exp_33_ram[752] = 35;
    exp_33_ram[753] = 3;
    exp_33_ram[754] = 131;
    exp_33_ram[755] = 19;
    exp_33_ram[756] = 131;
    exp_33_ram[757] = 231;
    exp_33_ram[758] = 131;
    exp_33_ram[759] = 147;
    exp_33_ram[760] = 35;
    exp_33_ram[761] = 111;
    exp_33_ram[762] = 131;
    exp_33_ram[763] = 147;
    exp_33_ram[764] = 35;
    exp_33_ram[765] = 35;
    exp_33_ram[766] = 131;
    exp_33_ram[767] = 131;
    exp_33_ram[768] = 147;
    exp_33_ram[769] = 19;
    exp_33_ram[770] = 99;
    exp_33_ram[771] = 19;
    exp_33_ram[772] = 183;
    exp_33_ram[773] = 147;
    exp_33_ram[774] = 179;
    exp_33_ram[775] = 131;
    exp_33_ram[776] = 103;
    exp_33_ram[777] = 131;
    exp_33_ram[778] = 147;
    exp_33_ram[779] = 35;
    exp_33_ram[780] = 131;
    exp_33_ram[781] = 147;
    exp_33_ram[782] = 35;
    exp_33_ram[783] = 147;
    exp_33_ram[784] = 35;
    exp_33_ram[785] = 111;
    exp_33_ram[786] = 131;
    exp_33_ram[787] = 147;
    exp_33_ram[788] = 35;
    exp_33_ram[789] = 131;
    exp_33_ram[790] = 147;
    exp_33_ram[791] = 35;
    exp_33_ram[792] = 147;
    exp_33_ram[793] = 35;
    exp_33_ram[794] = 111;
    exp_33_ram[795] = 131;
    exp_33_ram[796] = 147;
    exp_33_ram[797] = 35;
    exp_33_ram[798] = 131;
    exp_33_ram[799] = 147;
    exp_33_ram[800] = 35;
    exp_33_ram[801] = 147;
    exp_33_ram[802] = 35;
    exp_33_ram[803] = 111;
    exp_33_ram[804] = 131;
    exp_33_ram[805] = 147;
    exp_33_ram[806] = 35;
    exp_33_ram[807] = 131;
    exp_33_ram[808] = 147;
    exp_33_ram[809] = 35;
    exp_33_ram[810] = 147;
    exp_33_ram[811] = 35;
    exp_33_ram[812] = 111;
    exp_33_ram[813] = 131;
    exp_33_ram[814] = 147;
    exp_33_ram[815] = 35;
    exp_33_ram[816] = 131;
    exp_33_ram[817] = 147;
    exp_33_ram[818] = 35;
    exp_33_ram[819] = 147;
    exp_33_ram[820] = 35;
    exp_33_ram[821] = 111;
    exp_33_ram[822] = 35;
    exp_33_ram[823] = 19;
    exp_33_ram[824] = 131;
    exp_33_ram[825] = 227;
    exp_33_ram[826] = 35;
    exp_33_ram[827] = 131;
    exp_33_ram[828] = 131;
    exp_33_ram[829] = 19;
    exp_33_ram[830] = 239;
    exp_33_ram[831] = 147;
    exp_33_ram[832] = 99;
    exp_33_ram[833] = 147;
    exp_33_ram[834] = 19;
    exp_33_ram[835] = 239;
    exp_33_ram[836] = 35;
    exp_33_ram[837] = 111;
    exp_33_ram[838] = 131;
    exp_33_ram[839] = 3;
    exp_33_ram[840] = 147;
    exp_33_ram[841] = 99;
    exp_33_ram[842] = 131;
    exp_33_ram[843] = 19;
    exp_33_ram[844] = 35;
    exp_33_ram[845] = 131;
    exp_33_ram[846] = 35;
    exp_33_ram[847] = 131;
    exp_33_ram[848] = 99;
    exp_33_ram[849] = 131;
    exp_33_ram[850] = 147;
    exp_33_ram[851] = 35;
    exp_33_ram[852] = 131;
    exp_33_ram[853] = 179;
    exp_33_ram[854] = 35;
    exp_33_ram[855] = 111;
    exp_33_ram[856] = 131;
    exp_33_ram[857] = 35;
    exp_33_ram[858] = 131;
    exp_33_ram[859] = 147;
    exp_33_ram[860] = 35;
    exp_33_ram[861] = 35;
    exp_33_ram[862] = 131;
    exp_33_ram[863] = 3;
    exp_33_ram[864] = 147;
    exp_33_ram[865] = 99;
    exp_33_ram[866] = 131;
    exp_33_ram[867] = 147;
    exp_33_ram[868] = 35;
    exp_33_ram[869] = 131;
    exp_33_ram[870] = 147;
    exp_33_ram[871] = 35;
    exp_33_ram[872] = 131;
    exp_33_ram[873] = 131;
    exp_33_ram[874] = 19;
    exp_33_ram[875] = 239;
    exp_33_ram[876] = 147;
    exp_33_ram[877] = 99;
    exp_33_ram[878] = 147;
    exp_33_ram[879] = 19;
    exp_33_ram[880] = 239;
    exp_33_ram[881] = 35;
    exp_33_ram[882] = 111;
    exp_33_ram[883] = 131;
    exp_33_ram[884] = 3;
    exp_33_ram[885] = 147;
    exp_33_ram[886] = 99;
    exp_33_ram[887] = 131;
    exp_33_ram[888] = 19;
    exp_33_ram[889] = 35;
    exp_33_ram[890] = 131;
    exp_33_ram[891] = 35;
    exp_33_ram[892] = 131;
    exp_33_ram[893] = 99;
    exp_33_ram[894] = 147;
    exp_33_ram[895] = 35;
    exp_33_ram[896] = 131;
    exp_33_ram[897] = 147;
    exp_33_ram[898] = 35;
    exp_33_ram[899] = 131;
    exp_33_ram[900] = 131;
    exp_33_ram[901] = 147;
    exp_33_ram[902] = 19;
    exp_33_ram[903] = 99;
    exp_33_ram[904] = 19;
    exp_33_ram[905] = 183;
    exp_33_ram[906] = 147;
    exp_33_ram[907] = 179;
    exp_33_ram[908] = 131;
    exp_33_ram[909] = 103;
    exp_33_ram[910] = 131;
    exp_33_ram[911] = 147;
    exp_33_ram[912] = 35;
    exp_33_ram[913] = 131;
    exp_33_ram[914] = 147;
    exp_33_ram[915] = 35;
    exp_33_ram[916] = 131;
    exp_33_ram[917] = 3;
    exp_33_ram[918] = 147;
    exp_33_ram[919] = 99;
    exp_33_ram[920] = 131;
    exp_33_ram[921] = 147;
    exp_33_ram[922] = 35;
    exp_33_ram[923] = 131;
    exp_33_ram[924] = 147;
    exp_33_ram[925] = 35;
    exp_33_ram[926] = 111;
    exp_33_ram[927] = 131;
    exp_33_ram[928] = 147;
    exp_33_ram[929] = 35;
    exp_33_ram[930] = 131;
    exp_33_ram[931] = 147;
    exp_33_ram[932] = 35;
    exp_33_ram[933] = 131;
    exp_33_ram[934] = 3;
    exp_33_ram[935] = 147;
    exp_33_ram[936] = 99;
    exp_33_ram[937] = 131;
    exp_33_ram[938] = 147;
    exp_33_ram[939] = 35;
    exp_33_ram[940] = 131;
    exp_33_ram[941] = 147;
    exp_33_ram[942] = 35;
    exp_33_ram[943] = 111;
    exp_33_ram[944] = 131;
    exp_33_ram[945] = 147;
    exp_33_ram[946] = 35;
    exp_33_ram[947] = 131;
    exp_33_ram[948] = 147;
    exp_33_ram[949] = 35;
    exp_33_ram[950] = 111;
    exp_33_ram[951] = 131;
    exp_33_ram[952] = 147;
    exp_33_ram[953] = 35;
    exp_33_ram[954] = 131;
    exp_33_ram[955] = 147;
    exp_33_ram[956] = 35;
    exp_33_ram[957] = 111;
    exp_33_ram[958] = 131;
    exp_33_ram[959] = 147;
    exp_33_ram[960] = 35;
    exp_33_ram[961] = 131;
    exp_33_ram[962] = 147;
    exp_33_ram[963] = 35;
    exp_33_ram[964] = 111;
    exp_33_ram[965] = 19;
    exp_33_ram[966] = 111;
    exp_33_ram[967] = 19;
    exp_33_ram[968] = 111;
    exp_33_ram[969] = 19;
    exp_33_ram[970] = 131;
    exp_33_ram[971] = 131;
    exp_33_ram[972] = 147;
    exp_33_ram[973] = 19;
    exp_33_ram[974] = 99;
    exp_33_ram[975] = 19;
    exp_33_ram[976] = 183;
    exp_33_ram[977] = 147;
    exp_33_ram[978] = 179;
    exp_33_ram[979] = 131;
    exp_33_ram[980] = 103;
    exp_33_ram[981] = 131;
    exp_33_ram[982] = 3;
    exp_33_ram[983] = 147;
    exp_33_ram[984] = 99;
    exp_33_ram[985] = 131;
    exp_33_ram[986] = 3;
    exp_33_ram[987] = 147;
    exp_33_ram[988] = 99;
    exp_33_ram[989] = 147;
    exp_33_ram[990] = 35;
    exp_33_ram[991] = 111;
    exp_33_ram[992] = 131;
    exp_33_ram[993] = 3;
    exp_33_ram[994] = 147;
    exp_33_ram[995] = 99;
    exp_33_ram[996] = 147;
    exp_33_ram[997] = 35;
    exp_33_ram[998] = 111;
    exp_33_ram[999] = 131;
    exp_33_ram[1000] = 3;
    exp_33_ram[1001] = 147;
    exp_33_ram[1002] = 99;
    exp_33_ram[1003] = 147;
    exp_33_ram[1004] = 35;
    exp_33_ram[1005] = 111;
    exp_33_ram[1006] = 147;
    exp_33_ram[1007] = 35;
    exp_33_ram[1008] = 131;
    exp_33_ram[1009] = 147;
    exp_33_ram[1010] = 35;
    exp_33_ram[1011] = 131;
    exp_33_ram[1012] = 3;
    exp_33_ram[1013] = 147;
    exp_33_ram[1014] = 99;
    exp_33_ram[1015] = 131;
    exp_33_ram[1016] = 147;
    exp_33_ram[1017] = 35;
    exp_33_ram[1018] = 131;
    exp_33_ram[1019] = 3;
    exp_33_ram[1020] = 147;
    exp_33_ram[1021] = 99;
    exp_33_ram[1022] = 131;
    exp_33_ram[1023] = 3;
    exp_33_ram[1024] = 147;
    exp_33_ram[1025] = 99;
    exp_33_ram[1026] = 131;
    exp_33_ram[1027] = 147;
    exp_33_ram[1028] = 35;
    exp_33_ram[1029] = 131;
    exp_33_ram[1030] = 147;
    exp_33_ram[1031] = 99;
    exp_33_ram[1032] = 131;
    exp_33_ram[1033] = 147;
    exp_33_ram[1034] = 35;
    exp_33_ram[1035] = 131;
    exp_33_ram[1036] = 3;
    exp_33_ram[1037] = 147;
    exp_33_ram[1038] = 99;
    exp_33_ram[1039] = 131;
    exp_33_ram[1040] = 3;
    exp_33_ram[1041] = 147;
    exp_33_ram[1042] = 99;
    exp_33_ram[1043] = 131;
    exp_33_ram[1044] = 147;
    exp_33_ram[1045] = 99;
    exp_33_ram[1046] = 131;
    exp_33_ram[1047] = 147;
    exp_33_ram[1048] = 99;
    exp_33_ram[1049] = 131;
    exp_33_ram[1050] = 19;
    exp_33_ram[1051] = 35;
    exp_33_ram[1052] = 131;
    exp_33_ram[1053] = 35;
    exp_33_ram[1054] = 131;
    exp_33_ram[1055] = 19;
    exp_33_ram[1056] = 131;
    exp_33_ram[1057] = 179;
    exp_33_ram[1058] = 179;
    exp_33_ram[1059] = 147;
    exp_33_ram[1060] = 131;
    exp_33_ram[1061] = 147;
    exp_33_ram[1062] = 19;
    exp_33_ram[1063] = 131;
    exp_33_ram[1064] = 35;
    exp_33_ram[1065] = 131;
    exp_33_ram[1066] = 35;
    exp_33_ram[1067] = 131;
    exp_33_ram[1068] = 3;
    exp_33_ram[1069] = 147;
    exp_33_ram[1070] = 19;
    exp_33_ram[1071] = 131;
    exp_33_ram[1072] = 3;
    exp_33_ram[1073] = 131;
    exp_33_ram[1074] = 3;
    exp_33_ram[1075] = 239;
    exp_33_ram[1076] = 35;
    exp_33_ram[1077] = 111;
    exp_33_ram[1078] = 131;
    exp_33_ram[1079] = 147;
    exp_33_ram[1080] = 99;
    exp_33_ram[1081] = 131;
    exp_33_ram[1082] = 19;
    exp_33_ram[1083] = 35;
    exp_33_ram[1084] = 131;
    exp_33_ram[1085] = 147;
    exp_33_ram[1086] = 111;
    exp_33_ram[1087] = 131;
    exp_33_ram[1088] = 147;
    exp_33_ram[1089] = 99;
    exp_33_ram[1090] = 131;
    exp_33_ram[1091] = 19;
    exp_33_ram[1092] = 35;
    exp_33_ram[1093] = 131;
    exp_33_ram[1094] = 147;
    exp_33_ram[1095] = 147;
    exp_33_ram[1096] = 111;
    exp_33_ram[1097] = 131;
    exp_33_ram[1098] = 19;
    exp_33_ram[1099] = 35;
    exp_33_ram[1100] = 131;
    exp_33_ram[1101] = 35;
    exp_33_ram[1102] = 131;
    exp_33_ram[1103] = 19;
    exp_33_ram[1104] = 131;
    exp_33_ram[1105] = 179;
    exp_33_ram[1106] = 179;
    exp_33_ram[1107] = 147;
    exp_33_ram[1108] = 131;
    exp_33_ram[1109] = 147;
    exp_33_ram[1110] = 19;
    exp_33_ram[1111] = 131;
    exp_33_ram[1112] = 35;
    exp_33_ram[1113] = 131;
    exp_33_ram[1114] = 35;
    exp_33_ram[1115] = 131;
    exp_33_ram[1116] = 3;
    exp_33_ram[1117] = 147;
    exp_33_ram[1118] = 19;
    exp_33_ram[1119] = 131;
    exp_33_ram[1120] = 3;
    exp_33_ram[1121] = 131;
    exp_33_ram[1122] = 3;
    exp_33_ram[1123] = 239;
    exp_33_ram[1124] = 35;
    exp_33_ram[1125] = 111;
    exp_33_ram[1126] = 131;
    exp_33_ram[1127] = 147;
    exp_33_ram[1128] = 99;
    exp_33_ram[1129] = 131;
    exp_33_ram[1130] = 147;
    exp_33_ram[1131] = 99;
    exp_33_ram[1132] = 131;
    exp_33_ram[1133] = 19;
    exp_33_ram[1134] = 35;
    exp_33_ram[1135] = 3;
    exp_33_ram[1136] = 131;
    exp_33_ram[1137] = 35;
    exp_33_ram[1138] = 131;
    exp_33_ram[1139] = 35;
    exp_33_ram[1140] = 131;
    exp_33_ram[1141] = 3;
    exp_33_ram[1142] = 147;
    exp_33_ram[1143] = 131;
    exp_33_ram[1144] = 3;
    exp_33_ram[1145] = 131;
    exp_33_ram[1146] = 3;
    exp_33_ram[1147] = 239;
    exp_33_ram[1148] = 35;
    exp_33_ram[1149] = 111;
    exp_33_ram[1150] = 131;
    exp_33_ram[1151] = 147;
    exp_33_ram[1152] = 99;
    exp_33_ram[1153] = 131;
    exp_33_ram[1154] = 19;
    exp_33_ram[1155] = 35;
    exp_33_ram[1156] = 131;
    exp_33_ram[1157] = 147;
    exp_33_ram[1158] = 111;
    exp_33_ram[1159] = 131;
    exp_33_ram[1160] = 147;
    exp_33_ram[1161] = 99;
    exp_33_ram[1162] = 131;
    exp_33_ram[1163] = 19;
    exp_33_ram[1164] = 35;
    exp_33_ram[1165] = 131;
    exp_33_ram[1166] = 147;
    exp_33_ram[1167] = 147;
    exp_33_ram[1168] = 111;
    exp_33_ram[1169] = 131;
    exp_33_ram[1170] = 19;
    exp_33_ram[1171] = 35;
    exp_33_ram[1172] = 131;
    exp_33_ram[1173] = 35;
    exp_33_ram[1174] = 131;
    exp_33_ram[1175] = 35;
    exp_33_ram[1176] = 131;
    exp_33_ram[1177] = 35;
    exp_33_ram[1178] = 131;
    exp_33_ram[1179] = 3;
    exp_33_ram[1180] = 147;
    exp_33_ram[1181] = 3;
    exp_33_ram[1182] = 131;
    exp_33_ram[1183] = 3;
    exp_33_ram[1184] = 131;
    exp_33_ram[1185] = 3;
    exp_33_ram[1186] = 239;
    exp_33_ram[1187] = 35;
    exp_33_ram[1188] = 131;
    exp_33_ram[1189] = 147;
    exp_33_ram[1190] = 35;
    exp_33_ram[1191] = 111;
    exp_33_ram[1192] = 147;
    exp_33_ram[1193] = 35;
    exp_33_ram[1194] = 131;
    exp_33_ram[1195] = 147;
    exp_33_ram[1196] = 99;
    exp_33_ram[1197] = 111;
    exp_33_ram[1198] = 131;
    exp_33_ram[1199] = 19;
    exp_33_ram[1200] = 35;
    exp_33_ram[1201] = 3;
    exp_33_ram[1202] = 131;
    exp_33_ram[1203] = 19;
    exp_33_ram[1204] = 131;
    exp_33_ram[1205] = 19;
    exp_33_ram[1206] = 231;
    exp_33_ram[1207] = 131;
    exp_33_ram[1208] = 19;
    exp_33_ram[1209] = 35;
    exp_33_ram[1210] = 3;
    exp_33_ram[1211] = 227;
    exp_33_ram[1212] = 131;
    exp_33_ram[1213] = 19;
    exp_33_ram[1214] = 35;
    exp_33_ram[1215] = 131;
    exp_33_ram[1216] = 19;
    exp_33_ram[1217] = 131;
    exp_33_ram[1218] = 19;
    exp_33_ram[1219] = 35;
    exp_33_ram[1220] = 3;
    exp_33_ram[1221] = 131;
    exp_33_ram[1222] = 19;
    exp_33_ram[1223] = 131;
    exp_33_ram[1224] = 231;
    exp_33_ram[1225] = 131;
    exp_33_ram[1226] = 147;
    exp_33_ram[1227] = 99;
    exp_33_ram[1228] = 111;
    exp_33_ram[1229] = 131;
    exp_33_ram[1230] = 19;
    exp_33_ram[1231] = 35;
    exp_33_ram[1232] = 3;
    exp_33_ram[1233] = 131;
    exp_33_ram[1234] = 19;
    exp_33_ram[1235] = 131;
    exp_33_ram[1236] = 19;
    exp_33_ram[1237] = 231;
    exp_33_ram[1238] = 131;
    exp_33_ram[1239] = 19;
    exp_33_ram[1240] = 35;
    exp_33_ram[1241] = 3;
    exp_33_ram[1242] = 227;
    exp_33_ram[1243] = 131;
    exp_33_ram[1244] = 147;
    exp_33_ram[1245] = 35;
    exp_33_ram[1246] = 111;
    exp_33_ram[1247] = 131;
    exp_33_ram[1248] = 19;
    exp_33_ram[1249] = 35;
    exp_33_ram[1250] = 131;
    exp_33_ram[1251] = 35;
    exp_33_ram[1252] = 131;
    exp_33_ram[1253] = 99;
    exp_33_ram[1254] = 131;
    exp_33_ram[1255] = 111;
    exp_33_ram[1256] = 147;
    exp_33_ram[1257] = 147;
    exp_33_ram[1258] = 3;
    exp_33_ram[1259] = 239;
    exp_33_ram[1260] = 35;
    exp_33_ram[1261] = 131;
    exp_33_ram[1262] = 147;
    exp_33_ram[1263] = 99;
    exp_33_ram[1264] = 3;
    exp_33_ram[1265] = 131;
    exp_33_ram[1266] = 99;
    exp_33_ram[1267] = 147;
    exp_33_ram[1268] = 35;
    exp_33_ram[1269] = 131;
    exp_33_ram[1270] = 147;
    exp_33_ram[1271] = 99;
    exp_33_ram[1272] = 111;
    exp_33_ram[1273] = 131;
    exp_33_ram[1274] = 19;
    exp_33_ram[1275] = 35;
    exp_33_ram[1276] = 3;
    exp_33_ram[1277] = 131;
    exp_33_ram[1278] = 19;
    exp_33_ram[1279] = 131;
    exp_33_ram[1280] = 19;
    exp_33_ram[1281] = 231;
    exp_33_ram[1282] = 131;
    exp_33_ram[1283] = 19;
    exp_33_ram[1284] = 35;
    exp_33_ram[1285] = 3;
    exp_33_ram[1286] = 227;
    exp_33_ram[1287] = 111;
    exp_33_ram[1288] = 131;
    exp_33_ram[1289] = 19;
    exp_33_ram[1290] = 35;
    exp_33_ram[1291] = 3;
    exp_33_ram[1292] = 131;
    exp_33_ram[1293] = 19;
    exp_33_ram[1294] = 35;
    exp_33_ram[1295] = 3;
    exp_33_ram[1296] = 131;
    exp_33_ram[1297] = 19;
    exp_33_ram[1298] = 131;
    exp_33_ram[1299] = 231;
    exp_33_ram[1300] = 131;
    exp_33_ram[1301] = 131;
    exp_33_ram[1302] = 99;
    exp_33_ram[1303] = 131;
    exp_33_ram[1304] = 147;
    exp_33_ram[1305] = 227;
    exp_33_ram[1306] = 131;
    exp_33_ram[1307] = 19;
    exp_33_ram[1308] = 35;
    exp_33_ram[1309] = 227;
    exp_33_ram[1310] = 131;
    exp_33_ram[1311] = 147;
    exp_33_ram[1312] = 99;
    exp_33_ram[1313] = 111;
    exp_33_ram[1314] = 131;
    exp_33_ram[1315] = 19;
    exp_33_ram[1316] = 35;
    exp_33_ram[1317] = 3;
    exp_33_ram[1318] = 131;
    exp_33_ram[1319] = 19;
    exp_33_ram[1320] = 131;
    exp_33_ram[1321] = 19;
    exp_33_ram[1322] = 231;
    exp_33_ram[1323] = 131;
    exp_33_ram[1324] = 19;
    exp_33_ram[1325] = 35;
    exp_33_ram[1326] = 3;
    exp_33_ram[1327] = 227;
    exp_33_ram[1328] = 131;
    exp_33_ram[1329] = 147;
    exp_33_ram[1330] = 35;
    exp_33_ram[1331] = 111;
    exp_33_ram[1332] = 147;
    exp_33_ram[1333] = 35;
    exp_33_ram[1334] = 131;
    exp_33_ram[1335] = 147;
    exp_33_ram[1336] = 35;
    exp_33_ram[1337] = 131;
    exp_33_ram[1338] = 19;
    exp_33_ram[1339] = 35;
    exp_33_ram[1340] = 131;
    exp_33_ram[1341] = 19;
    exp_33_ram[1342] = 131;
    exp_33_ram[1343] = 35;
    exp_33_ram[1344] = 131;
    exp_33_ram[1345] = 35;
    exp_33_ram[1346] = 131;
    exp_33_ram[1347] = 19;
    exp_33_ram[1348] = 147;
    exp_33_ram[1349] = 131;
    exp_33_ram[1350] = 3;
    exp_33_ram[1351] = 131;
    exp_33_ram[1352] = 3;
    exp_33_ram[1353] = 239;
    exp_33_ram[1354] = 35;
    exp_33_ram[1355] = 131;
    exp_33_ram[1356] = 147;
    exp_33_ram[1357] = 35;
    exp_33_ram[1358] = 111;
    exp_33_ram[1359] = 131;
    exp_33_ram[1360] = 19;
    exp_33_ram[1361] = 35;
    exp_33_ram[1362] = 3;
    exp_33_ram[1363] = 131;
    exp_33_ram[1364] = 19;
    exp_33_ram[1365] = 131;
    exp_33_ram[1366] = 19;
    exp_33_ram[1367] = 231;
    exp_33_ram[1368] = 131;
    exp_33_ram[1369] = 147;
    exp_33_ram[1370] = 35;
    exp_33_ram[1371] = 111;
    exp_33_ram[1372] = 131;
    exp_33_ram[1373] = 3;
    exp_33_ram[1374] = 131;
    exp_33_ram[1375] = 19;
    exp_33_ram[1376] = 35;
    exp_33_ram[1377] = 3;
    exp_33_ram[1378] = 131;
    exp_33_ram[1379] = 19;
    exp_33_ram[1380] = 131;
    exp_33_ram[1381] = 231;
    exp_33_ram[1382] = 131;
    exp_33_ram[1383] = 147;
    exp_33_ram[1384] = 35;
    exp_33_ram[1385] = 19;
    exp_33_ram[1386] = 131;
    exp_33_ram[1387] = 131;
    exp_33_ram[1388] = 99;
    exp_33_ram[1389] = 3;
    exp_33_ram[1390] = 131;
    exp_33_ram[1391] = 99;
    exp_33_ram[1392] = 131;
    exp_33_ram[1393] = 147;
    exp_33_ram[1394] = 111;
    exp_33_ram[1395] = 131;
    exp_33_ram[1396] = 3;
    exp_33_ram[1397] = 131;
    exp_33_ram[1398] = 19;
    exp_33_ram[1399] = 131;
    exp_33_ram[1400] = 19;
    exp_33_ram[1401] = 231;
    exp_33_ram[1402] = 131;
    exp_33_ram[1403] = 19;
    exp_33_ram[1404] = 131;
    exp_33_ram[1405] = 3;
    exp_33_ram[1406] = 19;
    exp_33_ram[1407] = 103;
    exp_33_ram[1408] = 19;
    exp_33_ram[1409] = 35;
    exp_33_ram[1410] = 35;
    exp_33_ram[1411] = 19;
    exp_33_ram[1412] = 35;
    exp_33_ram[1413] = 35;
    exp_33_ram[1414] = 35;
    exp_33_ram[1415] = 35;
    exp_33_ram[1416] = 35;
    exp_33_ram[1417] = 35;
    exp_33_ram[1418] = 35;
    exp_33_ram[1419] = 35;
    exp_33_ram[1420] = 147;
    exp_33_ram[1421] = 35;
    exp_33_ram[1422] = 131;
    exp_33_ram[1423] = 147;
    exp_33_ram[1424] = 35;
    exp_33_ram[1425] = 3;
    exp_33_ram[1426] = 147;
    exp_33_ram[1427] = 131;
    exp_33_ram[1428] = 19;
    exp_33_ram[1429] = 147;
    exp_33_ram[1430] = 19;
    exp_33_ram[1431] = 239;
    exp_33_ram[1432] = 35;
    exp_33_ram[1433] = 131;
    exp_33_ram[1434] = 19;
    exp_33_ram[1435] = 131;
    exp_33_ram[1436] = 3;
    exp_33_ram[1437] = 19;
    exp_33_ram[1438] = 103;
    exp_33_ram[1439] = 19;
    exp_33_ram[1440] = 35;
    exp_33_ram[1441] = 35;
    exp_33_ram[1442] = 19;
    exp_33_ram[1443] = 147;
    exp_33_ram[1444] = 163;
    exp_33_ram[1445] = 3;
    exp_33_ram[1446] = 183;
    exp_33_ram[1447] = 131;
    exp_33_ram[1448] = 147;
    exp_33_ram[1449] = 19;
    exp_33_ram[1450] = 239;
    exp_33_ram[1451] = 19;
    exp_33_ram[1452] = 131;
    exp_33_ram[1453] = 3;
    exp_33_ram[1454] = 19;
    exp_33_ram[1455] = 103;
    exp_33_ram[1456] = 19;
    exp_33_ram[1457] = 35;
    exp_33_ram[1458] = 35;
    exp_33_ram[1459] = 19;
    exp_33_ram[1460] = 19;
    exp_33_ram[1461] = 239;
    exp_33_ram[1462] = 3;
    exp_33_ram[1463] = 131;
    exp_33_ram[1464] = 19;
    exp_33_ram[1465] = 147;
    exp_33_ram[1466] = 19;
    exp_33_ram[1467] = 239;
    exp_33_ram[1468] = 3;
    exp_33_ram[1469] = 131;
    exp_33_ram[1470] = 19;
    exp_33_ram[1471] = 147;
    exp_33_ram[1472] = 19;
    exp_33_ram[1473] = 239;
    exp_33_ram[1474] = 3;
    exp_33_ram[1475] = 131;
    exp_33_ram[1476] = 19;
    exp_33_ram[1477] = 147;
    exp_33_ram[1478] = 19;
    exp_33_ram[1479] = 239;
    exp_33_ram[1480] = 3;
    exp_33_ram[1481] = 131;
    exp_33_ram[1482] = 19;
    exp_33_ram[1483] = 147;
    exp_33_ram[1484] = 19;
    exp_33_ram[1485] = 239;
    exp_33_ram[1486] = 3;
    exp_33_ram[1487] = 131;
    exp_33_ram[1488] = 19;
    exp_33_ram[1489] = 147;
    exp_33_ram[1490] = 19;
    exp_33_ram[1491] = 239;
    exp_33_ram[1492] = 3;
    exp_33_ram[1493] = 131;
    exp_33_ram[1494] = 19;
    exp_33_ram[1495] = 147;
    exp_33_ram[1496] = 19;
    exp_33_ram[1497] = 239;
    exp_33_ram[1498] = 19;
    exp_33_ram[1499] = 147;
    exp_33_ram[1500] = 19;
    exp_33_ram[1501] = 239;
    exp_33_ram[1502] = 3;
    exp_33_ram[1503] = 131;
    exp_33_ram[1504] = 19;
    exp_33_ram[1505] = 147;
    exp_33_ram[1506] = 19;
    exp_33_ram[1507] = 239;
    exp_33_ram[1508] = 3;
    exp_33_ram[1509] = 131;
    exp_33_ram[1510] = 19;
    exp_33_ram[1511] = 147;
    exp_33_ram[1512] = 19;
    exp_33_ram[1513] = 239;
    exp_33_ram[1514] = 3;
    exp_33_ram[1515] = 131;
    exp_33_ram[1516] = 19;
    exp_33_ram[1517] = 147;
    exp_33_ram[1518] = 19;
    exp_33_ram[1519] = 239;
    exp_33_ram[1520] = 3;
    exp_33_ram[1521] = 131;
    exp_33_ram[1522] = 19;
    exp_33_ram[1523] = 147;
    exp_33_ram[1524] = 19;
    exp_33_ram[1525] = 239;
    exp_33_ram[1526] = 3;
    exp_33_ram[1527] = 131;
    exp_33_ram[1528] = 19;
    exp_33_ram[1529] = 147;
    exp_33_ram[1530] = 19;
    exp_33_ram[1531] = 239;
    exp_33_ram[1532] = 3;
    exp_33_ram[1533] = 131;
    exp_33_ram[1534] = 19;
    exp_33_ram[1535] = 147;
    exp_33_ram[1536] = 19;
    exp_33_ram[1537] = 239;
    exp_33_ram[1538] = 3;
    exp_33_ram[1539] = 131;
    exp_33_ram[1540] = 19;
    exp_33_ram[1541] = 147;
    exp_33_ram[1542] = 19;
    exp_33_ram[1543] = 239;
    exp_33_ram[1544] = 3;
    exp_33_ram[1545] = 131;
    exp_33_ram[1546] = 19;
    exp_33_ram[1547] = 147;
    exp_33_ram[1548] = 19;
    exp_33_ram[1549] = 239;
    exp_33_ram[1550] = 3;
    exp_33_ram[1551] = 131;
    exp_33_ram[1552] = 19;
    exp_33_ram[1553] = 147;
    exp_33_ram[1554] = 19;
    exp_33_ram[1555] = 239;
    exp_33_ram[1556] = 3;
    exp_33_ram[1557] = 131;
    exp_33_ram[1558] = 19;
    exp_33_ram[1559] = 147;
    exp_33_ram[1560] = 19;
    exp_33_ram[1561] = 239;
    exp_33_ram[1562] = 3;
    exp_33_ram[1563] = 131;
    exp_33_ram[1564] = 19;
    exp_33_ram[1565] = 147;
    exp_33_ram[1566] = 19;
    exp_33_ram[1567] = 239;
    exp_33_ram[1568] = 3;
    exp_33_ram[1569] = 131;
    exp_33_ram[1570] = 19;
    exp_33_ram[1571] = 147;
    exp_33_ram[1572] = 19;
    exp_33_ram[1573] = 239;
    exp_33_ram[1574] = 19;
    exp_33_ram[1575] = 147;
    exp_33_ram[1576] = 19;
    exp_33_ram[1577] = 239;
    exp_33_ram[1578] = 3;
    exp_33_ram[1579] = 131;
    exp_33_ram[1580] = 19;
    exp_33_ram[1581] = 147;
    exp_33_ram[1582] = 19;
    exp_33_ram[1583] = 239;
    exp_33_ram[1584] = 3;
    exp_33_ram[1585] = 131;
    exp_33_ram[1586] = 19;
    exp_33_ram[1587] = 147;
    exp_33_ram[1588] = 19;
    exp_33_ram[1589] = 239;
    exp_33_ram[1590] = 3;
    exp_33_ram[1591] = 131;
    exp_33_ram[1592] = 19;
    exp_33_ram[1593] = 147;
    exp_33_ram[1594] = 19;
    exp_33_ram[1595] = 239;
    exp_33_ram[1596] = 3;
    exp_33_ram[1597] = 131;
    exp_33_ram[1598] = 19;
    exp_33_ram[1599] = 147;
    exp_33_ram[1600] = 19;
    exp_33_ram[1601] = 239;
    exp_33_ram[1602] = 3;
    exp_33_ram[1603] = 131;
    exp_33_ram[1604] = 19;
    exp_33_ram[1605] = 147;
    exp_33_ram[1606] = 19;
    exp_33_ram[1607] = 239;
    exp_33_ram[1608] = 3;
    exp_33_ram[1609] = 131;
    exp_33_ram[1610] = 19;
    exp_33_ram[1611] = 147;
    exp_33_ram[1612] = 19;
    exp_33_ram[1613] = 239;
    exp_33_ram[1614] = 3;
    exp_33_ram[1615] = 131;
    exp_33_ram[1616] = 19;
    exp_33_ram[1617] = 147;
    exp_33_ram[1618] = 19;
    exp_33_ram[1619] = 239;
    exp_33_ram[1620] = 3;
    exp_33_ram[1621] = 131;
    exp_33_ram[1622] = 19;
    exp_33_ram[1623] = 147;
    exp_33_ram[1624] = 19;
    exp_33_ram[1625] = 239;
    exp_33_ram[1626] = 3;
    exp_33_ram[1627] = 131;
    exp_33_ram[1628] = 19;
    exp_33_ram[1629] = 147;
    exp_33_ram[1630] = 19;
    exp_33_ram[1631] = 239;
    exp_33_ram[1632] = 3;
    exp_33_ram[1633] = 131;
    exp_33_ram[1634] = 19;
    exp_33_ram[1635] = 147;
    exp_33_ram[1636] = 19;
    exp_33_ram[1637] = 239;
    exp_33_ram[1638] = 3;
    exp_33_ram[1639] = 131;
    exp_33_ram[1640] = 19;
    exp_33_ram[1641] = 147;
    exp_33_ram[1642] = 19;
    exp_33_ram[1643] = 239;
    exp_33_ram[1644] = 3;
    exp_33_ram[1645] = 131;
    exp_33_ram[1646] = 19;
    exp_33_ram[1647] = 147;
    exp_33_ram[1648] = 19;
    exp_33_ram[1649] = 239;
    exp_33_ram[1650] = 19;
    exp_33_ram[1651] = 147;
    exp_33_ram[1652] = 19;
    exp_33_ram[1653] = 239;
    exp_33_ram[1654] = 3;
    exp_33_ram[1655] = 131;
    exp_33_ram[1656] = 19;
    exp_33_ram[1657] = 147;
    exp_33_ram[1658] = 19;
    exp_33_ram[1659] = 239;
    exp_33_ram[1660] = 3;
    exp_33_ram[1661] = 131;
    exp_33_ram[1662] = 19;
    exp_33_ram[1663] = 147;
    exp_33_ram[1664] = 19;
    exp_33_ram[1665] = 239;
    exp_33_ram[1666] = 3;
    exp_33_ram[1667] = 131;
    exp_33_ram[1668] = 19;
    exp_33_ram[1669] = 147;
    exp_33_ram[1670] = 19;
    exp_33_ram[1671] = 239;
    exp_33_ram[1672] = 3;
    exp_33_ram[1673] = 131;
    exp_33_ram[1674] = 19;
    exp_33_ram[1675] = 147;
    exp_33_ram[1676] = 19;
    exp_33_ram[1677] = 239;
    exp_33_ram[1678] = 3;
    exp_33_ram[1679] = 131;
    exp_33_ram[1680] = 19;
    exp_33_ram[1681] = 147;
    exp_33_ram[1682] = 19;
    exp_33_ram[1683] = 239;
    exp_33_ram[1684] = 3;
    exp_33_ram[1685] = 131;
    exp_33_ram[1686] = 19;
    exp_33_ram[1687] = 147;
    exp_33_ram[1688] = 19;
    exp_33_ram[1689] = 239;
    exp_33_ram[1690] = 3;
    exp_33_ram[1691] = 131;
    exp_33_ram[1692] = 19;
    exp_33_ram[1693] = 147;
    exp_33_ram[1694] = 19;
    exp_33_ram[1695] = 239;
    exp_33_ram[1696] = 3;
    exp_33_ram[1697] = 131;
    exp_33_ram[1698] = 19;
    exp_33_ram[1699] = 147;
    exp_33_ram[1700] = 19;
    exp_33_ram[1701] = 239;
    exp_33_ram[1702] = 3;
    exp_33_ram[1703] = 131;
    exp_33_ram[1704] = 19;
    exp_33_ram[1705] = 147;
    exp_33_ram[1706] = 19;
    exp_33_ram[1707] = 239;
    exp_33_ram[1708] = 3;
    exp_33_ram[1709] = 131;
    exp_33_ram[1710] = 19;
    exp_33_ram[1711] = 147;
    exp_33_ram[1712] = 19;
    exp_33_ram[1713] = 239;
    exp_33_ram[1714] = 3;
    exp_33_ram[1715] = 131;
    exp_33_ram[1716] = 19;
    exp_33_ram[1717] = 147;
    exp_33_ram[1718] = 19;
    exp_33_ram[1719] = 239;
    exp_33_ram[1720] = 3;
    exp_33_ram[1721] = 131;
    exp_33_ram[1722] = 19;
    exp_33_ram[1723] = 147;
    exp_33_ram[1724] = 19;
    exp_33_ram[1725] = 239;
    exp_33_ram[1726] = 19;
    exp_33_ram[1727] = 147;
    exp_33_ram[1728] = 19;
    exp_33_ram[1729] = 239;
    exp_33_ram[1730] = 3;
    exp_33_ram[1731] = 131;
    exp_33_ram[1732] = 19;
    exp_33_ram[1733] = 147;
    exp_33_ram[1734] = 19;
    exp_33_ram[1735] = 239;
    exp_33_ram[1736] = 3;
    exp_33_ram[1737] = 131;
    exp_33_ram[1738] = 19;
    exp_33_ram[1739] = 147;
    exp_33_ram[1740] = 19;
    exp_33_ram[1741] = 239;
    exp_33_ram[1742] = 3;
    exp_33_ram[1743] = 131;
    exp_33_ram[1744] = 19;
    exp_33_ram[1745] = 147;
    exp_33_ram[1746] = 19;
    exp_33_ram[1747] = 239;
    exp_33_ram[1748] = 3;
    exp_33_ram[1749] = 131;
    exp_33_ram[1750] = 19;
    exp_33_ram[1751] = 147;
    exp_33_ram[1752] = 19;
    exp_33_ram[1753] = 239;
    exp_33_ram[1754] = 3;
    exp_33_ram[1755] = 131;
    exp_33_ram[1756] = 19;
    exp_33_ram[1757] = 147;
    exp_33_ram[1758] = 19;
    exp_33_ram[1759] = 239;
    exp_33_ram[1760] = 3;
    exp_33_ram[1761] = 131;
    exp_33_ram[1762] = 19;
    exp_33_ram[1763] = 147;
    exp_33_ram[1764] = 19;
    exp_33_ram[1765] = 239;
    exp_33_ram[1766] = 3;
    exp_33_ram[1767] = 131;
    exp_33_ram[1768] = 19;
    exp_33_ram[1769] = 147;
    exp_33_ram[1770] = 19;
    exp_33_ram[1771] = 239;
    exp_33_ram[1772] = 3;
    exp_33_ram[1773] = 131;
    exp_33_ram[1774] = 19;
    exp_33_ram[1775] = 147;
    exp_33_ram[1776] = 19;
    exp_33_ram[1777] = 239;
    exp_33_ram[1778] = 3;
    exp_33_ram[1779] = 131;
    exp_33_ram[1780] = 19;
    exp_33_ram[1781] = 147;
    exp_33_ram[1782] = 19;
    exp_33_ram[1783] = 239;
    exp_33_ram[1784] = 3;
    exp_33_ram[1785] = 131;
    exp_33_ram[1786] = 19;
    exp_33_ram[1787] = 147;
    exp_33_ram[1788] = 19;
    exp_33_ram[1789] = 239;
    exp_33_ram[1790] = 3;
    exp_33_ram[1791] = 131;
    exp_33_ram[1792] = 19;
    exp_33_ram[1793] = 147;
    exp_33_ram[1794] = 19;
    exp_33_ram[1795] = 239;
    exp_33_ram[1796] = 3;
    exp_33_ram[1797] = 131;
    exp_33_ram[1798] = 19;
    exp_33_ram[1799] = 147;
    exp_33_ram[1800] = 19;
    exp_33_ram[1801] = 239;
    exp_33_ram[1802] = 3;
    exp_33_ram[1803] = 131;
    exp_33_ram[1804] = 19;
    exp_33_ram[1805] = 147;
    exp_33_ram[1806] = 19;
    exp_33_ram[1807] = 239;
    exp_33_ram[1808] = 3;
    exp_33_ram[1809] = 131;
    exp_33_ram[1810] = 19;
    exp_33_ram[1811] = 147;
    exp_33_ram[1812] = 19;
    exp_33_ram[1813] = 239;
    exp_33_ram[1814] = 3;
    exp_33_ram[1815] = 131;
    exp_33_ram[1816] = 19;
    exp_33_ram[1817] = 147;
    exp_33_ram[1818] = 19;
    exp_33_ram[1819] = 239;
    exp_33_ram[1820] = 3;
    exp_33_ram[1821] = 131;
    exp_33_ram[1822] = 19;
    exp_33_ram[1823] = 147;
    exp_33_ram[1824] = 19;
    exp_33_ram[1825] = 239;
    exp_33_ram[1826] = 3;
    exp_33_ram[1827] = 131;
    exp_33_ram[1828] = 19;
    exp_33_ram[1829] = 147;
    exp_33_ram[1830] = 19;
    exp_33_ram[1831] = 239;
    exp_33_ram[1832] = 3;
    exp_33_ram[1833] = 131;
    exp_33_ram[1834] = 19;
    exp_33_ram[1835] = 147;
    exp_33_ram[1836] = 19;
    exp_33_ram[1837] = 239;
    exp_33_ram[1838] = 3;
    exp_33_ram[1839] = 131;
    exp_33_ram[1840] = 19;
    exp_33_ram[1841] = 147;
    exp_33_ram[1842] = 19;
    exp_33_ram[1843] = 239;
    exp_33_ram[1844] = 3;
    exp_33_ram[1845] = 131;
    exp_33_ram[1846] = 19;
    exp_33_ram[1847] = 147;
    exp_33_ram[1848] = 19;
    exp_33_ram[1849] = 239;
    exp_33_ram[1850] = 3;
    exp_33_ram[1851] = 131;
    exp_33_ram[1852] = 19;
    exp_33_ram[1853] = 147;
    exp_33_ram[1854] = 19;
    exp_33_ram[1855] = 239;
    exp_33_ram[1856] = 3;
    exp_33_ram[1857] = 131;
    exp_33_ram[1858] = 19;
    exp_33_ram[1859] = 147;
    exp_33_ram[1860] = 19;
    exp_33_ram[1861] = 239;
    exp_33_ram[1862] = 3;
    exp_33_ram[1863] = 131;
    exp_33_ram[1864] = 19;
    exp_33_ram[1865] = 147;
    exp_33_ram[1866] = 19;
    exp_33_ram[1867] = 239;
    exp_33_ram[1868] = 3;
    exp_33_ram[1869] = 131;
    exp_33_ram[1870] = 19;
    exp_33_ram[1871] = 147;
    exp_33_ram[1872] = 19;
    exp_33_ram[1873] = 239;
    exp_33_ram[1874] = 3;
    exp_33_ram[1875] = 131;
    exp_33_ram[1876] = 19;
    exp_33_ram[1877] = 147;
    exp_33_ram[1878] = 19;
    exp_33_ram[1879] = 239;
    exp_33_ram[1880] = 3;
    exp_33_ram[1881] = 131;
    exp_33_ram[1882] = 19;
    exp_33_ram[1883] = 147;
    exp_33_ram[1884] = 19;
    exp_33_ram[1885] = 239;
    exp_33_ram[1886] = 19;
    exp_33_ram[1887] = 239;
    exp_33_ram[1888] = 19;
    exp_33_ram[1889] = 131;
    exp_33_ram[1890] = 3;
    exp_33_ram[1891] = 19;
    exp_33_ram[1892] = 103;
    exp_33_ram[1893] = 19;
    exp_33_ram[1894] = 35;
    exp_33_ram[1895] = 35;
    exp_33_ram[1896] = 19;
    exp_33_ram[1897] = 239;
    exp_33_ram[1898] = 19;
    exp_33_ram[1899] = 131;
    exp_33_ram[1900] = 3;
    exp_33_ram[1901] = 19;
    exp_33_ram[1902] = 103;
    exp_33_ram[1903] = 8;
    exp_33_ram[1904] = 144;
    exp_33_ram[1905] = 216;
    exp_33_ram[1906] = 216;
    exp_33_ram[1907] = 180;
    exp_33_ram[1908] = 216;
    exp_33_ram[1909] = 216;
    exp_33_ram[1910] = 216;
    exp_33_ram[1911] = 216;
    exp_33_ram[1912] = 216;
    exp_33_ram[1913] = 216;
    exp_33_ram[1914] = 216;
    exp_33_ram[1915] = 108;
    exp_33_ram[1916] = 216;
    exp_33_ram[1917] = 72;
    exp_33_ram[1918] = 216;
    exp_33_ram[1919] = 216;
    exp_33_ram[1920] = 36;
    exp_33_ram[1921] = 124;
    exp_33_ram[1922] = 20;
    exp_33_ram[1923] = 220;
    exp_33_ram[1924] = 20;
    exp_33_ram[1925] = 56;
    exp_33_ram[1926] = 20;
    exp_33_ram[1927] = 20;
    exp_33_ram[1928] = 20;
    exp_33_ram[1929] = 20;
    exp_33_ram[1930] = 20;
    exp_33_ram[1931] = 20;
    exp_33_ram[1932] = 20;
    exp_33_ram[1933] = 192;
    exp_33_ram[1934] = 20;
    exp_33_ram[1935] = 20;
    exp_33_ram[1936] = 20;
    exp_33_ram[1937] = 20;
    exp_33_ram[1938] = 20;
    exp_33_ram[1939] = 248;
    exp_33_ram[1940] = 60;
    exp_33_ram[1941] = 112;
    exp_33_ram[1942] = 112;
    exp_33_ram[1943] = 112;
    exp_33_ram[1944] = 112;
    exp_33_ram[1945] = 112;
    exp_33_ram[1946] = 112;
    exp_33_ram[1947] = 112;
    exp_33_ram[1948] = 112;
    exp_33_ram[1949] = 112;
    exp_33_ram[1950] = 112;
    exp_33_ram[1951] = 112;
    exp_33_ram[1952] = 112;
    exp_33_ram[1953] = 112;
    exp_33_ram[1954] = 112;
    exp_33_ram[1955] = 112;
    exp_33_ram[1956] = 112;
    exp_33_ram[1957] = 112;
    exp_33_ram[1958] = 112;
    exp_33_ram[1959] = 112;
    exp_33_ram[1960] = 112;
    exp_33_ram[1961] = 112;
    exp_33_ram[1962] = 112;
    exp_33_ram[1963] = 112;
    exp_33_ram[1964] = 112;
    exp_33_ram[1965] = 112;
    exp_33_ram[1966] = 112;
    exp_33_ram[1967] = 112;
    exp_33_ram[1968] = 112;
    exp_33_ram[1969] = 112;
    exp_33_ram[1970] = 112;
    exp_33_ram[1971] = 112;
    exp_33_ram[1972] = 112;
    exp_33_ram[1973] = 112;
    exp_33_ram[1974] = 112;
    exp_33_ram[1975] = 112;
    exp_33_ram[1976] = 112;
    exp_33_ram[1977] = 112;
    exp_33_ram[1978] = 112;
    exp_33_ram[1979] = 112;
    exp_33_ram[1980] = 112;
    exp_33_ram[1981] = 112;
    exp_33_ram[1982] = 112;
    exp_33_ram[1983] = 112;
    exp_33_ram[1984] = 112;
    exp_33_ram[1985] = 112;
    exp_33_ram[1986] = 112;
    exp_33_ram[1987] = 112;
    exp_33_ram[1988] = 112;
    exp_33_ram[1989] = 112;
    exp_33_ram[1990] = 112;
    exp_33_ram[1991] = 84;
    exp_33_ram[1992] = 112;
    exp_33_ram[1993] = 112;
    exp_33_ram[1994] = 112;
    exp_33_ram[1995] = 112;
    exp_33_ram[1996] = 112;
    exp_33_ram[1997] = 112;
    exp_33_ram[1998] = 112;
    exp_33_ram[1999] = 112;
    exp_33_ram[2000] = 112;
    exp_33_ram[2001] = 84;
    exp_33_ram[2002] = 160;
    exp_33_ram[2003] = 84;
    exp_33_ram[2004] = 112;
    exp_33_ram[2005] = 112;
    exp_33_ram[2006] = 112;
    exp_33_ram[2007] = 112;
    exp_33_ram[2008] = 84;
    exp_33_ram[2009] = 112;
    exp_33_ram[2010] = 112;
    exp_33_ram[2011] = 112;
    exp_33_ram[2012] = 112;
    exp_33_ram[2013] = 112;
    exp_33_ram[2014] = 84;
    exp_33_ram[2015] = 208;
    exp_33_ram[2016] = 112;
    exp_33_ram[2017] = 112;
    exp_33_ram[2018] = 124;
    exp_33_ram[2019] = 112;
    exp_33_ram[2020] = 84;
    exp_33_ram[2021] = 112;
    exp_33_ram[2022] = 112;
    exp_33_ram[2023] = 84;
    exp_33_ram[2024] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_179;

  reg [31:0] exp_179_reg;
  always@(*) begin
    case (exp_177)
      0:exp_179_reg <= exp_157;
      1:exp_179_reg <= exp_167;
      default:exp_179_reg <= exp_178;
    endcase
  end
  assign exp_179 = exp_179_reg;
  assign exp_177 = exp_139[2:2];
  assign exp_139 = exp_1;
  assign exp_178 = 0;

      reg [31:0] exp_157_reg = 0;
      always@(posedge clk) begin
        if (exp_156) begin
          exp_157_reg <= exp_164;
        end
      end
      assign exp_157 = exp_157_reg;
    
  reg [31:0] exp_164_reg;
  always@(*) begin
    case (exp_159)
      0:exp_164_reg <= exp_161;
      1:exp_164_reg <= exp_162;
      default:exp_164_reg <= exp_163;
    endcase
  end
  assign exp_164 = exp_164_reg;
  assign exp_159 = exp_157 == exp_158;
  assign exp_158 = 4294967295;
  assign exp_163 = 0;
  assign exp_161 = exp_157 + exp_160;
  assign exp_160 = 1;
  assign exp_162 = 0;
  assign exp_156 = 1;

      reg [31:0] exp_167_reg = 0;
      always@(posedge clk) begin
        if (exp_166) begin
          exp_167_reg <= exp_174;
        end
      end
      assign exp_167 = exp_167_reg;
    
  reg [31:0] exp_174_reg;
  always@(*) begin
    case (exp_169)
      0:exp_174_reg <= exp_171;
      1:exp_174_reg <= exp_172;
      default:exp_174_reg <= exp_173;
    endcase
  end
  assign exp_174 = exp_174_reg;
  assign exp_169 = exp_167 == exp_168;
  assign exp_168 = 4294967295;
  assign exp_173 = 0;
  assign exp_171 = exp_167 + exp_170;
  assign exp_170 = 1;
  assign exp_172 = 0;
  assign exp_166 = exp_159 & exp_165;
  assign exp_165 = 1;
  assign exp_182 = exp_201;
  assign exp_201 = 0;
  assign exp_204 = exp_222;
  assign exp_222 = 0;
  assign exp_226 = exp_241;
  assign exp_241 = stdin_in;
  assign exp_461 = exp_248[15:8];
  assign exp_462 = exp_248[23:16];
  assign exp_463 = exp_248[31:24];
  assign exp_475 = $signed(exp_474);
  assign exp_474 = exp_473 + exp_469;
  assign exp_473 = 0;

  reg [15:0] exp_469_reg;
  always@(*) begin
    case (exp_459)
      0:exp_469_reg <= exp_466;
      1:exp_469_reg <= exp_467;
      default:exp_469_reg <= exp_468;
    endcase
  end
  assign exp_469 = exp_469_reg;
  assign exp_468 = 0;
  assign exp_466 = exp_248[15:0];
  assign exp_467 = exp_248[31:16];
  assign exp_476 = 0;
  assign exp_477 = exp_465;
  assign exp_478 = exp_469;
  assign exp_479 = 0;
  assign exp_480 = 0;

  reg [31:0] exp_839_reg;
  always@(*) begin
    case (exp_629)
      0:exp_839_reg <= exp_835;
      1:exp_839_reg <= exp_837;
      default:exp_839_reg <= exp_838;
    endcase
  end
  assign exp_839 = exp_839_reg;
  assign exp_838 = 0;

  reg [31:0] exp_835_reg;
  always@(*) begin
    case (exp_606)
      0:exp_835_reg <= exp_830;
      1:exp_835_reg <= exp_831;
      default:exp_835_reg <= exp_834;
    endcase
  end
  assign exp_835 = exp_835_reg;
  assign exp_606 = exp_605 & exp_603;
  assign exp_605 = exp_598 == exp_604;
  assign exp_604 = 0;
  assign exp_834 = 0;
  assign exp_830 = exp_829[63:32];

  reg [63:0] exp_829_reg;
  always@(*) begin
    case (exp_826)
      0:exp_829_reg <= exp_825;
      1:exp_829_reg <= exp_827;
      default:exp_829_reg <= exp_828;
    endcase
  end
  assign exp_829 = exp_829_reg;

      reg [0:0] exp_826_reg = 0;
      always@(posedge clk) begin
        if (exp_811) begin
          exp_826_reg <= exp_809;
        end
      end
      assign exp_826 = exp_826_reg;
    
      reg [0:0] exp_809_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_809_reg <= exp_786;
        end
      end
      assign exp_809 = exp_809_reg;
    
      reg [0:0] exp_786_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_786_reg <= exp_783;
        end
      end
      assign exp_786 = exp_786_reg;
      assign exp_783 = exp_781 ^ exp_782;
  assign exp_781 = exp_763 & exp_746;
  assign exp_763 = exp_762 + exp_761;
  assign exp_762 = 0;
  assign exp_761 = exp_759[31:31];

      reg [31:0] exp_759_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_759_reg <= exp_376;
        end
      end
      assign exp_759 = exp_759_reg;
      assign exp_758 = exp_748 == exp_757;
  assign exp_757 = 0;
  assign exp_746 = exp_745 | exp_612;
  assign exp_745 = exp_606 | exp_609;
  assign exp_609 = exp_608 & exp_603;
  assign exp_608 = exp_598 == exp_607;
  assign exp_607 = 1;
  assign exp_612 = exp_611 & exp_603;
  assign exp_611 = exp_598 == exp_610;
  assign exp_610 = 2;
  assign exp_782 = exp_766 & exp_747;
  assign exp_766 = exp_765 + exp_764;
  assign exp_765 = 0;
  assign exp_764 = exp_760[31:31];

      reg [31:0] exp_760_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_760_reg <= exp_377;
        end
      end
      assign exp_760 = exp_760_reg;
      assign exp_747 = exp_606 | exp_609;
  assign exp_768 = exp_748 == exp_767;
  assign exp_767 = 1;
  assign exp_788 = exp_748 == exp_787;
  assign exp_787 = 2;
  assign exp_811 = exp_748 == exp_810;
  assign exp_810 = 3;
  assign exp_828 = 0;

      reg [63:0] exp_825_reg = 0;
      always@(posedge clk) begin
        if (exp_811) begin
          exp_825_reg <= exp_824;
        end
      end
      assign exp_825 = exp_825_reg;
      assign exp_824 = exp_820 + exp_823;
  assign exp_820 = exp_816 + exp_819;
  assign exp_816 = exp_812 + exp_815;
  assign exp_812 = exp_805;

      reg [31:0] exp_805_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_805_reg <= exp_792;
        end
      end
      assign exp_805 = exp_805_reg;
      assign exp_792 = exp_790 * exp_791;
  assign exp_790 = exp_789;
  assign exp_789 = exp_784[15:0];

      reg [31:0] exp_784_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_784_reg <= exp_774;
        end
      end
      assign exp_784 = exp_784_reg;
      assign exp_774 = exp_773 + exp_772;
  assign exp_773 = 0;

  reg [31:0] exp_772_reg;
  always@(*) begin
    case (exp_769)
      0:exp_772_reg <= exp_759;
      1:exp_772_reg <= exp_770;
      default:exp_772_reg <= exp_771;
    endcase
  end
  assign exp_772 = exp_772_reg;
  assign exp_769 = exp_763 & exp_746;
  assign exp_771 = 0;
  assign exp_770 = -exp_759;
  assign exp_791 = exp_785[15:0];

      reg [31:0] exp_785_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_785_reg <= exp_780;
        end
      end
      assign exp_785 = exp_785_reg;
      assign exp_780 = exp_779 + exp_778;
  assign exp_779 = 0;

  reg [31:0] exp_778_reg;
  always@(*) begin
    case (exp_775)
      0:exp_778_reg <= exp_760;
      1:exp_778_reg <= exp_776;
      default:exp_778_reg <= exp_777;
    endcase
  end
  assign exp_778 = exp_778_reg;
  assign exp_775 = exp_766 & exp_747;
  assign exp_777 = 0;
  assign exp_776 = -exp_760;
  assign exp_815 = exp_813 << exp_814;
  assign exp_813 = exp_806;

      reg [31:0] exp_806_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_806_reg <= exp_796;
        end
      end
      assign exp_806 = exp_806_reg;
      assign exp_796 = exp_794 * exp_795;
  assign exp_794 = exp_793;
  assign exp_793 = exp_784[15:0];
  assign exp_795 = exp_785[31:16];
  assign exp_814 = 16;
  assign exp_819 = exp_817 << exp_818;
  assign exp_817 = exp_807;

      reg [31:0] exp_807_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_807_reg <= exp_800;
        end
      end
      assign exp_807 = exp_807_reg;
      assign exp_800 = exp_798 * exp_799;
  assign exp_798 = exp_797;
  assign exp_797 = exp_784[31:16];
  assign exp_799 = exp_785[15:0];
  assign exp_818 = 16;
  assign exp_823 = exp_821 << exp_822;
  assign exp_821 = exp_808;

      reg [31:0] exp_808_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_808_reg <= exp_804;
        end
      end
      assign exp_808 = exp_808_reg;
      assign exp_804 = exp_802 * exp_803;
  assign exp_802 = exp_801;
  assign exp_801 = exp_784[31:16];
  assign exp_803 = exp_785[31:16];
  assign exp_822 = 32;
  assign exp_827 = -exp_825;
  assign exp_831 = exp_829[31:0];

  reg [31:0] exp_837_reg;
  always@(*) begin
    case (exp_630)
      0:exp_837_reg <= exp_740;
      1:exp_837_reg <= exp_741;
      default:exp_837_reg <= exp_836;
    endcase
  end
  assign exp_837 = exp_837_reg;
  assign exp_630 = exp_598[1:1];
  assign exp_836 = 0;

      reg [31:0] exp_740_reg = 0;
      always@(posedge clk) begin
        if (exp_649) begin
          exp_740_reg <= exp_734;
        end
      end
      assign exp_740 = exp_740_reg;
    
  reg [31:0] exp_734_reg;
  always@(*) begin
    case (exp_730)
      0:exp_734_reg <= exp_721;
      1:exp_734_reg <= exp_732;
      default:exp_734_reg <= exp_733;
    endcase
  end
  assign exp_734 = exp_734_reg;
  assign exp_730 = exp_729 & exp_632;
  assign exp_729 = exp_678 == exp_728;

      reg [31:0] exp_678_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_678_reg <= exp_675;
        end
      end
      assign exp_678 = exp_678_reg;
      assign exp_675 = exp_674 + exp_673;
  assign exp_674 = 0;

  reg [31:0] exp_673_reg;
  always@(*) begin
    case (exp_670)
      0:exp_673_reg <= exp_655;
      1:exp_673_reg <= exp_671;
      default:exp_673_reg <= exp_672;
    endcase
  end
  assign exp_673 = exp_673_reg;
  assign exp_670 = exp_661 & exp_632;
  assign exp_661 = exp_660 + exp_659;
  assign exp_660 = 0;
  assign exp_659 = exp_655[31:31];

      reg [31:0] exp_655_reg = 0;
      always@(posedge clk) begin
        if (exp_653) begin
          exp_655_reg <= exp_377;
        end
      end
      assign exp_655 = exp_655_reg;
      assign exp_653 = exp_635 == exp_652;
  assign exp_652 = 0;
  assign exp_632 = ~exp_631;
  assign exp_631 = exp_598[0:0];
  assign exp_672 = 0;
  assign exp_671 = -exp_655;
  assign exp_663 = exp_635 == exp_662;
  assign exp_662 = 1;
  assign exp_728 = 0;
  assign exp_733 = 0;
  assign exp_721 = exp_720 + exp_719;
  assign exp_720 = 0;

  reg [31:0] exp_719_reg;
  always@(*) begin
    case (exp_716)
      0:exp_719_reg <= exp_714;
      1:exp_719_reg <= exp_717;
      default:exp_719_reg <= exp_718;
    endcase
  end
  assign exp_719 = exp_719_reg;
  assign exp_716 = exp_680 & exp_632;

      reg [0:0] exp_680_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_680_reg <= exp_676;
        end
      end
      assign exp_680 = exp_680_reg;
      assign exp_676 = exp_658 ^ exp_661;
  assign exp_658 = exp_657 + exp_656;
  assign exp_657 = 0;
  assign exp_656 = exp_654[31:31];

      reg [31:0] exp_654_reg = 0;
      always@(posedge clk) begin
        if (exp_653) begin
          exp_654_reg <= exp_376;
        end
      end
      assign exp_654 = exp_654_reg;
      assign exp_718 = 0;

      reg [31:0] exp_714_reg = 0;
      always@(posedge clk) begin
        if (exp_647) begin
          exp_714_reg <= exp_684;
        end
      end
      assign exp_714 = exp_714_reg;
    
      reg [31:0] exp_684_reg = 0;
      always@(posedge clk) begin
        if (exp_683) begin
          exp_684_reg <= exp_711;
        end
      end
      assign exp_684 = exp_684_reg;
    
  reg [31:0] exp_711_reg;
  always@(*) begin
    case (exp_645)
      0:exp_711_reg <= exp_703;
      1:exp_711_reg <= exp_709;
      default:exp_711_reg <= exp_710;
    endcase
  end
  assign exp_711 = exp_711_reg;
  assign exp_645 = exp_635 == exp_644;
  assign exp_644 = 2;
  assign exp_710 = 0;

  reg [31:0] exp_703_reg;
  always@(*) begin
    case (exp_693)
      0:exp_703_reg <= exp_697;
      1:exp_703_reg <= exp_701;
      default:exp_703_reg <= exp_702;
    endcase
  end
  assign exp_703 = exp_703_reg;
  assign exp_693 = ~exp_692;
  assign exp_692 = exp_691[32:32];
  assign exp_691 = exp_690 - exp_678;
  assign exp_690 = exp_689;
  assign exp_689 = {exp_687, exp_688};  assign exp_687 = exp_682[31:0];

      reg [31:0] exp_682_reg = 0;
      always@(posedge clk) begin
        if (exp_681) begin
          exp_682_reg <= exp_708;
        end
      end
      assign exp_682 = exp_682_reg;
    
  reg [32:0] exp_708_reg;
  always@(*) begin
    case (exp_645)
      0:exp_708_reg <= exp_695;
      1:exp_708_reg <= exp_706;
      default:exp_708_reg <= exp_707;
    endcase
  end
  assign exp_708 = exp_708_reg;
  assign exp_707 = 0;

  reg [32:0] exp_695_reg;
  always@(*) begin
    case (exp_693)
      0:exp_695_reg <= exp_689;
      1:exp_695_reg <= exp_691;
      default:exp_695_reg <= exp_694;
    endcase
  end
  assign exp_695 = exp_695_reg;
  assign exp_694 = 0;
  assign exp_706 = 0;
  assign exp_681 = 1;
  assign exp_688 = exp_686[31:31];

      reg [31:0] exp_686_reg = 0;
      always@(posedge clk) begin
        if (exp_685) begin
          exp_686_reg <= exp_713;
        end
      end
      assign exp_686 = exp_686_reg;
    
  reg [31:0] exp_713_reg;
  always@(*) begin
    case (exp_645)
      0:exp_713_reg <= exp_705;
      1:exp_713_reg <= exp_677;
      default:exp_713_reg <= exp_712;
    endcase
  end
  assign exp_713 = exp_713_reg;
  assign exp_712 = 0;
  assign exp_705 = exp_686 << exp_704;
  assign exp_704 = 1;

      reg [31:0] exp_677_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_677_reg <= exp_669;
        end
      end
      assign exp_677 = exp_677_reg;
      assign exp_669 = exp_668 + exp_667;
  assign exp_668 = 0;

  reg [31:0] exp_667_reg;
  always@(*) begin
    case (exp_664)
      0:exp_667_reg <= exp_654;
      1:exp_667_reg <= exp_665;
      default:exp_667_reg <= exp_666;
    endcase
  end
  assign exp_667 = exp_667_reg;
  assign exp_664 = exp_658 & exp_632;
  assign exp_666 = 0;
  assign exp_665 = -exp_654;
  assign exp_685 = 1;
  assign exp_702 = 0;
  assign exp_697 = exp_684 << exp_696;
  assign exp_696 = 1;
  assign exp_701 = exp_699 | exp_700;
  assign exp_699 = exp_684 << exp_698;
  assign exp_698 = 1;
  assign exp_700 = 1;
  assign exp_709 = 0;
  assign exp_683 = 1;
  assign exp_647 = exp_635 == exp_646;
  assign exp_646 = 35;
  assign exp_717 = -exp_714;
  assign exp_732 = $signed(exp_731);
  assign exp_731 = -1;
  assign exp_649 = exp_635 == exp_648;
  assign exp_648 = 36;

      reg [31:0] exp_741_reg = 0;
      always@(posedge clk) begin
        if (exp_649) begin
          exp_741_reg <= exp_739;
        end
      end
      assign exp_741 = exp_741_reg;
    
  reg [31:0] exp_739_reg;
  always@(*) begin
    case (exp_737)
      0:exp_739_reg <= exp_727;
      1:exp_739_reg <= exp_654;
      default:exp_739_reg <= exp_738;
    endcase
  end
  assign exp_739 = exp_739_reg;
  assign exp_737 = exp_736 & exp_632;
  assign exp_736 = exp_678 == exp_735;
  assign exp_735 = 0;
  assign exp_738 = 0;
  assign exp_727 = exp_726 + exp_725;
  assign exp_726 = 0;

  reg [31:0] exp_725_reg;
  always@(*) begin
    case (exp_722)
      0:exp_725_reg <= exp_715;
      1:exp_725_reg <= exp_723;
      default:exp_725_reg <= exp_724;
    endcase
  end
  assign exp_725 = exp_725_reg;
  assign exp_722 = exp_679 & exp_632;

      reg [0:0] exp_679_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_679_reg <= exp_658;
        end
      end
      assign exp_679 = exp_679_reg;
      assign exp_724 = 0;

      reg [31:0] exp_715_reg = 0;
      always@(posedge clk) begin
        if (exp_647) begin
          exp_715_reg <= exp_682;
        end
      end
      assign exp_715 = exp_715_reg;
      assign exp_723 = -exp_715;
  assign exp_310 = $signed(exp_309);
  assign exp_309 = 0;
  assign exp_539 = exp_374 != exp_375;
  assign exp_552 = 0;
  assign exp_553 = 0;
  assign exp_540 = $signed(exp_374) < $signed(exp_375);
  assign exp_541 = $signed(exp_374) >= $signed(exp_375);
  assign exp_546 = exp_543 < exp_545;
  assign exp_543 = exp_542 + exp_374;
  assign exp_542 = 0;
  assign exp_545 = exp_544 + exp_375;
  assign exp_544 = 0;
  assign exp_551 = exp_548 >= exp_550;
  assign exp_548 = exp_547 + exp_374;
  assign exp_547 = 0;
  assign exp_550 = exp_549 + exp_375;
  assign exp_549 = 0;
  assign exp_866 = 0;
  assign exp_865 = exp_264 + exp_864;
  assign exp_864 = 4;

  reg [32:0] exp_596_reg;
  always@(*) begin
    case (exp_397)
      0:exp_596_reg <= exp_586;
      1:exp_596_reg <= exp_594;
      default:exp_596_reg <= exp_595;
    endcase
  end
  assign exp_596 = exp_596_reg;
  assign exp_595 = 0;
  assign exp_586 = exp_585 + exp_383;

  reg [31:0] exp_585_reg;
  always@(*) begin
    case (exp_395)
      0:exp_585_reg <= exp_571;
      1:exp_585_reg <= exp_583;
      default:exp_585_reg <= exp_584;
    endcase
  end
  assign exp_585 = exp_585_reg;
  assign exp_584 = 0;
  assign exp_571 = $signed(exp_570);
  assign exp_570 = exp_569 + exp_568;
  assign exp_569 = 0;
  assign exp_568 = {exp_567, exp_564};  assign exp_567 = {exp_566, exp_563};  assign exp_566 = {exp_565, exp_562};  assign exp_565 = {exp_560, exp_561};  assign exp_560 = exp_382[31:31];
  assign exp_561 = exp_382[7:7];
  assign exp_562 = exp_382[30:25];
  assign exp_563 = exp_382[11:8];
  assign exp_564 = 0;
  assign exp_583 = $signed(exp_582);
  assign exp_582 = exp_581 + exp_580;
  assign exp_581 = 0;
  assign exp_580 = {exp_579, exp_576};  assign exp_579 = {exp_578, exp_575};  assign exp_578 = {exp_577, exp_574};  assign exp_577 = {exp_572, exp_573};  assign exp_572 = exp_382[31:31];
  assign exp_573 = exp_382[19:12];
  assign exp_574 = exp_382[20:20];
  assign exp_575 = exp_382[30:21];
  assign exp_576 = 0;

      reg [31:0] exp_383_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_383_reg <= exp_266;
        end
      end
      assign exp_383 = exp_383_reg;
      assign exp_594 = exp_593 & exp_592;
  assign exp_593 = $signed(exp_591);
  assign exp_591 = exp_374 + exp_590;
  assign exp_590 = $signed(exp_589);
  assign exp_589 = exp_588 + exp_587;
  assign exp_588 = 0;
  assign exp_587 = exp_382[31:20];
  assign exp_592 = 4294967294;
  assign exp_263 = exp_256 & exp_254;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_265;
  assign exp_398 = 3;
  assign exp_244 = ~exp_229;
  assign exp_229 = exp_6;
  assign exp_200 = exp_184 & exp_185;
  assign exp_184 = exp_192;
  assign exp_192 = exp_5 & exp_191;
  assign exp_185 = exp_6;
  assign exp_181 = exp_2;

      reg [31:0] exp_221_reg = 0;
      always@(posedge clk) begin
        if (exp_220) begin
          exp_221_reg <= exp_203;
        end
      end
      assign exp_221 = exp_221_reg;
      assign exp_203 = exp_2;
  assign exp_220 = exp_206 & exp_207;
  assign exp_206 = exp_214;
  assign exp_214 = exp_5 & exp_213;
  assign exp_207 = exp_6;
  assign stdin_ready_out = exp_245;
  assign stdout_valid_out = exp_200;
  assign stdout_out = exp_181;
  assign leds_out = exp_221;

endmodule