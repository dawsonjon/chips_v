
module test(clk, debug_ready_in, stdout_ready_in, spare_ready_in, debug_valid_out, debug_out, stdout_valid_out, stdout_out, spare_valid_out, spare_out);
  input [0:0] debug_ready_in;
  input [0:0] stdout_ready_in;
  input [0:0] spare_ready_in;
  input [0:0] clk;
  output [0:0] debug_valid_out;
  output [31:0] debug_out;
  output [0:0] stdout_valid_out;
  output [31:0] stdout_out;
  output [0:0] spare_valid_out;
  output [31:0] spare_out;
  wire [0:0] exp_159;
  wire [0:0] exp_143;
  wire [0:0] exp_151;
  wire [0:0] exp_5;
  wire [0:0] exp_243;
  wire [0:0] exp_527;
  wire [0:0] exp_392;
  wire [6:0] exp_377;
  wire [31:0] exp_375;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [11:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_257;
  wire [32:0] exp_859;
  wire [0:0] exp_855;
  wire [0:0] exp_552;
  wire [0:0] exp_530;
  wire [0:0] exp_388;
  wire [6:0] exp_387;
  wire [0:0] exp_390;
  wire [6:0] exp_389;
  wire [0:0] exp_551;
  wire [0:0] exp_396;
  wire [6:0] exp_395;
  wire [0:0] exp_550;
  wire [0:0] exp_549;
  wire [0:0] exp_548;
  wire [2:0] exp_378;
  wire [0:0] exp_547;
  wire [0:0] exp_531;
  wire [31:0] exp_367;
  wire [31:0] exp_305;
  wire [0:0] exp_301;
  wire [4:0] exp_281;
  wire [0:0] exp_300;
  wire [0:0] exp_304;
  wire [31:0] exp_297;
  wire [0:0] exp_278;
  wire [0:0] exp_850;
  wire [0:0] exp_849;
  wire [0:0] exp_848;
  wire [0:0] exp_847;
  wire [4:0] exp_260;
  wire [4:0] exp_842;
  wire [0:0] exp_841;
  wire [0:0] exp_434;
  wire [0:0] exp_433;
  wire [0:0] exp_432;
  wire [0:0] exp_431;
  wire [0:0] exp_430;
  wire [0:0] exp_429;
  wire [0:0] exp_380;
  wire [4:0] exp_379;
  wire [0:0] exp_382;
  wire [5:0] exp_381;
  wire [0:0] exp_384;
  wire [5:0] exp_383;
  wire [0:0] exp_386;
  wire [4:0] exp_385;
  wire [0:0] exp_836;
  wire [0:0] exp_835;
  wire [0:0] exp_621;
  wire [0:0] exp_595;
  wire [0:0] exp_593;
  wire [6:0] exp_591;
  wire [5:0] exp_592;
  wire [0:0] exp_594;
  wire [0:0] exp_620;
  wire [2:0] exp_590;
  wire [0:0] exp_834;
  wire [0:0] exp_832;
  wire [0:0] exp_825;
  wire [2:0] exp_740;
  wire [2:0] exp_747;
  wire [0:0] exp_742;
  wire [2:0] exp_741;
  wire [0:0] exp_746;
  wire [2:0] exp_744;
  wire [0:0] exp_743;
  wire [0:0] exp_745;
  wire [0:0] exp_736;
  wire [0:0] exp_735;
  wire [0:0] exp_734;
  wire [2:0] exp_824;
  wire [0:0] exp_833;
  wire [0:0] exp_643;
  wire [5:0] exp_627;
  wire [5:0] exp_634;
  wire [0:0] exp_629;
  wire [5:0] exp_628;
  wire [0:0] exp_633;
  wire [5:0] exp_631;
  wire [0:0] exp_630;
  wire [0:0] exp_632;
  wire [5:0] exp_642;
  wire [0:0] exp_255;
  wire [0:0] exp_254;
  wire [0:0] exp_252;
  wire [0:0] exp_251;
  wire [0:0] exp_249;
  wire [0:0] exp_250;
  wire [0:0] exp_248;
  wire [0:0] exp_860;
  wire [0:0] exp_247;
  wire [0:0] exp_246;
  wire [0:0] exp_864;
  wire [0:0] exp_863;
  wire [0:0] exp_862;
  wire [0:0] exp_861;
  wire [0:0] exp_242;
  wire [0:0] exp_233;
  wire [0:0] exp_228;
  wire [0:0] exp_225;
  wire [31:0] exp_1;
  wire [31:0] exp_239;
  wire [31:0] exp_446;
  wire [31:0] exp_445;
  wire [31:0] exp_444;
  wire [31:0] exp_443;
  wire [11:0] exp_442;
  wire [11:0] exp_441;
  wire [11:0] exp_440;
  wire [0:0] exp_394;
  wire [5:0] exp_393;
  wire [0:0] exp_439;
  wire [11:0] exp_435;
  wire [11:0] exp_438;
  wire [6:0] exp_436;
  wire [4:0] exp_437;
  wire [35:0] exp_224;
  wire [0:0] exp_227;
  wire [35:0] exp_226;
  wire [0:0] exp_232;
  wire [0:0] exp_211;
  wire [0:0] exp_206;
  wire [0:0] exp_203;
  wire [35:0] exp_202;
  wire [0:0] exp_205;
  wire [35:0] exp_204;
  wire [0:0] exp_210;
  wire [0:0] exp_177;
  wire [0:0] exp_172;
  wire [0:0] exp_169;
  wire [31:0] exp_168;
  wire [0:0] exp_171;
  wire [31:0] exp_170;
  wire [0:0] exp_176;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [28:0] exp_146;
  wire [0:0] exp_149;
  wire [28:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [13:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_244;
  wire [0:0] exp_529;
  wire [0:0] exp_528;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_157;
  wire [0:0] exp_164;
  wire [0:0] exp_189;
  wire [0:0] exp_198;
  wire [0:0] exp_213;
  wire [0:0] exp_220;
  wire [0:0] exp_235;
  wire [0:0] exp_838;
  wire [0:0] exp_837;
  wire [0:0] exp_253;
  wire [0:0] exp_296;
  wire [31:0] exp_268;
  wire [0:0] exp_267;
  wire [1:0] exp_276;
  wire [4:0] exp_263;
  wire [0:0] exp_266;
  wire [0:0] exp_844;
  wire [0:0] exp_843;
  wire [4:0] exp_262;
  wire [31:0] exp_264;
  wire [31:0] exp_840;
  wire [0:0] exp_839;
  wire [31:0] exp_477;
  wire [0:0] exp_476;
  wire [31:0] exp_428;
  wire [2:0] exp_371;
  wire [2:0] exp_362;
  wire [0:0] exp_359;
  wire [0:0] exp_293;
  wire [6:0] exp_283;
  wire [6:0] exp_292;
  wire [0:0] exp_295;
  wire [6:0] exp_294;
  wire [0:0] exp_361;
  wire [2:0] exp_349;
  wire [0:0] exp_291;
  wire [4:0] exp_290;
  wire [0:0] exp_348;
  wire [2:0] exp_336;
  wire [0:0] exp_289;
  wire [5:0] exp_288;
  wire [0:0] exp_335;
  wire [2:0] exp_285;
  wire [0:0] exp_334;
  wire [0:0] exp_347;
  wire [0:0] exp_360;
  wire [0:0] exp_366;
  wire [0:0] exp_427;
  wire [31:0] exp_407;
  wire [0:0] exp_373;
  wire [0:0] exp_365;
  wire [0:0] exp_351;
  wire [0:0] exp_338;
  wire [0:0] exp_324;
  wire [0:0] exp_322;
  wire [0:0] exp_323;
  wire [0:0] exp_287;
  wire [4:0] exp_286;
  wire [0:0] exp_337;
  wire [0:0] exp_350;
  wire [0:0] exp_364;
  wire [0:0] exp_363;
  wire [0:0] exp_406;
  wire [31:0] exp_404;
  wire [31:0] exp_369;
  wire [31:0] exp_355;
  wire [0:0] exp_352;
  wire [0:0] exp_354;
  wire [31:0] exp_344;
  wire [0:0] exp_343;
  wire [31:0] exp_330;
  wire [0:0] exp_329;
  wire [31:0] exp_328;
  wire [31:0] exp_326;
  wire [19:0] exp_325;
  wire [3:0] exp_327;
  wire [31:0] exp_342;
  wire [31:0] exp_340;
  wire [19:0] exp_339;
  wire [3:0] exp_341;
  wire [31:0] exp_353;
  wire [31:0] exp_370;
  wire [31:0] exp_358;
  wire [0:0] exp_356;
  wire [0:0] exp_357;
  wire [31:0] exp_346;
  wire [0:0] exp_345;
  wire [31:0] exp_333;
  wire [0:0] exp_332;
  wire [31:0] exp_317;
  wire [0:0] exp_316;
  wire [31:0] exp_311;
  wire [0:0] exp_307;
  wire [4:0] exp_282;
  wire [0:0] exp_306;
  wire [0:0] exp_310;
  wire [31:0] exp_299;
  wire [0:0] exp_279;
  wire [0:0] exp_854;
  wire [0:0] exp_853;
  wire [0:0] exp_852;
  wire [0:0] exp_851;
  wire [4:0] exp_261;
  wire [0:0] exp_298;
  wire [31:0] exp_275;
  wire [0:0] exp_274;
  wire [1:0] exp_277;
  wire [4:0] exp_270;
  wire [0:0] exp_273;
  wire [0:0] exp_846;
  wire [0:0] exp_845;
  wire [4:0] exp_269;
  wire [31:0] exp_271;
  wire [31:0] exp_280;
  wire [31:0] exp_309;
  wire [0:0] exp_308;
  wire [31:0] exp_315;
  wire [31:0] exp_312;
  wire [31:0] exp_314;
  wire [11:0] exp_313;
  wire [31:0] exp_331;
  wire [31:0] exp_259;
  wire [0:0] exp_258;
  wire [31:0] exp_405;
  wire [31:0] exp_409;
  wire [31:0] exp_408;
  wire [5:0] exp_403;
  wire [5:0] exp_402;
  wire [5:0] exp_401;
  wire [4:0] exp_372;
  wire [4:0] exp_321;
  wire [0:0] exp_320;
  wire [4:0] exp_319;
  wire [4:0] exp_284;
  wire [31:0] exp_425;
  wire [1:0] exp_411;
  wire [0:0] exp_410;
  wire [31:0] exp_426;
  wire [1:0] exp_417;
  wire [0:0] exp_416;
  wire [31:0] exp_413;
  wire [31:0] exp_412;
  wire [31:0] exp_415;
  wire [31:0] exp_414;
  wire [31:0] exp_418;
  wire [31:0] exp_422;
  wire [32:0] exp_421;
  wire [32:0] exp_419;
  wire [0:0] exp_400;
  wire [0:0] exp_374;
  wire [0:0] exp_318;
  wire [0:0] exp_399;
  wire [0:0] exp_398;
  wire [0:0] exp_397;
  wire [32:0] exp_420;
  wire [31:0] exp_423;
  wire [31:0] exp_424;
  wire [31:0] exp_475;
  wire [0:0] exp_474;
  wire [31:0] exp_465;
  wire [7:0] exp_464;
  wire [7:0] exp_463;
  wire [7:0] exp_458;
  wire [1:0] exp_449;
  wire [1:0] exp_448;
  wire [1:0] exp_447;
  wire [0:0] exp_457;
  wire [7:0] exp_453;
  wire [31:0] exp_241;
  wire [31:0] exp_231;
  wire [0:0] exp_230;
  wire [31:0] exp_209;
  wire [0:0] exp_208;
  wire [31:0] exp_175;
  wire [0:0] exp_174;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [11:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_245;
  wire [3:0] exp_526;
  wire [0:0] exp_525;
  wire [3:0] exp_513;
  wire [3:0] exp_509;
  wire [1:0] exp_512;
  wire [1:0] exp_511;
  wire [1:0] exp_510;
  wire [3:0] exp_518;
  wire [3:0] exp_514;
  wire [0:0] exp_517;
  wire [0:0] exp_516;
  wire [0:0] exp_515;
  wire [3:0] exp_519;
  wire [3:0] exp_520;
  wire [3:0] exp_521;
  wire [3:0] exp_522;
  wire [3:0] exp_523;
  wire [3:0] exp_524;
  wire [11:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_240;
  wire [31:0] exp_508;
  wire [0:0] exp_507;
  wire [31:0] exp_495;
  wire [0:0] exp_494;
  wire [31:0] exp_481;
  wire [7:0] exp_480;
  wire [7:0] exp_479;
  wire [7:0] exp_478;
  wire [31:0] exp_368;
  wire [31:0] exp_489;
  wire [3:0] exp_488;
  wire [31:0] exp_491;
  wire [4:0] exp_490;
  wire [31:0] exp_493;
  wire [4:0] exp_492;
  wire [31:0] exp_499;
  wire [0:0] exp_452;
  wire [0:0] exp_451;
  wire [0:0] exp_450;
  wire [0:0] exp_498;
  wire [31:0] exp_485;
  wire [15:0] exp_484;
  wire [15:0] exp_483;
  wire [15:0] exp_482;
  wire [31:0] exp_497;
  wire [4:0] exp_496;
  wire [31:0] exp_501;
  wire [31:0] exp_500;
  wire [31:0] exp_487;
  wire [31:0] exp_486;
  wire [31:0] exp_502;
  wire [31:0] exp_503;
  wire [31:0] exp_504;
  wire [31:0] exp_505;
  wire [31:0] exp_506;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [11:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [11:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [11:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [11:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [11:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [11:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [11:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [11:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [11:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [11:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [11:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [11:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_160;
  wire [31:0] exp_163;
  wire [31:0] exp_194;
  wire [0:0] exp_190;
  wire [31:0] exp_161;
  wire [0:0] exp_193;
  wire [31:0] exp_191;
  wire [63:0] exp_179;
  wire [63:0] exp_186;
  wire [0:0] exp_181;
  wire [63:0] exp_180;
  wire [0:0] exp_185;
  wire [63:0] exp_183;
  wire [0:0] exp_182;
  wire [0:0] exp_184;
  wire [0:0] exp_178;
  wire [31:0] exp_192;
  wire [31:0] exp_197;
  wire [31:0] exp_216;
  wire [31:0] exp_219;
  wire [31:0] exp_238;
  wire [7:0] exp_454;
  wire [7:0] exp_455;
  wire [7:0] exp_456;
  wire [31:0] exp_468;
  wire [15:0] exp_467;
  wire [15:0] exp_466;
  wire [15:0] exp_462;
  wire [0:0] exp_461;
  wire [15:0] exp_459;
  wire [15:0] exp_460;
  wire [31:0] exp_469;
  wire [31:0] exp_470;
  wire [31:0] exp_471;
  wire [31:0] exp_472;
  wire [31:0] exp_473;
  wire [31:0] exp_831;
  wire [0:0] exp_830;
  wire [31:0] exp_827;
  wire [0:0] exp_598;
  wire [0:0] exp_597;
  wire [0:0] exp_596;
  wire [0:0] exp_826;
  wire [31:0] exp_822;
  wire [63:0] exp_821;
  wire [0:0] exp_818;
  wire [0:0] exp_801;
  wire [0:0] exp_778;
  wire [0:0] exp_775;
  wire [0:0] exp_773;
  wire [0:0] exp_755;
  wire [0:0] exp_754;
  wire [0:0] exp_753;
  wire [31:0] exp_751;
  wire [0:0] exp_750;
  wire [0:0] exp_749;
  wire [0:0] exp_738;
  wire [0:0] exp_737;
  wire [0:0] exp_601;
  wire [0:0] exp_600;
  wire [0:0] exp_599;
  wire [0:0] exp_604;
  wire [0:0] exp_603;
  wire [1:0] exp_602;
  wire [0:0] exp_774;
  wire [0:0] exp_758;
  wire [0:0] exp_757;
  wire [0:0] exp_756;
  wire [31:0] exp_752;
  wire [0:0] exp_739;
  wire [0:0] exp_760;
  wire [0:0] exp_759;
  wire [0:0] exp_780;
  wire [1:0] exp_779;
  wire [0:0] exp_803;
  wire [1:0] exp_802;
  wire [0:0] exp_820;
  wire [63:0] exp_817;
  wire [63:0] exp_816;
  wire [63:0] exp_812;
  wire [63:0] exp_808;
  wire [63:0] exp_804;
  wire [31:0] exp_797;
  wire [31:0] exp_784;
  wire [31:0] exp_782;
  wire [15:0] exp_781;
  wire [31:0] exp_776;
  wire [31:0] exp_766;
  wire [31:0] exp_765;
  wire [31:0] exp_764;
  wire [0:0] exp_761;
  wire [0:0] exp_763;
  wire [31:0] exp_762;
  wire [15:0] exp_783;
  wire [31:0] exp_777;
  wire [31:0] exp_772;
  wire [31:0] exp_771;
  wire [31:0] exp_770;
  wire [0:0] exp_767;
  wire [0:0] exp_769;
  wire [31:0] exp_768;
  wire [63:0] exp_807;
  wire [63:0] exp_805;
  wire [31:0] exp_798;
  wire [31:0] exp_788;
  wire [31:0] exp_786;
  wire [15:0] exp_785;
  wire [15:0] exp_787;
  wire [4:0] exp_806;
  wire [63:0] exp_811;
  wire [63:0] exp_809;
  wire [31:0] exp_799;
  wire [31:0] exp_792;
  wire [31:0] exp_790;
  wire [15:0] exp_789;
  wire [15:0] exp_791;
  wire [4:0] exp_810;
  wire [63:0] exp_815;
  wire [63:0] exp_813;
  wire [31:0] exp_800;
  wire [31:0] exp_796;
  wire [31:0] exp_794;
  wire [15:0] exp_793;
  wire [15:0] exp_795;
  wire [5:0] exp_814;
  wire [63:0] exp_819;
  wire [31:0] exp_823;
  wire [31:0] exp_829;
  wire [0:0] exp_622;
  wire [0:0] exp_828;
  wire [31:0] exp_732;
  wire [31:0] exp_726;
  wire [0:0] exp_722;
  wire [0:0] exp_721;
  wire [31:0] exp_670;
  wire [31:0] exp_667;
  wire [31:0] exp_666;
  wire [31:0] exp_665;
  wire [0:0] exp_662;
  wire [0:0] exp_653;
  wire [0:0] exp_652;
  wire [0:0] exp_651;
  wire [31:0] exp_647;
  wire [0:0] exp_645;
  wire [0:0] exp_644;
  wire [0:0] exp_624;
  wire [0:0] exp_623;
  wire [0:0] exp_664;
  wire [31:0] exp_663;
  wire [0:0] exp_655;
  wire [0:0] exp_654;
  wire [0:0] exp_720;
  wire [0:0] exp_725;
  wire [31:0] exp_713;
  wire [31:0] exp_712;
  wire [31:0] exp_711;
  wire [0:0] exp_708;
  wire [0:0] exp_672;
  wire [0:0] exp_668;
  wire [0:0] exp_650;
  wire [0:0] exp_649;
  wire [0:0] exp_648;
  wire [31:0] exp_646;
  wire [0:0] exp_710;
  wire [31:0] exp_706;
  wire [31:0] exp_676;
  wire [31:0] exp_703;
  wire [0:0] exp_637;
  wire [1:0] exp_636;
  wire [0:0] exp_702;
  wire [31:0] exp_695;
  wire [0:0] exp_685;
  wire [0:0] exp_684;
  wire [32:0] exp_683;
  wire [32:0] exp_682;
  wire [32:0] exp_681;
  wire [31:0] exp_679;
  wire [31:0] exp_674;
  wire [32:0] exp_700;
  wire [0:0] exp_699;
  wire [32:0] exp_687;
  wire [0:0] exp_686;
  wire [0:0] exp_698;
  wire [0:0] exp_673;
  wire [0:0] exp_680;
  wire [31:0] exp_678;
  wire [31:0] exp_705;
  wire [0:0] exp_704;
  wire [31:0] exp_697;
  wire [0:0] exp_696;
  wire [31:0] exp_669;
  wire [31:0] exp_661;
  wire [31:0] exp_660;
  wire [31:0] exp_659;
  wire [0:0] exp_656;
  wire [0:0] exp_658;
  wire [31:0] exp_657;
  wire [0:0] exp_677;
  wire [0:0] exp_694;
  wire [31:0] exp_689;
  wire [0:0] exp_688;
  wire [31:0] exp_693;
  wire [31:0] exp_691;
  wire [0:0] exp_690;
  wire [0:0] exp_692;
  wire [0:0] exp_701;
  wire [0:0] exp_675;
  wire [0:0] exp_639;
  wire [5:0] exp_638;
  wire [31:0] exp_709;
  wire [31:0] exp_724;
  wire [0:0] exp_723;
  wire [0:0] exp_641;
  wire [5:0] exp_640;
  wire [31:0] exp_733;
  wire [31:0] exp_731;
  wire [0:0] exp_729;
  wire [0:0] exp_728;
  wire [0:0] exp_727;
  wire [0:0] exp_730;
  wire [31:0] exp_719;
  wire [31:0] exp_718;
  wire [31:0] exp_717;
  wire [0:0] exp_714;
  wire [0:0] exp_671;
  wire [0:0] exp_716;
  wire [31:0] exp_707;
  wire [31:0] exp_715;
  wire [31:0] exp_303;
  wire [0:0] exp_302;
  wire [0:0] exp_532;
  wire [0:0] exp_545;
  wire [0:0] exp_546;
  wire [0:0] exp_533;
  wire [0:0] exp_534;
  wire [0:0] exp_539;
  wire [31:0] exp_536;
  wire [31:0] exp_535;
  wire [31:0] exp_538;
  wire [31:0] exp_537;
  wire [0:0] exp_544;
  wire [31:0] exp_541;
  wire [31:0] exp_540;
  wire [31:0] exp_543;
  wire [31:0] exp_542;
  wire [0:0] exp_858;
  wire [31:0] exp_857;
  wire [2:0] exp_856;
  wire [32:0] exp_589;
  wire [0:0] exp_588;
  wire [31:0] exp_579;
  wire [31:0] exp_578;
  wire [0:0] exp_577;
  wire [31:0] exp_564;
  wire [12:0] exp_563;
  wire [12:0] exp_562;
  wire [12:0] exp_561;
  wire [11:0] exp_560;
  wire [7:0] exp_559;
  wire [1:0] exp_558;
  wire [0:0] exp_553;
  wire [0:0] exp_554;
  wire [5:0] exp_555;
  wire [3:0] exp_556;
  wire [0:0] exp_557;
  wire [31:0] exp_576;
  wire [20:0] exp_575;
  wire [20:0] exp_574;
  wire [20:0] exp_573;
  wire [19:0] exp_572;
  wire [9:0] exp_571;
  wire [8:0] exp_570;
  wire [0:0] exp_565;
  wire [7:0] exp_566;
  wire [0:0] exp_567;
  wire [9:0] exp_568;
  wire [0:0] exp_569;
  wire [31:0] exp_376;
  wire [32:0] exp_587;
  wire [32:0] exp_586;
  wire [31:0] exp_584;
  wire [31:0] exp_583;
  wire [11:0] exp_582;
  wire [11:0] exp_581;
  wire [11:0] exp_580;
  wire [32:0] exp_585;
  wire [0:0] exp_256;
  wire [0:0] exp_80;
  wire [11:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_391;
  wire [0:0] exp_144;
  wire [31:0] exp_140;
  wire [0:0] exp_215;
  wire [0:0] exp_199;
  wire [0:0] exp_207;
  wire [0:0] exp_200;
  wire [31:0] exp_196;
  wire [0:0] exp_237;
  wire [0:0] exp_221;
  wire [0:0] exp_229;
  wire [0:0] exp_222;
  wire [31:0] exp_218;

  assign exp_159 = exp_143 & exp_144;
  assign exp_143 = exp_151;
  assign exp_151 = exp_5 & exp_150;
  assign exp_5 = exp_243;
  assign exp_243 = exp_527;
  assign exp_527 = exp_392 | exp_394;
  assign exp_392 = exp_377 == exp_391;
  assign exp_377 = exp_375[6:0];

      reg [31:0] exp_375_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_375_reg <= exp_96;
        end
      end
      assign exp_375 = exp_375_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};

  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_257;

      reg [31:0] exp_257_reg = 0;
      always@(posedge clk) begin
        if (exp_256) begin
          exp_257_reg <= exp_859;
        end
      end
      assign exp_257 = exp_257_reg;
    
  reg [32:0] exp_859_reg;
  always@(*) begin
    case (exp_855)
      0:exp_859_reg <= exp_857;
      1:exp_859_reg <= exp_589;
      default:exp_859_reg <= exp_858;
    endcase
  end
  assign exp_859 = exp_859_reg;
  assign exp_855 = exp_552 & exp_255;
  assign exp_552 = exp_530 | exp_551;
  assign exp_530 = exp_388 | exp_390;
  assign exp_388 = exp_377 == exp_387;
  assign exp_387 = 111;
  assign exp_390 = exp_377 == exp_389;
  assign exp_389 = 103;

  reg [0:0] exp_551_reg;
  always@(*) begin
    case (exp_396)
      0:exp_551_reg <= exp_549;
      1:exp_551_reg <= exp_548;
      default:exp_551_reg <= exp_550;
    endcase
  end
  assign exp_551 = exp_551_reg;
  assign exp_396 = exp_377 == exp_395;
  assign exp_395 = 99;
  assign exp_550 = 0;
  assign exp_549 = 0;

  reg [0:0] exp_548_reg;
  always@(*) begin
    case (exp_378)
      0:exp_548_reg <= exp_531;
      1:exp_548_reg <= exp_532;
      2:exp_548_reg <= exp_545;
      3:exp_548_reg <= exp_546;
      4:exp_548_reg <= exp_533;
      5:exp_548_reg <= exp_534;
      6:exp_548_reg <= exp_539;
      7:exp_548_reg <= exp_544;
      default:exp_548_reg <= exp_547;
    endcase
  end
  assign exp_548 = exp_548_reg;
  assign exp_378 = exp_375[14:12];
  assign exp_547 = 0;
  assign exp_531 = exp_367 == exp_368;

      reg [31:0] exp_367_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_367_reg <= exp_305;
        end
      end
      assign exp_367 = exp_367_reg;
    
  reg [31:0] exp_305_reg;
  always@(*) begin
    case (exp_301)
      0:exp_305_reg <= exp_297;
      1:exp_305_reg <= exp_303;
      default:exp_305_reg <= exp_304;
    endcase
  end
  assign exp_305 = exp_305_reg;
  assign exp_301 = exp_281 == exp_300;
  assign exp_281 = exp_96[19:15];
  assign exp_300 = 0;
  assign exp_304 = 0;

  reg [31:0] exp_297_reg;
  always@(*) begin
    case (exp_278)
      0:exp_297_reg <= exp_268;
      1:exp_297_reg <= exp_280;
      default:exp_297_reg <= exp_296;
    endcase
  end
  assign exp_297 = exp_297_reg;
  assign exp_278 = exp_850;
  assign exp_850 = exp_849 & exp_247;
  assign exp_849 = exp_848 & exp_255;
  assign exp_848 = exp_847 & exp_841;
  assign exp_847 = exp_260 == exp_842;
  assign exp_260 = exp_96[19:15];
  assign exp_842 = exp_375[11:7];
  assign exp_841 = exp_434 | exp_836;
  assign exp_434 = exp_433 | exp_392;
  assign exp_433 = exp_432 | exp_386;
  assign exp_432 = exp_431 | exp_384;
  assign exp_431 = exp_430 | exp_390;
  assign exp_430 = exp_429 | exp_388;
  assign exp_429 = exp_380 | exp_382;
  assign exp_380 = exp_377 == exp_379;
  assign exp_379 = 19;
  assign exp_382 = exp_377 == exp_381;
  assign exp_381 = 51;
  assign exp_384 = exp_377 == exp_383;
  assign exp_383 = 55;
  assign exp_386 = exp_377 == exp_385;
  assign exp_385 = 23;
  assign exp_836 = exp_835 & exp_595;

  reg [0:0] exp_835_reg;
  always@(*) begin
    case (exp_621)
      0:exp_835_reg <= exp_832;
      1:exp_835_reg <= exp_833;
      default:exp_835_reg <= exp_834;
    endcase
  end
  assign exp_835 = exp_835_reg;
  assign exp_621 = exp_595 & exp_620;
  assign exp_595 = exp_593 & exp_594;
  assign exp_593 = exp_591 == exp_592;
  assign exp_591 = exp_375[6:0];
  assign exp_592 = 51;
  assign exp_594 = exp_375[25:25];
  assign exp_620 = exp_590[2:2];
  assign exp_590 = exp_375[14:12];
  assign exp_834 = 0;
  assign exp_832 = exp_825 & exp_595;
  assign exp_825 = exp_740 == exp_824;

      reg [2:0] exp_740_reg = 0;
      always@(posedge clk) begin
        if (exp_736) begin
          exp_740_reg <= exp_747;
        end
      end
      assign exp_740 = exp_740_reg;
    
  reg [2:0] exp_747_reg;
  always@(*) begin
    case (exp_742)
      0:exp_747_reg <= exp_744;
      1:exp_747_reg <= exp_745;
      default:exp_747_reg <= exp_746;
    endcase
  end
  assign exp_747 = exp_747_reg;
  assign exp_742 = exp_740 == exp_741;
  assign exp_741 = 4;
  assign exp_746 = 0;
  assign exp_744 = exp_740 + exp_743;
  assign exp_743 = 1;
  assign exp_745 = 0;
  assign exp_736 = exp_595 & exp_735;
  assign exp_735 = ~exp_734;
  assign exp_734 = exp_590[2:2];
  assign exp_824 = 4;
  assign exp_833 = exp_643 & exp_595;
  assign exp_643 = exp_627 == exp_642;

      reg [5:0] exp_627_reg = 0;
      always@(posedge clk) begin
        if (exp_621) begin
          exp_627_reg <= exp_634;
        end
      end
      assign exp_627 = exp_627_reg;
    
  reg [5:0] exp_634_reg;
  always@(*) begin
    case (exp_629)
      0:exp_634_reg <= exp_631;
      1:exp_634_reg <= exp_632;
      default:exp_634_reg <= exp_633;
    endcase
  end
  assign exp_634 = exp_634_reg;
  assign exp_629 = exp_627 == exp_628;
  assign exp_628 = 37;
  assign exp_633 = 0;
  assign exp_631 = exp_627 + exp_630;
  assign exp_630 = 1;
  assign exp_632 = 0;
  assign exp_642 = 37;

      reg [0:0] exp_255_reg = 0;
      always@(posedge clk) begin
        if (exp_247) begin
          exp_255_reg <= exp_254;
        end
      end
      assign exp_255 = exp_255_reg;
      assign exp_254 = exp_252 & exp_253;

      reg [0:0] exp_252_reg = 0;
      always@(posedge clk) begin
        if (exp_247) begin
          exp_252_reg <= exp_251;
        end
      end
      assign exp_252 = exp_252_reg;
      assign exp_251 = exp_249 & exp_250;
  assign exp_249 = 1;
  assign exp_250 = ~exp_248;
  assign exp_248 = exp_860;
  assign exp_860 = exp_255 & exp_552;
  assign exp_247 = ~exp_246;
  assign exp_246 = exp_864;
  assign exp_864 = exp_255 & exp_863;
  assign exp_863 = exp_862 | exp_838;
  assign exp_862 = exp_243 & exp_861;
  assign exp_861 = ~exp_242;
  assign exp_242 = exp_233;

  reg [0:0] exp_233_reg;
  always@(*) begin
    case (exp_228)
      0:exp_233_reg <= exp_211;
      1:exp_233_reg <= exp_220;
      default:exp_233_reg <= exp_232;
    endcase
  end
  assign exp_233 = exp_233_reg;
  assign exp_228 = exp_225 & exp_227;
  assign exp_225 = exp_1 >= exp_224;
  assign exp_1 = exp_239;
  assign exp_239 = exp_446;
  assign exp_446 = exp_445 + exp_444;
  assign exp_445 = 0;
  assign exp_444 = exp_367 + exp_443;
  assign exp_443 = $signed(exp_442);
  assign exp_442 = exp_441 + exp_440;
  assign exp_441 = 0;

  reg [11:0] exp_440_reg;
  always@(*) begin
    case (exp_394)
      0:exp_440_reg <= exp_435;
      1:exp_440_reg <= exp_438;
      default:exp_440_reg <= exp_439;
    endcase
  end
  assign exp_440 = exp_440_reg;
  assign exp_394 = exp_377 == exp_393;
  assign exp_393 = 35;
  assign exp_439 = 0;
  assign exp_435 = exp_375[31:20];
  assign exp_438 = {exp_436, exp_437};  assign exp_436 = exp_375[31:25];
  assign exp_437 = exp_375[11:7];
  assign exp_224 = 34359738380;
  assign exp_227 = exp_1 <= exp_226;
  assign exp_226 = 34359738380;
  assign exp_232 = 0;

  reg [0:0] exp_211_reg;
  always@(*) begin
    case (exp_206)
      0:exp_211_reg <= exp_177;
      1:exp_211_reg <= exp_198;
      default:exp_211_reg <= exp_210;
    endcase
  end
  assign exp_211 = exp_211_reg;
  assign exp_206 = exp_203 & exp_205;
  assign exp_203 = exp_1 >= exp_202;
  assign exp_202 = 34359738376;
  assign exp_205 = exp_1 <= exp_204;
  assign exp_204 = 34359738376;
  assign exp_210 = 0;

  reg [0:0] exp_177_reg;
  always@(*) begin
    case (exp_172)
      0:exp_177_reg <= exp_155;
      1:exp_177_reg <= exp_164;
      default:exp_177_reg <= exp_176;
    endcase
  end
  assign exp_177 = exp_177_reg;
  assign exp_172 = exp_169 & exp_171;
  assign exp_169 = exp_1 >= exp_168;
  assign exp_168 = 2147483648;
  assign exp_171 = exp_1 <= exp_170;
  assign exp_170 = 2147483652;
  assign exp_176 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 305419896;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 305419896;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 16380;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_244;
  assign exp_244 = exp_529;
  assign exp_529 = exp_528 + exp_394;
  assign exp_528 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_157;
  assign exp_157 = debug_ready_in;
  assign exp_164 = exp_189;
  assign exp_189 = 1;
  assign exp_198 = exp_213;
  assign exp_213 = stdout_ready_in;
  assign exp_220 = exp_235;
  assign exp_235 = spare_ready_in;
  assign exp_838 = exp_595 & exp_837;
  assign exp_837 = ~exp_835;
  assign exp_253 = ~exp_248;
  assign exp_296 = 0;

  //Create RAM
  reg [31:0] exp_268_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_266) begin
      exp_268_ram[exp_262] <= exp_264;
    end
  end
  assign exp_268 = exp_268_ram[exp_263];
  assign exp_267 = exp_276;
  assign exp_276 = 1;
  assign exp_263 = exp_260;
  assign exp_266 = exp_844;
  assign exp_844 = exp_843 & exp_247;
  assign exp_843 = exp_841 & exp_255;
  assign exp_262 = exp_842;
  assign exp_264 = exp_840;

  reg [31:0] exp_840_reg;
  always@(*) begin
    case (exp_836)
      0:exp_840_reg <= exp_477;
      1:exp_840_reg <= exp_831;
      default:exp_840_reg <= exp_839;
    endcase
  end
  assign exp_840 = exp_840_reg;
  assign exp_839 = 0;

  reg [31:0] exp_477_reg;
  always@(*) begin
    case (exp_392)
      0:exp_477_reg <= exp_428;
      1:exp_477_reg <= exp_475;
      default:exp_477_reg <= exp_476;
    endcase
  end
  assign exp_477 = exp_477_reg;
  assign exp_476 = 0;

  reg [31:0] exp_428_reg;
  always@(*) begin
    case (exp_371)
      0:exp_428_reg <= exp_407;
      1:exp_428_reg <= exp_409;
      2:exp_428_reg <= exp_425;
      3:exp_428_reg <= exp_426;
      4:exp_428_reg <= exp_418;
      5:exp_428_reg <= exp_422;
      6:exp_428_reg <= exp_423;
      7:exp_428_reg <= exp_424;
      default:exp_428_reg <= exp_427;
    endcase
  end
  assign exp_428 = exp_428_reg;

      reg [2:0] exp_371_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_371_reg <= exp_362;
        end
      end
      assign exp_371 = exp_371_reg;
    
  reg [2:0] exp_362_reg;
  always@(*) begin
    case (exp_359)
      0:exp_362_reg <= exp_349;
      1:exp_362_reg <= exp_360;
      default:exp_362_reg <= exp_361;
    endcase
  end
  assign exp_362 = exp_362_reg;
  assign exp_359 = exp_293 | exp_295;
  assign exp_293 = exp_283 == exp_292;
  assign exp_283 = exp_96[6:0];
  assign exp_292 = 111;
  assign exp_295 = exp_283 == exp_294;
  assign exp_294 = 103;
  assign exp_361 = 0;

  reg [2:0] exp_349_reg;
  always@(*) begin
    case (exp_291)
      0:exp_349_reg <= exp_336;
      1:exp_349_reg <= exp_347;
      default:exp_349_reg <= exp_348;
    endcase
  end
  assign exp_349 = exp_349_reg;
  assign exp_291 = exp_283 == exp_290;
  assign exp_290 = 23;
  assign exp_348 = 0;

  reg [2:0] exp_336_reg;
  always@(*) begin
    case (exp_289)
      0:exp_336_reg <= exp_285;
      1:exp_336_reg <= exp_334;
      default:exp_336_reg <= exp_335;
    endcase
  end
  assign exp_336 = exp_336_reg;
  assign exp_289 = exp_283 == exp_288;
  assign exp_288 = 55;
  assign exp_335 = 0;
  assign exp_285 = exp_96[14:12];
  assign exp_334 = 0;
  assign exp_347 = 0;
  assign exp_360 = 0;
  assign exp_366 = exp_247 & exp_252;
  assign exp_427 = 0;

  reg [31:0] exp_407_reg;
  always@(*) begin
    case (exp_373)
      0:exp_407_reg <= exp_404;
      1:exp_407_reg <= exp_405;
      default:exp_407_reg <= exp_406;
    endcase
  end
  assign exp_407 = exp_407_reg;

      reg [0:0] exp_373_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_373_reg <= exp_365;
        end
      end
      assign exp_373 = exp_373_reg;
      assign exp_365 = exp_351 & exp_364;
  assign exp_351 = exp_338 & exp_350;
  assign exp_338 = exp_324 & exp_337;
  assign exp_324 = exp_322 & exp_323;
  assign exp_322 = exp_96[30:30];
  assign exp_323 = ~exp_287;
  assign exp_287 = exp_283 == exp_286;
  assign exp_286 = 19;
  assign exp_337 = ~exp_289;
  assign exp_350 = ~exp_291;
  assign exp_364 = ~exp_363;
  assign exp_363 = exp_293 | exp_295;
  assign exp_406 = 0;
  assign exp_404 = exp_369 + exp_370;

      reg [31:0] exp_369_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_369_reg <= exp_355;
        end
      end
      assign exp_369 = exp_369_reg;
    
  reg [31:0] exp_355_reg;
  always@(*) begin
    case (exp_352)
      0:exp_355_reg <= exp_344;
      1:exp_355_reg <= exp_353;
      default:exp_355_reg <= exp_354;
    endcase
  end
  assign exp_355 = exp_355_reg;
  assign exp_352 = exp_293 | exp_295;
  assign exp_354 = 0;

  reg [31:0] exp_344_reg;
  always@(*) begin
    case (exp_291)
      0:exp_344_reg <= exp_330;
      1:exp_344_reg <= exp_342;
      default:exp_344_reg <= exp_343;
    endcase
  end
  assign exp_344 = exp_344_reg;
  assign exp_343 = 0;

  reg [31:0] exp_330_reg;
  always@(*) begin
    case (exp_289)
      0:exp_330_reg <= exp_305;
      1:exp_330_reg <= exp_328;
      default:exp_330_reg <= exp_329;
    endcase
  end
  assign exp_330 = exp_330_reg;
  assign exp_329 = 0;
  assign exp_328 = exp_326 << exp_327;
  assign exp_326 = exp_325;
  assign exp_325 = exp_96[31:12];
  assign exp_327 = 12;
  assign exp_342 = exp_340 << exp_341;
  assign exp_340 = exp_339;
  assign exp_339 = exp_96[31:12];
  assign exp_341 = 12;
  assign exp_353 = 4;

      reg [31:0] exp_370_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_370_reg <= exp_358;
        end
      end
      assign exp_370 = exp_370_reg;
    
  reg [31:0] exp_358_reg;
  always@(*) begin
    case (exp_356)
      0:exp_358_reg <= exp_346;
      1:exp_358_reg <= exp_259;
      default:exp_358_reg <= exp_357;
    endcase
  end
  assign exp_358 = exp_358_reg;
  assign exp_356 = exp_293 | exp_295;
  assign exp_357 = 0;

  reg [31:0] exp_346_reg;
  always@(*) begin
    case (exp_291)
      0:exp_346_reg <= exp_333;
      1:exp_346_reg <= exp_259;
      default:exp_346_reg <= exp_345;
    endcase
  end
  assign exp_346 = exp_346_reg;
  assign exp_345 = 0;

  reg [31:0] exp_333_reg;
  always@(*) begin
    case (exp_289)
      0:exp_333_reg <= exp_317;
      1:exp_333_reg <= exp_331;
      default:exp_333_reg <= exp_332;
    endcase
  end
  assign exp_333 = exp_333_reg;
  assign exp_332 = 0;

  reg [31:0] exp_317_reg;
  always@(*) begin
    case (exp_287)
      0:exp_317_reg <= exp_311;
      1:exp_317_reg <= exp_315;
      default:exp_317_reg <= exp_316;
    endcase
  end
  assign exp_317 = exp_317_reg;
  assign exp_316 = 0;

  reg [31:0] exp_311_reg;
  always@(*) begin
    case (exp_307)
      0:exp_311_reg <= exp_299;
      1:exp_311_reg <= exp_309;
      default:exp_311_reg <= exp_310;
    endcase
  end
  assign exp_311 = exp_311_reg;
  assign exp_307 = exp_282 == exp_306;
  assign exp_282 = exp_96[24:20];
  assign exp_306 = 0;
  assign exp_310 = 0;

  reg [31:0] exp_299_reg;
  always@(*) begin
    case (exp_279)
      0:exp_299_reg <= exp_275;
      1:exp_299_reg <= exp_280;
      default:exp_299_reg <= exp_298;
    endcase
  end
  assign exp_299 = exp_299_reg;
  assign exp_279 = exp_854;
  assign exp_854 = exp_853 & exp_247;
  assign exp_853 = exp_852 & exp_255;
  assign exp_852 = exp_851 & exp_841;
  assign exp_851 = exp_261 == exp_842;
  assign exp_261 = exp_96[24:20];
  assign exp_298 = 0;

  //Create RAM
  reg [31:0] exp_275_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_273) begin
      exp_275_ram[exp_269] <= exp_271;
    end
  end
  assign exp_275 = exp_275_ram[exp_270];
  assign exp_274 = exp_277;
  assign exp_277 = 1;
  assign exp_270 = exp_261;
  assign exp_273 = exp_846;
  assign exp_846 = exp_845 & exp_247;
  assign exp_845 = exp_841 & exp_255;
  assign exp_269 = exp_842;
  assign exp_271 = exp_840;
  assign exp_280 = exp_840;
  assign exp_309 = $signed(exp_308);
  assign exp_308 = 0;
  assign exp_315 = exp_312 + exp_314;
  assign exp_312 = 0;
  assign exp_314 = $signed(exp_313);
  assign exp_313 = exp_96[31:20];
  assign exp_331 = 0;

      reg [31:0] exp_259_reg = 0;
      always@(posedge clk) begin
        if (exp_258) begin
          exp_259_reg <= exp_257;
        end
      end
      assign exp_259 = exp_259_reg;
      assign exp_258 = exp_249 & exp_247;
  assign exp_405 = exp_369 - exp_370;
  assign exp_409 = exp_369 << exp_408;
  assign exp_408 = $signed(exp_403);
  assign exp_403 = exp_402 + exp_401;
  assign exp_402 = 0;
  assign exp_401 = exp_372;

      reg [4:0] exp_372_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_372_reg <= exp_321;
        end
      end
      assign exp_372 = exp_372_reg;
    
  reg [4:0] exp_321_reg;
  always@(*) begin
    case (exp_287)
      0:exp_321_reg <= exp_319;
      1:exp_321_reg <= exp_284;
      default:exp_321_reg <= exp_320;
    endcase
  end
  assign exp_321 = exp_321_reg;
  assign exp_320 = 0;
  assign exp_319 = exp_317[4:0];
  assign exp_284 = exp_96[24:20];
  assign exp_425 = $signed(exp_411);
  assign exp_411 = exp_410;
  assign exp_410 = $signed(exp_369) < $signed(exp_370);
  assign exp_426 = $signed(exp_417);
  assign exp_417 = exp_416;
  assign exp_416 = exp_413 < exp_415;
  assign exp_413 = exp_412 + exp_369;
  assign exp_412 = 0;
  assign exp_415 = exp_414 + exp_370;
  assign exp_414 = 0;
  assign exp_418 = exp_369 ^ exp_370;
  assign exp_422 = exp_421[31:0];
  assign exp_421 = $signed(exp_419) >>> $signed(exp_420);
  assign exp_419 = {exp_400, exp_369};
  reg [0:0] exp_400_reg;
  always@(*) begin
    case (exp_374)
      0:exp_400_reg <= exp_398;
      1:exp_400_reg <= exp_397;
      default:exp_400_reg <= exp_399;
    endcase
  end
  assign exp_400 = exp_400_reg;

      reg [0:0] exp_374_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_374_reg <= exp_318;
        end
      end
      assign exp_374 = exp_374_reg;
      assign exp_318 = exp_96[30:30];
  assign exp_399 = 0;
  assign exp_398 = 0;
  assign exp_397 = exp_369[31:31];
  assign exp_420 = $signed(exp_403);
  assign exp_423 = exp_369 | exp_370;
  assign exp_424 = exp_369 & exp_370;

  reg [31:0] exp_475_reg;
  always@(*) begin
    case (exp_378)
      0:exp_475_reg <= exp_465;
      1:exp_475_reg <= exp_468;
      2:exp_475_reg <= exp_241;
      3:exp_475_reg <= exp_469;
      4:exp_475_reg <= exp_470;
      5:exp_475_reg <= exp_471;
      6:exp_475_reg <= exp_472;
      7:exp_475_reg <= exp_473;
      default:exp_475_reg <= exp_474;
    endcase
  end
  assign exp_475 = exp_475_reg;
  assign exp_474 = 0;
  assign exp_465 = $signed(exp_464);
  assign exp_464 = exp_463 + exp_458;
  assign exp_463 = 0;

  reg [7:0] exp_458_reg;
  always@(*) begin
    case (exp_449)
      0:exp_458_reg <= exp_453;
      1:exp_458_reg <= exp_454;
      2:exp_458_reg <= exp_455;
      3:exp_458_reg <= exp_456;
      default:exp_458_reg <= exp_457;
    endcase
  end
  assign exp_458 = exp_458_reg;
  assign exp_449 = exp_448 + exp_447;
  assign exp_448 = 0;
  assign exp_447 = exp_446[1:0];
  assign exp_457 = 0;
  assign exp_453 = exp_241[7:0];
  assign exp_241 = exp_231;

  reg [31:0] exp_231_reg;
  always@(*) begin
    case (exp_228)
      0:exp_231_reg <= exp_209;
      1:exp_231_reg <= exp_219;
      default:exp_231_reg <= exp_230;
    endcase
  end
  assign exp_231 = exp_231_reg;
  assign exp_230 = 0;

  reg [31:0] exp_209_reg;
  always@(*) begin
    case (exp_206)
      0:exp_209_reg <= exp_175;
      1:exp_209_reg <= exp_197;
      default:exp_209_reg <= exp_208;
    endcase
  end
  assign exp_209 = exp_209_reg;
  assign exp_208 = 0;

  reg [31:0] exp_175_reg;
  always@(*) begin
    case (exp_172)
      0:exp_175_reg <= exp_153;
      1:exp_175_reg <= exp_163;
      default:exp_175_reg <= exp_174;
    endcase
  end
  assign exp_175 = exp_175_reg;
  assign exp_174 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 127;
    exp_54_ram[32] = 3;
    exp_54_ram[33] = 0;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 0;
    exp_54_ram[36] = 0;
    exp_54_ram[37] = 0;
    exp_54_ram[38] = 0;
    exp_54_ram[39] = 0;
    exp_54_ram[40] = 0;
    exp_54_ram[41] = 0;
    exp_54_ram[42] = 254;
    exp_54_ram[43] = 128;
    exp_54_ram[44] = 0;
    exp_54_ram[45] = 253;
    exp_54_ram[46] = 12;
    exp_54_ram[47] = 255;
    exp_54_ram[48] = 108;
    exp_54_ram[49] = 111;
    exp_54_ram[50] = 33;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_245;
  assign exp_245 = exp_526;

  reg [3:0] exp_526_reg;
  always@(*) begin
    case (exp_378)
      0:exp_526_reg <= exp_513;
      1:exp_526_reg <= exp_518;
      2:exp_526_reg <= exp_519;
      3:exp_526_reg <= exp_520;
      4:exp_526_reg <= exp_521;
      5:exp_526_reg <= exp_522;
      6:exp_526_reg <= exp_523;
      7:exp_526_reg <= exp_524;
      default:exp_526_reg <= exp_525;
    endcase
  end
  assign exp_526 = exp_526_reg;
  assign exp_525 = 0;
  assign exp_513 = exp_509 << exp_512;
  assign exp_509 = 1;
  assign exp_512 = exp_511 + exp_510;
  assign exp_511 = 0;
  assign exp_510 = exp_446[1:0];
  assign exp_518 = exp_514 << exp_517;
  assign exp_514 = 3;
  assign exp_517 = exp_516 + exp_515;
  assign exp_516 = 0;
  assign exp_515 = exp_446[1:1];
  assign exp_519 = 15;
  assign exp_520 = 0;
  assign exp_521 = 0;
  assign exp_522 = 0;
  assign exp_523 = 0;
  assign exp_524 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_240;
  assign exp_240 = exp_508;

  reg [31:0] exp_508_reg;
  always@(*) begin
    case (exp_378)
      0:exp_508_reg <= exp_495;
      1:exp_508_reg <= exp_499;
      2:exp_508_reg <= exp_501;
      3:exp_508_reg <= exp_502;
      4:exp_508_reg <= exp_503;
      5:exp_508_reg <= exp_504;
      6:exp_508_reg <= exp_505;
      7:exp_508_reg <= exp_506;
      default:exp_508_reg <= exp_507;
    endcase
  end
  assign exp_508 = exp_508_reg;
  assign exp_507 = 0;

  reg [31:0] exp_495_reg;
  always@(*) begin
    case (exp_449)
      0:exp_495_reg <= exp_481;
      1:exp_495_reg <= exp_489;
      2:exp_495_reg <= exp_491;
      3:exp_495_reg <= exp_493;
      default:exp_495_reg <= exp_494;
    endcase
  end
  assign exp_495 = exp_495_reg;
  assign exp_494 = 0;
  assign exp_481 = exp_480;
  assign exp_480 = exp_479 + exp_478;
  assign exp_479 = 0;
  assign exp_478 = exp_368[7:0];

      reg [31:0] exp_368_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_368_reg <= exp_311;
        end
      end
      assign exp_368 = exp_368_reg;
      assign exp_489 = exp_481 << exp_488;
  assign exp_488 = 8;
  assign exp_491 = exp_481 << exp_490;
  assign exp_490 = 16;
  assign exp_493 = exp_481 << exp_492;
  assign exp_492 = 24;

  reg [31:0] exp_499_reg;
  always@(*) begin
    case (exp_452)
      0:exp_499_reg <= exp_485;
      1:exp_499_reg <= exp_497;
      default:exp_499_reg <= exp_498;
    endcase
  end
  assign exp_499 = exp_499_reg;
  assign exp_452 = exp_451 + exp_450;
  assign exp_451 = 0;
  assign exp_450 = exp_446[1:1];
  assign exp_498 = 0;
  assign exp_485 = exp_484;
  assign exp_484 = exp_483 + exp_482;
  assign exp_483 = 0;
  assign exp_482 = exp_368[15:0];
  assign exp_497 = exp_485 << exp_496;
  assign exp_496 = 16;
  assign exp_501 = exp_500 + exp_487;
  assign exp_500 = 0;
  assign exp_487 = exp_486 + exp_368;
  assign exp_486 = 0;
  assign exp_502 = 0;
  assign exp_503 = 0;
  assign exp_504 = 0;
  assign exp_505 = 0;
  assign exp_506 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 192;
    exp_47_ram[32] = 128;
    exp_47_ram[33] = 0;
    exp_47_ram[34] = 5;
    exp_47_ram[35] = 0;
    exp_47_ram[36] = 167;
    exp_47_ram[37] = 7;
    exp_47_ram[38] = 7;
    exp_47_ram[39] = 0;
    exp_47_ram[40] = 21;
    exp_47_ram[41] = 229;
    exp_47_ram[42] = 159;
    exp_47_ram[43] = 0;
    exp_47_ram[44] = 133;
    exp_47_ram[45] = 95;
    exp_47_ram[46] = 0;
    exp_47_ram[47] = 31;
    exp_47_ram[48] = 108;
    exp_47_ram[49] = 87;
    exp_47_ram[50] = 100;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 1;
    exp_40_ram[32] = 0;
    exp_40_ram[33] = 0;
    exp_40_ram[34] = 7;
    exp_40_ram[35] = 5;
    exp_40_ram[36] = 135;
    exp_40_ram[37] = 71;
    exp_40_ram[38] = 20;
    exp_40_ram[39] = 128;
    exp_40_ram[40] = 5;
    exp_40_ram[41] = 160;
    exp_40_ram[42] = 240;
    exp_40_ram[43] = 5;
    exp_40_ram[44] = 133;
    exp_40_ram[45] = 240;
    exp_40_ram[46] = 5;
    exp_40_ram[47] = 240;
    exp_40_ram[48] = 101;
    exp_40_ram[49] = 32;
    exp_40_ram[50] = 108;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 19;
    exp_33_ram[32] = 239;
    exp_33_ram[33] = 111;
    exp_33_ram[34] = 147;
    exp_33_ram[35] = 19;
    exp_33_ram[36] = 51;
    exp_33_ram[37] = 3;
    exp_33_ram[38] = 99;
    exp_33_ram[39] = 103;
    exp_33_ram[40] = 19;
    exp_33_ram[41] = 35;
    exp_33_ram[42] = 111;
    exp_33_ram[43] = 183;
    exp_33_ram[44] = 147;
    exp_33_ram[45] = 111;
    exp_33_ram[46] = 19;
    exp_33_ram[47] = 111;
    exp_33_ram[48] = 72;
    exp_33_ram[49] = 111;
    exp_33_ram[50] = 114;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_160;
  assign exp_160 = 0;
  assign exp_163 = exp_194;

  reg [31:0] exp_194_reg;
  always@(*) begin
    case (exp_190)
      0:exp_194_reg <= exp_191;
      1:exp_194_reg <= exp_192;
      default:exp_194_reg <= exp_193;
    endcase
  end
  assign exp_194 = exp_194_reg;
  assign exp_190 = exp_161[2:2];
  assign exp_161 = exp_1;
  assign exp_193 = 0;
  assign exp_191 = exp_179[31:0];

      reg [63:0] exp_179_reg = 0;
      always@(posedge clk) begin
        if (exp_178) begin
          exp_179_reg <= exp_186;
        end
      end
      assign exp_179 = exp_179_reg;
    
  reg [63:0] exp_186_reg;
  always@(*) begin
    case (exp_181)
      0:exp_186_reg <= exp_183;
      1:exp_186_reg <= exp_184;
      default:exp_186_reg <= exp_185;
    endcase
  end
  assign exp_186 = exp_186_reg;
  assign exp_181 = exp_179 == exp_180;
  assign exp_180 = 18446744073709551616;
  assign exp_185 = 0;
  assign exp_183 = exp_179 + exp_182;
  assign exp_182 = 1;
  assign exp_184 = 0;
  assign exp_178 = 1;
  assign exp_192 = exp_179[63:32];
  assign exp_197 = exp_216;
  assign exp_216 = 0;
  assign exp_219 = exp_238;
  assign exp_238 = 0;
  assign exp_454 = exp_241[15:8];
  assign exp_455 = exp_241[23:16];
  assign exp_456 = exp_241[31:24];
  assign exp_468 = $signed(exp_467);
  assign exp_467 = exp_466 + exp_462;
  assign exp_466 = 0;

  reg [15:0] exp_462_reg;
  always@(*) begin
    case (exp_452)
      0:exp_462_reg <= exp_459;
      1:exp_462_reg <= exp_460;
      default:exp_462_reg <= exp_461;
    endcase
  end
  assign exp_462 = exp_462_reg;
  assign exp_461 = 0;
  assign exp_459 = exp_241[15:0];
  assign exp_460 = exp_241[31:16];
  assign exp_469 = 0;
  assign exp_470 = exp_458;
  assign exp_471 = exp_462;
  assign exp_472 = 0;
  assign exp_473 = 0;

  reg [31:0] exp_831_reg;
  always@(*) begin
    case (exp_621)
      0:exp_831_reg <= exp_827;
      1:exp_831_reg <= exp_829;
      default:exp_831_reg <= exp_830;
    endcase
  end
  assign exp_831 = exp_831_reg;
  assign exp_830 = 0;

  reg [31:0] exp_827_reg;
  always@(*) begin
    case (exp_598)
      0:exp_827_reg <= exp_822;
      1:exp_827_reg <= exp_823;
      default:exp_827_reg <= exp_826;
    endcase
  end
  assign exp_827 = exp_827_reg;
  assign exp_598 = exp_597 & exp_595;
  assign exp_597 = exp_590 == exp_596;
  assign exp_596 = 0;
  assign exp_826 = 0;
  assign exp_822 = exp_821[63:32];

  reg [63:0] exp_821_reg;
  always@(*) begin
    case (exp_818)
      0:exp_821_reg <= exp_817;
      1:exp_821_reg <= exp_819;
      default:exp_821_reg <= exp_820;
    endcase
  end
  assign exp_821 = exp_821_reg;

      reg [0:0] exp_818_reg = 0;
      always@(posedge clk) begin
        if (exp_803) begin
          exp_818_reg <= exp_801;
        end
      end
      assign exp_818 = exp_818_reg;
    
      reg [0:0] exp_801_reg = 0;
      always@(posedge clk) begin
        if (exp_780) begin
          exp_801_reg <= exp_778;
        end
      end
      assign exp_801 = exp_801_reg;
    
      reg [0:0] exp_778_reg = 0;
      always@(posedge clk) begin
        if (exp_760) begin
          exp_778_reg <= exp_775;
        end
      end
      assign exp_778 = exp_778_reg;
      assign exp_775 = exp_773 ^ exp_774;
  assign exp_773 = exp_755 & exp_738;
  assign exp_755 = exp_754 + exp_753;
  assign exp_754 = 0;
  assign exp_753 = exp_751[31:31];

      reg [31:0] exp_751_reg = 0;
      always@(posedge clk) begin
        if (exp_750) begin
          exp_751_reg <= exp_369;
        end
      end
      assign exp_751 = exp_751_reg;
      assign exp_750 = exp_740 == exp_749;
  assign exp_749 = 0;
  assign exp_738 = exp_737 | exp_604;
  assign exp_737 = exp_598 | exp_601;
  assign exp_601 = exp_600 & exp_595;
  assign exp_600 = exp_590 == exp_599;
  assign exp_599 = 1;
  assign exp_604 = exp_603 & exp_595;
  assign exp_603 = exp_590 == exp_602;
  assign exp_602 = 2;
  assign exp_774 = exp_758 & exp_739;
  assign exp_758 = exp_757 + exp_756;
  assign exp_757 = 0;
  assign exp_756 = exp_752[31:31];

      reg [31:0] exp_752_reg = 0;
      always@(posedge clk) begin
        if (exp_750) begin
          exp_752_reg <= exp_370;
        end
      end
      assign exp_752 = exp_752_reg;
      assign exp_739 = exp_598 | exp_601;
  assign exp_760 = exp_740 == exp_759;
  assign exp_759 = 1;
  assign exp_780 = exp_740 == exp_779;
  assign exp_779 = 2;
  assign exp_803 = exp_740 == exp_802;
  assign exp_802 = 3;
  assign exp_820 = 0;

      reg [63:0] exp_817_reg = 0;
      always@(posedge clk) begin
        if (exp_803) begin
          exp_817_reg <= exp_816;
        end
      end
      assign exp_817 = exp_817_reg;
      assign exp_816 = exp_812 + exp_815;
  assign exp_812 = exp_808 + exp_811;
  assign exp_808 = exp_804 + exp_807;
  assign exp_804 = exp_797;

      reg [31:0] exp_797_reg = 0;
      always@(posedge clk) begin
        if (exp_780) begin
          exp_797_reg <= exp_784;
        end
      end
      assign exp_797 = exp_797_reg;
      assign exp_784 = exp_782 * exp_783;
  assign exp_782 = exp_781;
  assign exp_781 = exp_776[15:0];

      reg [31:0] exp_776_reg = 0;
      always@(posedge clk) begin
        if (exp_760) begin
          exp_776_reg <= exp_766;
        end
      end
      assign exp_776 = exp_776_reg;
      assign exp_766 = exp_765 + exp_764;
  assign exp_765 = 0;

  reg [31:0] exp_764_reg;
  always@(*) begin
    case (exp_761)
      0:exp_764_reg <= exp_751;
      1:exp_764_reg <= exp_762;
      default:exp_764_reg <= exp_763;
    endcase
  end
  assign exp_764 = exp_764_reg;
  assign exp_761 = exp_755 & exp_738;
  assign exp_763 = 0;
  assign exp_762 = -exp_751;
  assign exp_783 = exp_777[15:0];

      reg [31:0] exp_777_reg = 0;
      always@(posedge clk) begin
        if (exp_760) begin
          exp_777_reg <= exp_772;
        end
      end
      assign exp_777 = exp_777_reg;
      assign exp_772 = exp_771 + exp_770;
  assign exp_771 = 0;

  reg [31:0] exp_770_reg;
  always@(*) begin
    case (exp_767)
      0:exp_770_reg <= exp_752;
      1:exp_770_reg <= exp_768;
      default:exp_770_reg <= exp_769;
    endcase
  end
  assign exp_770 = exp_770_reg;
  assign exp_767 = exp_758 & exp_739;
  assign exp_769 = 0;
  assign exp_768 = -exp_752;
  assign exp_807 = exp_805 << exp_806;
  assign exp_805 = exp_798;

      reg [31:0] exp_798_reg = 0;
      always@(posedge clk) begin
        if (exp_780) begin
          exp_798_reg <= exp_788;
        end
      end
      assign exp_798 = exp_798_reg;
      assign exp_788 = exp_786 * exp_787;
  assign exp_786 = exp_785;
  assign exp_785 = exp_776[15:0];
  assign exp_787 = exp_777[31:16];
  assign exp_806 = 16;
  assign exp_811 = exp_809 << exp_810;
  assign exp_809 = exp_799;

      reg [31:0] exp_799_reg = 0;
      always@(posedge clk) begin
        if (exp_780) begin
          exp_799_reg <= exp_792;
        end
      end
      assign exp_799 = exp_799_reg;
      assign exp_792 = exp_790 * exp_791;
  assign exp_790 = exp_789;
  assign exp_789 = exp_776[31:16];
  assign exp_791 = exp_777[15:0];
  assign exp_810 = 16;
  assign exp_815 = exp_813 << exp_814;
  assign exp_813 = exp_800;

      reg [31:0] exp_800_reg = 0;
      always@(posedge clk) begin
        if (exp_780) begin
          exp_800_reg <= exp_796;
        end
      end
      assign exp_800 = exp_800_reg;
      assign exp_796 = exp_794 * exp_795;
  assign exp_794 = exp_793;
  assign exp_793 = exp_776[31:16];
  assign exp_795 = exp_777[31:16];
  assign exp_814 = 32;
  assign exp_819 = -exp_817;
  assign exp_823 = exp_821[31:0];

  reg [31:0] exp_829_reg;
  always@(*) begin
    case (exp_622)
      0:exp_829_reg <= exp_732;
      1:exp_829_reg <= exp_733;
      default:exp_829_reg <= exp_828;
    endcase
  end
  assign exp_829 = exp_829_reg;
  assign exp_622 = exp_590[1:1];
  assign exp_828 = 0;

      reg [31:0] exp_732_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_732_reg <= exp_726;
        end
      end
      assign exp_732 = exp_732_reg;
    
  reg [31:0] exp_726_reg;
  always@(*) begin
    case (exp_722)
      0:exp_726_reg <= exp_713;
      1:exp_726_reg <= exp_724;
      default:exp_726_reg <= exp_725;
    endcase
  end
  assign exp_726 = exp_726_reg;
  assign exp_722 = exp_721 & exp_624;
  assign exp_721 = exp_670 == exp_720;

      reg [31:0] exp_670_reg = 0;
      always@(posedge clk) begin
        if (exp_655) begin
          exp_670_reg <= exp_667;
        end
      end
      assign exp_670 = exp_670_reg;
      assign exp_667 = exp_666 + exp_665;
  assign exp_666 = 0;

  reg [31:0] exp_665_reg;
  always@(*) begin
    case (exp_662)
      0:exp_665_reg <= exp_647;
      1:exp_665_reg <= exp_663;
      default:exp_665_reg <= exp_664;
    endcase
  end
  assign exp_665 = exp_665_reg;
  assign exp_662 = exp_653 & exp_624;
  assign exp_653 = exp_652 + exp_651;
  assign exp_652 = 0;
  assign exp_651 = exp_647[31:31];

      reg [31:0] exp_647_reg = 0;
      always@(posedge clk) begin
        if (exp_645) begin
          exp_647_reg <= exp_370;
        end
      end
      assign exp_647 = exp_647_reg;
      assign exp_645 = exp_627 == exp_644;
  assign exp_644 = 0;
  assign exp_624 = ~exp_623;
  assign exp_623 = exp_590[0:0];
  assign exp_664 = 0;
  assign exp_663 = -exp_647;
  assign exp_655 = exp_627 == exp_654;
  assign exp_654 = 1;
  assign exp_720 = 0;
  assign exp_725 = 0;
  assign exp_713 = exp_712 + exp_711;
  assign exp_712 = 0;

  reg [31:0] exp_711_reg;
  always@(*) begin
    case (exp_708)
      0:exp_711_reg <= exp_706;
      1:exp_711_reg <= exp_709;
      default:exp_711_reg <= exp_710;
    endcase
  end
  assign exp_711 = exp_711_reg;
  assign exp_708 = exp_672 & exp_624;

      reg [0:0] exp_672_reg = 0;
      always@(posedge clk) begin
        if (exp_655) begin
          exp_672_reg <= exp_668;
        end
      end
      assign exp_672 = exp_672_reg;
      assign exp_668 = exp_650 ^ exp_653;
  assign exp_650 = exp_649 + exp_648;
  assign exp_649 = 0;
  assign exp_648 = exp_646[31:31];

      reg [31:0] exp_646_reg = 0;
      always@(posedge clk) begin
        if (exp_645) begin
          exp_646_reg <= exp_369;
        end
      end
      assign exp_646 = exp_646_reg;
      assign exp_710 = 0;

      reg [31:0] exp_706_reg = 0;
      always@(posedge clk) begin
        if (exp_639) begin
          exp_706_reg <= exp_676;
        end
      end
      assign exp_706 = exp_706_reg;
    
      reg [31:0] exp_676_reg = 0;
      always@(posedge clk) begin
        if (exp_675) begin
          exp_676_reg <= exp_703;
        end
      end
      assign exp_676 = exp_676_reg;
    
  reg [31:0] exp_703_reg;
  always@(*) begin
    case (exp_637)
      0:exp_703_reg <= exp_695;
      1:exp_703_reg <= exp_701;
      default:exp_703_reg <= exp_702;
    endcase
  end
  assign exp_703 = exp_703_reg;
  assign exp_637 = exp_627 == exp_636;
  assign exp_636 = 2;
  assign exp_702 = 0;

  reg [31:0] exp_695_reg;
  always@(*) begin
    case (exp_685)
      0:exp_695_reg <= exp_689;
      1:exp_695_reg <= exp_693;
      default:exp_695_reg <= exp_694;
    endcase
  end
  assign exp_695 = exp_695_reg;
  assign exp_685 = ~exp_684;
  assign exp_684 = exp_683[32:32];
  assign exp_683 = exp_682 - exp_670;
  assign exp_682 = exp_681;
  assign exp_681 = {exp_679, exp_680};  assign exp_679 = exp_674[31:0];

      reg [31:0] exp_674_reg = 0;
      always@(posedge clk) begin
        if (exp_673) begin
          exp_674_reg <= exp_700;
        end
      end
      assign exp_674 = exp_674_reg;
    
  reg [32:0] exp_700_reg;
  always@(*) begin
    case (exp_637)
      0:exp_700_reg <= exp_687;
      1:exp_700_reg <= exp_698;
      default:exp_700_reg <= exp_699;
    endcase
  end
  assign exp_700 = exp_700_reg;
  assign exp_699 = 0;

  reg [32:0] exp_687_reg;
  always@(*) begin
    case (exp_685)
      0:exp_687_reg <= exp_681;
      1:exp_687_reg <= exp_683;
      default:exp_687_reg <= exp_686;
    endcase
  end
  assign exp_687 = exp_687_reg;
  assign exp_686 = 0;
  assign exp_698 = 0;
  assign exp_673 = 1;
  assign exp_680 = exp_678[31:31];

      reg [31:0] exp_678_reg = 0;
      always@(posedge clk) begin
        if (exp_677) begin
          exp_678_reg <= exp_705;
        end
      end
      assign exp_678 = exp_678_reg;
    
  reg [31:0] exp_705_reg;
  always@(*) begin
    case (exp_637)
      0:exp_705_reg <= exp_697;
      1:exp_705_reg <= exp_669;
      default:exp_705_reg <= exp_704;
    endcase
  end
  assign exp_705 = exp_705_reg;
  assign exp_704 = 0;
  assign exp_697 = exp_678 << exp_696;
  assign exp_696 = 1;

      reg [31:0] exp_669_reg = 0;
      always@(posedge clk) begin
        if (exp_655) begin
          exp_669_reg <= exp_661;
        end
      end
      assign exp_669 = exp_669_reg;
      assign exp_661 = exp_660 + exp_659;
  assign exp_660 = 0;

  reg [31:0] exp_659_reg;
  always@(*) begin
    case (exp_656)
      0:exp_659_reg <= exp_646;
      1:exp_659_reg <= exp_657;
      default:exp_659_reg <= exp_658;
    endcase
  end
  assign exp_659 = exp_659_reg;
  assign exp_656 = exp_650 & exp_624;
  assign exp_658 = 0;
  assign exp_657 = -exp_646;
  assign exp_677 = 1;
  assign exp_694 = 0;
  assign exp_689 = exp_676 << exp_688;
  assign exp_688 = 1;
  assign exp_693 = exp_691 | exp_692;
  assign exp_691 = exp_676 << exp_690;
  assign exp_690 = 1;
  assign exp_692 = 1;
  assign exp_701 = 0;
  assign exp_675 = 1;
  assign exp_639 = exp_627 == exp_638;
  assign exp_638 = 35;
  assign exp_709 = -exp_706;
  assign exp_724 = $signed(exp_723);
  assign exp_723 = -1;
  assign exp_641 = exp_627 == exp_640;
  assign exp_640 = 36;

      reg [31:0] exp_733_reg = 0;
      always@(posedge clk) begin
        if (exp_641) begin
          exp_733_reg <= exp_731;
        end
      end
      assign exp_733 = exp_733_reg;
    
  reg [31:0] exp_731_reg;
  always@(*) begin
    case (exp_729)
      0:exp_731_reg <= exp_719;
      1:exp_731_reg <= exp_646;
      default:exp_731_reg <= exp_730;
    endcase
  end
  assign exp_731 = exp_731_reg;
  assign exp_729 = exp_728 & exp_624;
  assign exp_728 = exp_670 == exp_727;
  assign exp_727 = 0;
  assign exp_730 = 0;
  assign exp_719 = exp_718 + exp_717;
  assign exp_718 = 0;

  reg [31:0] exp_717_reg;
  always@(*) begin
    case (exp_714)
      0:exp_717_reg <= exp_707;
      1:exp_717_reg <= exp_715;
      default:exp_717_reg <= exp_716;
    endcase
  end
  assign exp_717 = exp_717_reg;
  assign exp_714 = exp_671 & exp_624;

      reg [0:0] exp_671_reg = 0;
      always@(posedge clk) begin
        if (exp_655) begin
          exp_671_reg <= exp_650;
        end
      end
      assign exp_671 = exp_671_reg;
      assign exp_716 = 0;

      reg [31:0] exp_707_reg = 0;
      always@(posedge clk) begin
        if (exp_639) begin
          exp_707_reg <= exp_674;
        end
      end
      assign exp_707 = exp_707_reg;
      assign exp_715 = -exp_707;
  assign exp_303 = $signed(exp_302);
  assign exp_302 = 0;
  assign exp_532 = exp_367 != exp_368;
  assign exp_545 = 0;
  assign exp_546 = 0;
  assign exp_533 = $signed(exp_367) < $signed(exp_368);
  assign exp_534 = $signed(exp_367) >= $signed(exp_368);
  assign exp_539 = exp_536 < exp_538;
  assign exp_536 = exp_535 + exp_367;
  assign exp_535 = 0;
  assign exp_538 = exp_537 + exp_368;
  assign exp_537 = 0;
  assign exp_544 = exp_541 >= exp_543;
  assign exp_541 = exp_540 + exp_367;
  assign exp_540 = 0;
  assign exp_543 = exp_542 + exp_368;
  assign exp_542 = 0;
  assign exp_858 = 0;
  assign exp_857 = exp_257 + exp_856;
  assign exp_856 = 4;

  reg [32:0] exp_589_reg;
  always@(*) begin
    case (exp_390)
      0:exp_589_reg <= exp_579;
      1:exp_589_reg <= exp_587;
      default:exp_589_reg <= exp_588;
    endcase
  end
  assign exp_589 = exp_589_reg;
  assign exp_588 = 0;
  assign exp_579 = exp_578 + exp_376;

  reg [31:0] exp_578_reg;
  always@(*) begin
    case (exp_388)
      0:exp_578_reg <= exp_564;
      1:exp_578_reg <= exp_576;
      default:exp_578_reg <= exp_577;
    endcase
  end
  assign exp_578 = exp_578_reg;
  assign exp_577 = 0;
  assign exp_564 = $signed(exp_563);
  assign exp_563 = exp_562 + exp_561;
  assign exp_562 = 0;
  assign exp_561 = {exp_560, exp_557};  assign exp_560 = {exp_559, exp_556};  assign exp_559 = {exp_558, exp_555};  assign exp_558 = {exp_553, exp_554};  assign exp_553 = exp_375[31:31];
  assign exp_554 = exp_375[7:7];
  assign exp_555 = exp_375[30:25];
  assign exp_556 = exp_375[11:8];
  assign exp_557 = 0;
  assign exp_576 = $signed(exp_575);
  assign exp_575 = exp_574 + exp_573;
  assign exp_574 = 0;
  assign exp_573 = {exp_572, exp_569};  assign exp_572 = {exp_571, exp_568};  assign exp_571 = {exp_570, exp_567};  assign exp_570 = {exp_565, exp_566};  assign exp_565 = exp_375[31:31];
  assign exp_566 = exp_375[19:12];
  assign exp_567 = exp_375[20:20];
  assign exp_568 = exp_375[30:21];
  assign exp_569 = 0;

      reg [31:0] exp_376_reg = 0;
      always@(posedge clk) begin
        if (exp_366) begin
          exp_376_reg <= exp_259;
        end
      end
      assign exp_376 = exp_376_reg;
      assign exp_587 = exp_586 & exp_585;
  assign exp_586 = $signed(exp_584);
  assign exp_584 = exp_367 + exp_583;
  assign exp_583 = $signed(exp_582);
  assign exp_582 = exp_581 + exp_580;
  assign exp_581 = 0;
  assign exp_580 = exp_375[31:20];
  assign exp_585 = 4294967294;
  assign exp_256 = exp_249 & exp_247;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_258;
  assign exp_391 = 3;
  assign exp_144 = exp_6;
  assign exp_140 = exp_2;
  assign exp_215 = exp_199 & exp_200;
  assign exp_199 = exp_207;
  assign exp_207 = exp_5 & exp_206;
  assign exp_200 = exp_6;
  assign exp_196 = exp_2;
  assign exp_237 = exp_221 & exp_222;
  assign exp_221 = exp_229;
  assign exp_229 = exp_5 & exp_228;
  assign exp_222 = exp_6;
  assign exp_218 = exp_2;
  assign debug_valid_out = exp_159;
  assign debug_out = exp_140;
  assign stdout_valid_out = exp_215;
  assign stdout_out = exp_196;
  assign spare_valid_out = exp_237;
  assign spare_out = exp_218;

endmodule