
module soc(clk, stdin_valid_in, stdin_in, stdout_ready_in, stdin_ready_out, stdout_valid_out, stdout_out, leds_out);
  input [0:0] stdin_valid_in;
  input [31:0] stdin_in;
  input [0:0] stdout_ready_in;
  input [0:0] clk;
  output [0:0] stdin_ready_out;
  output [0:0] stdout_valid_out;
  output [31:0] stdout_out;
  output [31:0] leds_out;
  wire [0:0] exp_245;
  wire [0:0] exp_228;
  wire [0:0] exp_236;
  wire [0:0] exp_5;
  wire [0:0] exp_250;
  wire [0:0] exp_597;
  wire [0:0] exp_534;
  wire [0:0] exp_399;
  wire [6:0] exp_384;
  wire [31:0] exp_382;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [11:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_264;
  wire [32:0] exp_867;
  wire [0:0] exp_863;
  wire [0:0] exp_559;
  wire [0:0] exp_537;
  wire [0:0] exp_395;
  wire [6:0] exp_394;
  wire [0:0] exp_397;
  wire [6:0] exp_396;
  wire [0:0] exp_558;
  wire [0:0] exp_403;
  wire [6:0] exp_402;
  wire [0:0] exp_557;
  wire [0:0] exp_556;
  wire [0:0] exp_555;
  wire [2:0] exp_385;
  wire [0:0] exp_554;
  wire [0:0] exp_538;
  wire [31:0] exp_374;
  wire [31:0] exp_312;
  wire [0:0] exp_308;
  wire [4:0] exp_288;
  wire [0:0] exp_307;
  wire [0:0] exp_311;
  wire [31:0] exp_304;
  wire [0:0] exp_285;
  wire [0:0] exp_858;
  wire [0:0] exp_857;
  wire [0:0] exp_856;
  wire [0:0] exp_855;
  wire [4:0] exp_267;
  wire [4:0] exp_850;
  wire [0:0] exp_849;
  wire [0:0] exp_441;
  wire [0:0] exp_440;
  wire [0:0] exp_439;
  wire [0:0] exp_438;
  wire [0:0] exp_437;
  wire [0:0] exp_436;
  wire [0:0] exp_387;
  wire [4:0] exp_386;
  wire [0:0] exp_389;
  wire [5:0] exp_388;
  wire [0:0] exp_391;
  wire [5:0] exp_390;
  wire [0:0] exp_393;
  wire [4:0] exp_392;
  wire [0:0] exp_844;
  wire [0:0] exp_843;
  wire [0:0] exp_629;
  wire [0:0] exp_603;
  wire [0:0] exp_601;
  wire [6:0] exp_599;
  wire [5:0] exp_600;
  wire [0:0] exp_602;
  wire [0:0] exp_628;
  wire [2:0] exp_598;
  wire [0:0] exp_842;
  wire [0:0] exp_840;
  wire [0:0] exp_833;
  wire [2:0] exp_748;
  wire [2:0] exp_755;
  wire [0:0] exp_750;
  wire [2:0] exp_749;
  wire [0:0] exp_754;
  wire [2:0] exp_752;
  wire [0:0] exp_751;
  wire [0:0] exp_753;
  wire [0:0] exp_744;
  wire [0:0] exp_743;
  wire [0:0] exp_742;
  wire [2:0] exp_832;
  wire [0:0] exp_841;
  wire [0:0] exp_651;
  wire [5:0] exp_635;
  wire [5:0] exp_642;
  wire [0:0] exp_637;
  wire [5:0] exp_636;
  wire [0:0] exp_641;
  wire [5:0] exp_639;
  wire [0:0] exp_638;
  wire [0:0] exp_640;
  wire [5:0] exp_650;
  wire [0:0] exp_262;
  wire [0:0] exp_261;
  wire [0:0] exp_259;
  wire [0:0] exp_258;
  wire [0:0] exp_256;
  wire [0:0] exp_257;
  wire [0:0] exp_255;
  wire [0:0] exp_868;
  wire [0:0] exp_254;
  wire [0:0] exp_253;
  wire [0:0] exp_872;
  wire [0:0] exp_871;
  wire [0:0] exp_870;
  wire [0:0] exp_869;
  wire [0:0] exp_249;
  wire [0:0] exp_240;
  wire [0:0] exp_235;
  wire [0:0] exp_232;
  wire [31:0] exp_1;
  wire [31:0] exp_246;
  wire [31:0] exp_453;
  wire [31:0] exp_452;
  wire [31:0] exp_451;
  wire [31:0] exp_450;
  wire [11:0] exp_449;
  wire [11:0] exp_448;
  wire [11:0] exp_447;
  wire [0:0] exp_401;
  wire [5:0] exp_400;
  wire [0:0] exp_446;
  wire [11:0] exp_442;
  wire [11:0] exp_445;
  wire [6:0] exp_443;
  wire [4:0] exp_444;
  wire [31:0] exp_231;
  wire [0:0] exp_234;
  wire [31:0] exp_233;
  wire [0:0] exp_239;
  wire [0:0] exp_218;
  wire [0:0] exp_213;
  wire [0:0] exp_210;
  wire [31:0] exp_209;
  wire [0:0] exp_212;
  wire [31:0] exp_211;
  wire [0:0] exp_217;
  wire [0:0] exp_196;
  wire [0:0] exp_191;
  wire [0:0] exp_188;
  wire [31:0] exp_187;
  wire [0:0] exp_190;
  wire [31:0] exp_189;
  wire [0:0] exp_195;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [31:0] exp_146;
  wire [0:0] exp_149;
  wire [31:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [13:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_251;
  wire [0:0] exp_536;
  wire [0:0] exp_535;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_176;
  wire [0:0] exp_183;
  wire [0:0] exp_198;
  wire [0:0] exp_205;
  wire [0:0] exp_223;
  wire [0:0] exp_227;
  wire [0:0] exp_243;
  wire [0:0] exp_846;
  wire [0:0] exp_845;
  wire [0:0] exp_260;
  wire [0:0] exp_303;
  wire [31:0] exp_275;
  wire [0:0] exp_274;
  wire [1:0] exp_283;
  wire [4:0] exp_270;
  wire [0:0] exp_273;
  wire [0:0] exp_852;
  wire [0:0] exp_851;
  wire [4:0] exp_269;
  wire [31:0] exp_271;
  wire [31:0] exp_848;
  wire [0:0] exp_847;
  wire [31:0] exp_484;
  wire [0:0] exp_483;
  wire [31:0] exp_435;
  wire [2:0] exp_378;
  wire [2:0] exp_369;
  wire [0:0] exp_366;
  wire [0:0] exp_300;
  wire [6:0] exp_290;
  wire [6:0] exp_299;
  wire [0:0] exp_302;
  wire [6:0] exp_301;
  wire [0:0] exp_368;
  wire [2:0] exp_356;
  wire [0:0] exp_298;
  wire [4:0] exp_297;
  wire [0:0] exp_355;
  wire [2:0] exp_343;
  wire [0:0] exp_296;
  wire [5:0] exp_295;
  wire [0:0] exp_342;
  wire [2:0] exp_292;
  wire [0:0] exp_341;
  wire [0:0] exp_354;
  wire [0:0] exp_367;
  wire [0:0] exp_373;
  wire [0:0] exp_434;
  wire [31:0] exp_414;
  wire [0:0] exp_380;
  wire [0:0] exp_372;
  wire [0:0] exp_358;
  wire [0:0] exp_345;
  wire [0:0] exp_331;
  wire [0:0] exp_329;
  wire [0:0] exp_330;
  wire [0:0] exp_294;
  wire [4:0] exp_293;
  wire [0:0] exp_344;
  wire [0:0] exp_357;
  wire [0:0] exp_371;
  wire [0:0] exp_370;
  wire [0:0] exp_413;
  wire [31:0] exp_411;
  wire [31:0] exp_376;
  wire [31:0] exp_362;
  wire [0:0] exp_359;
  wire [0:0] exp_361;
  wire [31:0] exp_351;
  wire [0:0] exp_350;
  wire [31:0] exp_337;
  wire [0:0] exp_336;
  wire [31:0] exp_335;
  wire [31:0] exp_333;
  wire [19:0] exp_332;
  wire [3:0] exp_334;
  wire [31:0] exp_349;
  wire [31:0] exp_347;
  wire [19:0] exp_346;
  wire [3:0] exp_348;
  wire [31:0] exp_360;
  wire [31:0] exp_377;
  wire [31:0] exp_365;
  wire [0:0] exp_363;
  wire [0:0] exp_364;
  wire [31:0] exp_353;
  wire [0:0] exp_352;
  wire [31:0] exp_340;
  wire [0:0] exp_339;
  wire [31:0] exp_324;
  wire [0:0] exp_323;
  wire [31:0] exp_318;
  wire [0:0] exp_314;
  wire [4:0] exp_289;
  wire [0:0] exp_313;
  wire [0:0] exp_317;
  wire [31:0] exp_306;
  wire [0:0] exp_286;
  wire [0:0] exp_862;
  wire [0:0] exp_861;
  wire [0:0] exp_860;
  wire [0:0] exp_859;
  wire [4:0] exp_268;
  wire [0:0] exp_305;
  wire [31:0] exp_282;
  wire [0:0] exp_281;
  wire [1:0] exp_284;
  wire [4:0] exp_277;
  wire [0:0] exp_280;
  wire [0:0] exp_854;
  wire [0:0] exp_853;
  wire [4:0] exp_276;
  wire [31:0] exp_278;
  wire [31:0] exp_287;
  wire [31:0] exp_316;
  wire [0:0] exp_315;
  wire [31:0] exp_322;
  wire [31:0] exp_319;
  wire [31:0] exp_321;
  wire [11:0] exp_320;
  wire [31:0] exp_338;
  wire [31:0] exp_266;
  wire [0:0] exp_265;
  wire [31:0] exp_412;
  wire [31:0] exp_416;
  wire [31:0] exp_415;
  wire [5:0] exp_410;
  wire [5:0] exp_409;
  wire [5:0] exp_408;
  wire [4:0] exp_379;
  wire [4:0] exp_328;
  wire [0:0] exp_327;
  wire [4:0] exp_326;
  wire [4:0] exp_291;
  wire [31:0] exp_432;
  wire [1:0] exp_418;
  wire [0:0] exp_417;
  wire [31:0] exp_433;
  wire [1:0] exp_424;
  wire [0:0] exp_423;
  wire [31:0] exp_420;
  wire [31:0] exp_419;
  wire [31:0] exp_422;
  wire [31:0] exp_421;
  wire [31:0] exp_425;
  wire [31:0] exp_429;
  wire [32:0] exp_428;
  wire [32:0] exp_426;
  wire [0:0] exp_407;
  wire [0:0] exp_381;
  wire [0:0] exp_325;
  wire [0:0] exp_406;
  wire [0:0] exp_405;
  wire [0:0] exp_404;
  wire [32:0] exp_427;
  wire [31:0] exp_430;
  wire [31:0] exp_431;
  wire [31:0] exp_482;
  wire [0:0] exp_481;
  wire [31:0] exp_472;
  wire [7:0] exp_471;
  wire [7:0] exp_470;
  wire [7:0] exp_465;
  wire [1:0] exp_456;
  wire [1:0] exp_455;
  wire [1:0] exp_454;
  wire [0:0] exp_464;
  wire [7:0] exp_460;
  wire [31:0] exp_248;
  wire [31:0] exp_238;
  wire [0:0] exp_237;
  wire [31:0] exp_216;
  wire [0:0] exp_215;
  wire [31:0] exp_194;
  wire [0:0] exp_193;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [11:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_252;
  wire [3:0] exp_533;
  wire [0:0] exp_532;
  wire [3:0] exp_520;
  wire [3:0] exp_516;
  wire [1:0] exp_519;
  wire [1:0] exp_518;
  wire [1:0] exp_517;
  wire [3:0] exp_525;
  wire [3:0] exp_521;
  wire [0:0] exp_524;
  wire [0:0] exp_523;
  wire [0:0] exp_522;
  wire [3:0] exp_526;
  wire [3:0] exp_527;
  wire [3:0] exp_528;
  wire [3:0] exp_529;
  wire [3:0] exp_530;
  wire [3:0] exp_531;
  wire [11:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_247;
  wire [31:0] exp_515;
  wire [0:0] exp_514;
  wire [31:0] exp_502;
  wire [0:0] exp_501;
  wire [31:0] exp_488;
  wire [7:0] exp_487;
  wire [7:0] exp_486;
  wire [7:0] exp_485;
  wire [31:0] exp_375;
  wire [31:0] exp_496;
  wire [3:0] exp_495;
  wire [31:0] exp_498;
  wire [4:0] exp_497;
  wire [31:0] exp_500;
  wire [4:0] exp_499;
  wire [31:0] exp_506;
  wire [0:0] exp_459;
  wire [0:0] exp_458;
  wire [0:0] exp_457;
  wire [0:0] exp_505;
  wire [31:0] exp_492;
  wire [15:0] exp_491;
  wire [15:0] exp_490;
  wire [15:0] exp_489;
  wire [31:0] exp_504;
  wire [4:0] exp_503;
  wire [31:0] exp_508;
  wire [31:0] exp_507;
  wire [31:0] exp_494;
  wire [31:0] exp_493;
  wire [31:0] exp_509;
  wire [31:0] exp_510;
  wire [31:0] exp_511;
  wire [31:0] exp_512;
  wire [31:0] exp_513;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [11:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [11:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [11:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [11:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [11:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [11:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [11:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [11:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [11:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [11:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [11:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [11:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_179;
  wire [0:0] exp_177;
  wire [31:0] exp_139;
  wire [0:0] exp_178;
  wire [31:0] exp_157;
  wire [31:0] exp_164;
  wire [0:0] exp_159;
  wire [31:0] exp_158;
  wire [0:0] exp_163;
  wire [31:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [31:0] exp_167;
  wire [31:0] exp_174;
  wire [0:0] exp_169;
  wire [31:0] exp_168;
  wire [0:0] exp_173;
  wire [31:0] exp_171;
  wire [0:0] exp_170;
  wire [0:0] exp_172;
  wire [0:0] exp_166;
  wire [0:0] exp_165;
  wire [31:0] exp_182;
  wire [31:0] exp_201;
  wire [31:0] exp_204;
  wire [31:0] exp_222;
  wire [31:0] exp_226;
  wire [31:0] exp_241;
  wire [7:0] exp_461;
  wire [7:0] exp_462;
  wire [7:0] exp_463;
  wire [31:0] exp_475;
  wire [15:0] exp_474;
  wire [15:0] exp_473;
  wire [15:0] exp_469;
  wire [0:0] exp_468;
  wire [15:0] exp_466;
  wire [15:0] exp_467;
  wire [31:0] exp_476;
  wire [31:0] exp_477;
  wire [31:0] exp_478;
  wire [31:0] exp_479;
  wire [31:0] exp_480;
  wire [31:0] exp_839;
  wire [0:0] exp_838;
  wire [31:0] exp_835;
  wire [0:0] exp_606;
  wire [0:0] exp_605;
  wire [0:0] exp_604;
  wire [0:0] exp_834;
  wire [31:0] exp_830;
  wire [63:0] exp_829;
  wire [0:0] exp_826;
  wire [0:0] exp_809;
  wire [0:0] exp_786;
  wire [0:0] exp_783;
  wire [0:0] exp_781;
  wire [0:0] exp_763;
  wire [0:0] exp_762;
  wire [0:0] exp_761;
  wire [31:0] exp_759;
  wire [0:0] exp_758;
  wire [0:0] exp_757;
  wire [0:0] exp_746;
  wire [0:0] exp_745;
  wire [0:0] exp_609;
  wire [0:0] exp_608;
  wire [0:0] exp_607;
  wire [0:0] exp_612;
  wire [0:0] exp_611;
  wire [1:0] exp_610;
  wire [0:0] exp_782;
  wire [0:0] exp_766;
  wire [0:0] exp_765;
  wire [0:0] exp_764;
  wire [31:0] exp_760;
  wire [0:0] exp_747;
  wire [0:0] exp_768;
  wire [0:0] exp_767;
  wire [0:0] exp_788;
  wire [1:0] exp_787;
  wire [0:0] exp_811;
  wire [1:0] exp_810;
  wire [0:0] exp_828;
  wire [63:0] exp_825;
  wire [63:0] exp_824;
  wire [63:0] exp_820;
  wire [63:0] exp_816;
  wire [63:0] exp_812;
  wire [31:0] exp_805;
  wire [31:0] exp_792;
  wire [31:0] exp_790;
  wire [15:0] exp_789;
  wire [31:0] exp_784;
  wire [31:0] exp_774;
  wire [31:0] exp_773;
  wire [31:0] exp_772;
  wire [0:0] exp_769;
  wire [0:0] exp_771;
  wire [31:0] exp_770;
  wire [15:0] exp_791;
  wire [31:0] exp_785;
  wire [31:0] exp_780;
  wire [31:0] exp_779;
  wire [31:0] exp_778;
  wire [0:0] exp_775;
  wire [0:0] exp_777;
  wire [31:0] exp_776;
  wire [63:0] exp_815;
  wire [63:0] exp_813;
  wire [31:0] exp_806;
  wire [31:0] exp_796;
  wire [31:0] exp_794;
  wire [15:0] exp_793;
  wire [15:0] exp_795;
  wire [4:0] exp_814;
  wire [63:0] exp_819;
  wire [63:0] exp_817;
  wire [31:0] exp_807;
  wire [31:0] exp_800;
  wire [31:0] exp_798;
  wire [15:0] exp_797;
  wire [15:0] exp_799;
  wire [4:0] exp_818;
  wire [63:0] exp_823;
  wire [63:0] exp_821;
  wire [31:0] exp_808;
  wire [31:0] exp_804;
  wire [31:0] exp_802;
  wire [15:0] exp_801;
  wire [15:0] exp_803;
  wire [5:0] exp_822;
  wire [63:0] exp_827;
  wire [31:0] exp_831;
  wire [31:0] exp_837;
  wire [0:0] exp_630;
  wire [0:0] exp_836;
  wire [31:0] exp_740;
  wire [31:0] exp_734;
  wire [0:0] exp_730;
  wire [0:0] exp_729;
  wire [31:0] exp_678;
  wire [31:0] exp_675;
  wire [31:0] exp_674;
  wire [31:0] exp_673;
  wire [0:0] exp_670;
  wire [0:0] exp_661;
  wire [0:0] exp_660;
  wire [0:0] exp_659;
  wire [31:0] exp_655;
  wire [0:0] exp_653;
  wire [0:0] exp_652;
  wire [0:0] exp_632;
  wire [0:0] exp_631;
  wire [0:0] exp_672;
  wire [31:0] exp_671;
  wire [0:0] exp_663;
  wire [0:0] exp_662;
  wire [0:0] exp_728;
  wire [0:0] exp_733;
  wire [31:0] exp_721;
  wire [31:0] exp_720;
  wire [31:0] exp_719;
  wire [0:0] exp_716;
  wire [0:0] exp_680;
  wire [0:0] exp_676;
  wire [0:0] exp_658;
  wire [0:0] exp_657;
  wire [0:0] exp_656;
  wire [31:0] exp_654;
  wire [0:0] exp_718;
  wire [31:0] exp_714;
  wire [31:0] exp_684;
  wire [31:0] exp_711;
  wire [0:0] exp_645;
  wire [1:0] exp_644;
  wire [0:0] exp_710;
  wire [31:0] exp_703;
  wire [0:0] exp_693;
  wire [0:0] exp_692;
  wire [32:0] exp_691;
  wire [32:0] exp_690;
  wire [32:0] exp_689;
  wire [31:0] exp_687;
  wire [31:0] exp_682;
  wire [32:0] exp_708;
  wire [0:0] exp_707;
  wire [32:0] exp_695;
  wire [0:0] exp_694;
  wire [0:0] exp_706;
  wire [0:0] exp_681;
  wire [0:0] exp_688;
  wire [31:0] exp_686;
  wire [31:0] exp_713;
  wire [0:0] exp_712;
  wire [31:0] exp_705;
  wire [0:0] exp_704;
  wire [31:0] exp_677;
  wire [31:0] exp_669;
  wire [31:0] exp_668;
  wire [31:0] exp_667;
  wire [0:0] exp_664;
  wire [0:0] exp_666;
  wire [31:0] exp_665;
  wire [0:0] exp_685;
  wire [0:0] exp_702;
  wire [31:0] exp_697;
  wire [0:0] exp_696;
  wire [31:0] exp_701;
  wire [31:0] exp_699;
  wire [0:0] exp_698;
  wire [0:0] exp_700;
  wire [0:0] exp_709;
  wire [0:0] exp_683;
  wire [0:0] exp_647;
  wire [5:0] exp_646;
  wire [31:0] exp_717;
  wire [31:0] exp_732;
  wire [0:0] exp_731;
  wire [0:0] exp_649;
  wire [5:0] exp_648;
  wire [31:0] exp_741;
  wire [31:0] exp_739;
  wire [0:0] exp_737;
  wire [0:0] exp_736;
  wire [0:0] exp_735;
  wire [0:0] exp_738;
  wire [31:0] exp_727;
  wire [31:0] exp_726;
  wire [31:0] exp_725;
  wire [0:0] exp_722;
  wire [0:0] exp_679;
  wire [0:0] exp_724;
  wire [31:0] exp_715;
  wire [31:0] exp_723;
  wire [31:0] exp_310;
  wire [0:0] exp_309;
  wire [0:0] exp_539;
  wire [0:0] exp_552;
  wire [0:0] exp_553;
  wire [0:0] exp_540;
  wire [0:0] exp_541;
  wire [0:0] exp_546;
  wire [31:0] exp_543;
  wire [31:0] exp_542;
  wire [31:0] exp_545;
  wire [31:0] exp_544;
  wire [0:0] exp_551;
  wire [31:0] exp_548;
  wire [31:0] exp_547;
  wire [31:0] exp_550;
  wire [31:0] exp_549;
  wire [0:0] exp_866;
  wire [31:0] exp_865;
  wire [2:0] exp_864;
  wire [32:0] exp_596;
  wire [0:0] exp_595;
  wire [31:0] exp_586;
  wire [31:0] exp_585;
  wire [0:0] exp_584;
  wire [31:0] exp_571;
  wire [12:0] exp_570;
  wire [12:0] exp_569;
  wire [12:0] exp_568;
  wire [11:0] exp_567;
  wire [7:0] exp_566;
  wire [1:0] exp_565;
  wire [0:0] exp_560;
  wire [0:0] exp_561;
  wire [5:0] exp_562;
  wire [3:0] exp_563;
  wire [0:0] exp_564;
  wire [31:0] exp_583;
  wire [20:0] exp_582;
  wire [20:0] exp_581;
  wire [20:0] exp_580;
  wire [19:0] exp_579;
  wire [9:0] exp_578;
  wire [8:0] exp_577;
  wire [0:0] exp_572;
  wire [7:0] exp_573;
  wire [0:0] exp_574;
  wire [9:0] exp_575;
  wire [0:0] exp_576;
  wire [31:0] exp_383;
  wire [32:0] exp_594;
  wire [32:0] exp_593;
  wire [31:0] exp_591;
  wire [31:0] exp_590;
  wire [11:0] exp_589;
  wire [11:0] exp_588;
  wire [11:0] exp_587;
  wire [32:0] exp_592;
  wire [0:0] exp_263;
  wire [0:0] exp_80;
  wire [11:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_398;
  wire [0:0] exp_244;
  wire [0:0] exp_229;
  wire [0:0] exp_200;
  wire [0:0] exp_184;
  wire [0:0] exp_192;
  wire [0:0] exp_185;
  wire [31:0] exp_181;
  wire [31:0] exp_221;
  wire [31:0] exp_203;
  wire [0:0] exp_220;
  wire [0:0] exp_206;
  wire [0:0] exp_214;
  wire [0:0] exp_207;

  assign exp_245 = exp_228 & exp_244;
  assign exp_228 = exp_236;
  assign exp_236 = exp_5 & exp_235;
  assign exp_5 = exp_250;
  assign exp_250 = exp_597;
  assign exp_597 = exp_534 & exp_262;
  assign exp_534 = exp_399 | exp_401;
  assign exp_399 = exp_384 == exp_398;
  assign exp_384 = exp_382[6:0];

      reg [31:0] exp_382_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_382_reg <= exp_96;
        end
      end
      assign exp_382 = exp_382_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_264;

      reg [31:0] exp_264_reg = 0;
      always@(posedge clk) begin
        if (exp_263) begin
          exp_264_reg <= exp_867;
        end
      end
      assign exp_264 = exp_264_reg;
    
  reg [32:0] exp_867_reg;
  always@(*) begin
    case (exp_863)
      0:exp_867_reg <= exp_865;
      1:exp_867_reg <= exp_596;
      default:exp_867_reg <= exp_866;
    endcase
  end
  assign exp_867 = exp_867_reg;
  assign exp_863 = exp_559 & exp_262;
  assign exp_559 = exp_537 | exp_558;
  assign exp_537 = exp_395 | exp_397;
  assign exp_395 = exp_384 == exp_394;
  assign exp_394 = 111;
  assign exp_397 = exp_384 == exp_396;
  assign exp_396 = 103;

  reg [0:0] exp_558_reg;
  always@(*) begin
    case (exp_403)
      0:exp_558_reg <= exp_556;
      1:exp_558_reg <= exp_555;
      default:exp_558_reg <= exp_557;
    endcase
  end
  assign exp_558 = exp_558_reg;
  assign exp_403 = exp_384 == exp_402;
  assign exp_402 = 99;
  assign exp_557 = 0;
  assign exp_556 = 0;

  reg [0:0] exp_555_reg;
  always@(*) begin
    case (exp_385)
      0:exp_555_reg <= exp_538;
      1:exp_555_reg <= exp_539;
      2:exp_555_reg <= exp_552;
      3:exp_555_reg <= exp_553;
      4:exp_555_reg <= exp_540;
      5:exp_555_reg <= exp_541;
      6:exp_555_reg <= exp_546;
      7:exp_555_reg <= exp_551;
      default:exp_555_reg <= exp_554;
    endcase
  end
  assign exp_555 = exp_555_reg;
  assign exp_385 = exp_382[14:12];
  assign exp_554 = 0;
  assign exp_538 = exp_374 == exp_375;

      reg [31:0] exp_374_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_374_reg <= exp_312;
        end
      end
      assign exp_374 = exp_374_reg;
    
  reg [31:0] exp_312_reg;
  always@(*) begin
    case (exp_308)
      0:exp_312_reg <= exp_304;
      1:exp_312_reg <= exp_310;
      default:exp_312_reg <= exp_311;
    endcase
  end
  assign exp_312 = exp_312_reg;
  assign exp_308 = exp_288 == exp_307;
  assign exp_288 = exp_96[19:15];
  assign exp_307 = 0;
  assign exp_311 = 0;

  reg [31:0] exp_304_reg;
  always@(*) begin
    case (exp_285)
      0:exp_304_reg <= exp_275;
      1:exp_304_reg <= exp_287;
      default:exp_304_reg <= exp_303;
    endcase
  end
  assign exp_304 = exp_304_reg;
  assign exp_285 = exp_858;
  assign exp_858 = exp_857 & exp_254;
  assign exp_857 = exp_856 & exp_262;
  assign exp_856 = exp_855 & exp_849;
  assign exp_855 = exp_267 == exp_850;
  assign exp_267 = exp_96[19:15];
  assign exp_850 = exp_382[11:7];
  assign exp_849 = exp_441 | exp_844;
  assign exp_441 = exp_440 | exp_399;
  assign exp_440 = exp_439 | exp_393;
  assign exp_439 = exp_438 | exp_391;
  assign exp_438 = exp_437 | exp_397;
  assign exp_437 = exp_436 | exp_395;
  assign exp_436 = exp_387 | exp_389;
  assign exp_387 = exp_384 == exp_386;
  assign exp_386 = 19;
  assign exp_389 = exp_384 == exp_388;
  assign exp_388 = 51;
  assign exp_391 = exp_384 == exp_390;
  assign exp_390 = 55;
  assign exp_393 = exp_384 == exp_392;
  assign exp_392 = 23;
  assign exp_844 = exp_843 & exp_603;

  reg [0:0] exp_843_reg;
  always@(*) begin
    case (exp_629)
      0:exp_843_reg <= exp_840;
      1:exp_843_reg <= exp_841;
      default:exp_843_reg <= exp_842;
    endcase
  end
  assign exp_843 = exp_843_reg;
  assign exp_629 = exp_603 & exp_628;
  assign exp_603 = exp_601 & exp_602;
  assign exp_601 = exp_599 == exp_600;
  assign exp_599 = exp_382[6:0];
  assign exp_600 = 51;
  assign exp_602 = exp_382[25:25];
  assign exp_628 = exp_598[2:2];
  assign exp_598 = exp_382[14:12];
  assign exp_842 = 0;
  assign exp_840 = exp_833 & exp_603;
  assign exp_833 = exp_748 == exp_832;

      reg [2:0] exp_748_reg = 0;
      always@(posedge clk) begin
        if (exp_744) begin
          exp_748_reg <= exp_755;
        end
      end
      assign exp_748 = exp_748_reg;
    
  reg [2:0] exp_755_reg;
  always@(*) begin
    case (exp_750)
      0:exp_755_reg <= exp_752;
      1:exp_755_reg <= exp_753;
      default:exp_755_reg <= exp_754;
    endcase
  end
  assign exp_755 = exp_755_reg;
  assign exp_750 = exp_748 == exp_749;
  assign exp_749 = 4;
  assign exp_754 = 0;
  assign exp_752 = exp_748 + exp_751;
  assign exp_751 = 1;
  assign exp_753 = 0;
  assign exp_744 = exp_603 & exp_743;
  assign exp_743 = ~exp_742;
  assign exp_742 = exp_598[2:2];
  assign exp_832 = 4;
  assign exp_841 = exp_651 & exp_603;
  assign exp_651 = exp_635 == exp_650;

      reg [5:0] exp_635_reg = 0;
      always@(posedge clk) begin
        if (exp_629) begin
          exp_635_reg <= exp_642;
        end
      end
      assign exp_635 = exp_635_reg;
    
  reg [5:0] exp_642_reg;
  always@(*) begin
    case (exp_637)
      0:exp_642_reg <= exp_639;
      1:exp_642_reg <= exp_640;
      default:exp_642_reg <= exp_641;
    endcase
  end
  assign exp_642 = exp_642_reg;
  assign exp_637 = exp_635 == exp_636;
  assign exp_636 = 37;
  assign exp_641 = 0;
  assign exp_639 = exp_635 + exp_638;
  assign exp_638 = 1;
  assign exp_640 = 0;
  assign exp_650 = 37;

      reg [0:0] exp_262_reg = 0;
      always@(posedge clk) begin
        if (exp_254) begin
          exp_262_reg <= exp_261;
        end
      end
      assign exp_262 = exp_262_reg;
      assign exp_261 = exp_259 & exp_260;

      reg [0:0] exp_259_reg = 0;
      always@(posedge clk) begin
        if (exp_254) begin
          exp_259_reg <= exp_258;
        end
      end
      assign exp_259 = exp_259_reg;
      assign exp_258 = exp_256 & exp_257;
  assign exp_256 = 1;
  assign exp_257 = ~exp_255;
  assign exp_255 = exp_868;
  assign exp_868 = exp_262 & exp_559;
  assign exp_254 = ~exp_253;
  assign exp_253 = exp_872;
  assign exp_872 = exp_262 & exp_871;
  assign exp_871 = exp_870 | exp_846;
  assign exp_870 = exp_250 & exp_869;
  assign exp_869 = ~exp_249;
  assign exp_249 = exp_240;

  reg [0:0] exp_240_reg;
  always@(*) begin
    case (exp_235)
      0:exp_240_reg <= exp_218;
      1:exp_240_reg <= exp_227;
      default:exp_240_reg <= exp_239;
    endcase
  end
  assign exp_240 = exp_240_reg;
  assign exp_235 = exp_232 & exp_234;
  assign exp_232 = exp_1 >= exp_231;
  assign exp_1 = exp_246;
  assign exp_246 = exp_453;
  assign exp_453 = exp_452 + exp_451;
  assign exp_452 = 0;
  assign exp_451 = exp_374 + exp_450;
  assign exp_450 = $signed(exp_449);
  assign exp_449 = exp_448 + exp_447;
  assign exp_448 = 0;

  reg [11:0] exp_447_reg;
  always@(*) begin
    case (exp_401)
      0:exp_447_reg <= exp_442;
      1:exp_447_reg <= exp_445;
      default:exp_447_reg <= exp_446;
    endcase
  end
  assign exp_447 = exp_447_reg;
  assign exp_401 = exp_384 == exp_400;
  assign exp_400 = 35;
  assign exp_446 = 0;
  assign exp_442 = exp_382[31:20];
  assign exp_445 = {exp_443, exp_444};  assign exp_443 = exp_382[31:25];
  assign exp_444 = exp_382[11:7];
  assign exp_231 = 2147483664;
  assign exp_234 = exp_1 <= exp_233;
  assign exp_233 = 2147483664;
  assign exp_239 = 0;

  reg [0:0] exp_218_reg;
  always@(*) begin
    case (exp_213)
      0:exp_218_reg <= exp_196;
      1:exp_218_reg <= exp_205;
      default:exp_218_reg <= exp_217;
    endcase
  end
  assign exp_218 = exp_218_reg;
  assign exp_213 = exp_210 & exp_212;
  assign exp_210 = exp_1 >= exp_209;
  assign exp_209 = 2147483660;
  assign exp_212 = exp_1 <= exp_211;
  assign exp_211 = 2147483660;
  assign exp_217 = 0;

  reg [0:0] exp_196_reg;
  always@(*) begin
    case (exp_191)
      0:exp_196_reg <= exp_155;
      1:exp_196_reg <= exp_183;
      default:exp_196_reg <= exp_195;
    endcase
  end
  assign exp_196 = exp_196_reg;
  assign exp_191 = exp_188 & exp_190;
  assign exp_188 = exp_1 >= exp_187;
  assign exp_187 = 2147483656;
  assign exp_190 = exp_1 <= exp_189;
  assign exp_189 = 2147483656;
  assign exp_195 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 2147483648;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 2147483652;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 16380;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_251;
  assign exp_251 = exp_536;
  assign exp_536 = exp_535 + exp_401;
  assign exp_535 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_176;
  assign exp_176 = 1;
  assign exp_183 = exp_198;
  assign exp_198 = stdout_ready_in;
  assign exp_205 = exp_223;
  assign exp_223 = 1;
  assign exp_227 = exp_243;
  assign exp_243 = stdin_valid_in;
  assign exp_846 = exp_603 & exp_845;
  assign exp_845 = ~exp_843;
  assign exp_260 = ~exp_255;
  assign exp_303 = 0;

  //Create RAM
  reg [31:0] exp_275_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_273) begin
      exp_275_ram[exp_269] <= exp_271;
    end
  end
  assign exp_275 = exp_275_ram[exp_270];
  assign exp_274 = exp_283;
  assign exp_283 = 1;
  assign exp_270 = exp_267;
  assign exp_273 = exp_852;
  assign exp_852 = exp_851 & exp_254;
  assign exp_851 = exp_849 & exp_262;
  assign exp_269 = exp_850;
  assign exp_271 = exp_848;

  reg [31:0] exp_848_reg;
  always@(*) begin
    case (exp_844)
      0:exp_848_reg <= exp_484;
      1:exp_848_reg <= exp_839;
      default:exp_848_reg <= exp_847;
    endcase
  end
  assign exp_848 = exp_848_reg;
  assign exp_847 = 0;

  reg [31:0] exp_484_reg;
  always@(*) begin
    case (exp_399)
      0:exp_484_reg <= exp_435;
      1:exp_484_reg <= exp_482;
      default:exp_484_reg <= exp_483;
    endcase
  end
  assign exp_484 = exp_484_reg;
  assign exp_483 = 0;

  reg [31:0] exp_435_reg;
  always@(*) begin
    case (exp_378)
      0:exp_435_reg <= exp_414;
      1:exp_435_reg <= exp_416;
      2:exp_435_reg <= exp_432;
      3:exp_435_reg <= exp_433;
      4:exp_435_reg <= exp_425;
      5:exp_435_reg <= exp_429;
      6:exp_435_reg <= exp_430;
      7:exp_435_reg <= exp_431;
      default:exp_435_reg <= exp_434;
    endcase
  end
  assign exp_435 = exp_435_reg;

      reg [2:0] exp_378_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_378_reg <= exp_369;
        end
      end
      assign exp_378 = exp_378_reg;
    
  reg [2:0] exp_369_reg;
  always@(*) begin
    case (exp_366)
      0:exp_369_reg <= exp_356;
      1:exp_369_reg <= exp_367;
      default:exp_369_reg <= exp_368;
    endcase
  end
  assign exp_369 = exp_369_reg;
  assign exp_366 = exp_300 | exp_302;
  assign exp_300 = exp_290 == exp_299;
  assign exp_290 = exp_96[6:0];
  assign exp_299 = 111;
  assign exp_302 = exp_290 == exp_301;
  assign exp_301 = 103;
  assign exp_368 = 0;

  reg [2:0] exp_356_reg;
  always@(*) begin
    case (exp_298)
      0:exp_356_reg <= exp_343;
      1:exp_356_reg <= exp_354;
      default:exp_356_reg <= exp_355;
    endcase
  end
  assign exp_356 = exp_356_reg;
  assign exp_298 = exp_290 == exp_297;
  assign exp_297 = 23;
  assign exp_355 = 0;

  reg [2:0] exp_343_reg;
  always@(*) begin
    case (exp_296)
      0:exp_343_reg <= exp_292;
      1:exp_343_reg <= exp_341;
      default:exp_343_reg <= exp_342;
    endcase
  end
  assign exp_343 = exp_343_reg;
  assign exp_296 = exp_290 == exp_295;
  assign exp_295 = 55;
  assign exp_342 = 0;
  assign exp_292 = exp_96[14:12];
  assign exp_341 = 0;
  assign exp_354 = 0;
  assign exp_367 = 0;
  assign exp_373 = exp_254 & exp_259;
  assign exp_434 = 0;

  reg [31:0] exp_414_reg;
  always@(*) begin
    case (exp_380)
      0:exp_414_reg <= exp_411;
      1:exp_414_reg <= exp_412;
      default:exp_414_reg <= exp_413;
    endcase
  end
  assign exp_414 = exp_414_reg;

      reg [0:0] exp_380_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_380_reg <= exp_372;
        end
      end
      assign exp_380 = exp_380_reg;
      assign exp_372 = exp_358 & exp_371;
  assign exp_358 = exp_345 & exp_357;
  assign exp_345 = exp_331 & exp_344;
  assign exp_331 = exp_329 & exp_330;
  assign exp_329 = exp_96[30:30];
  assign exp_330 = ~exp_294;
  assign exp_294 = exp_290 == exp_293;
  assign exp_293 = 19;
  assign exp_344 = ~exp_296;
  assign exp_357 = ~exp_298;
  assign exp_371 = ~exp_370;
  assign exp_370 = exp_300 | exp_302;
  assign exp_413 = 0;
  assign exp_411 = exp_376 + exp_377;

      reg [31:0] exp_376_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_376_reg <= exp_362;
        end
      end
      assign exp_376 = exp_376_reg;
    
  reg [31:0] exp_362_reg;
  always@(*) begin
    case (exp_359)
      0:exp_362_reg <= exp_351;
      1:exp_362_reg <= exp_360;
      default:exp_362_reg <= exp_361;
    endcase
  end
  assign exp_362 = exp_362_reg;
  assign exp_359 = exp_300 | exp_302;
  assign exp_361 = 0;

  reg [31:0] exp_351_reg;
  always@(*) begin
    case (exp_298)
      0:exp_351_reg <= exp_337;
      1:exp_351_reg <= exp_349;
      default:exp_351_reg <= exp_350;
    endcase
  end
  assign exp_351 = exp_351_reg;
  assign exp_350 = 0;

  reg [31:0] exp_337_reg;
  always@(*) begin
    case (exp_296)
      0:exp_337_reg <= exp_312;
      1:exp_337_reg <= exp_335;
      default:exp_337_reg <= exp_336;
    endcase
  end
  assign exp_337 = exp_337_reg;
  assign exp_336 = 0;
  assign exp_335 = exp_333 << exp_334;
  assign exp_333 = exp_332;
  assign exp_332 = exp_96[31:12];
  assign exp_334 = 12;
  assign exp_349 = exp_347 << exp_348;
  assign exp_347 = exp_346;
  assign exp_346 = exp_96[31:12];
  assign exp_348 = 12;
  assign exp_360 = 4;

      reg [31:0] exp_377_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_377_reg <= exp_365;
        end
      end
      assign exp_377 = exp_377_reg;
    
  reg [31:0] exp_365_reg;
  always@(*) begin
    case (exp_363)
      0:exp_365_reg <= exp_353;
      1:exp_365_reg <= exp_266;
      default:exp_365_reg <= exp_364;
    endcase
  end
  assign exp_365 = exp_365_reg;
  assign exp_363 = exp_300 | exp_302;
  assign exp_364 = 0;

  reg [31:0] exp_353_reg;
  always@(*) begin
    case (exp_298)
      0:exp_353_reg <= exp_340;
      1:exp_353_reg <= exp_266;
      default:exp_353_reg <= exp_352;
    endcase
  end
  assign exp_353 = exp_353_reg;
  assign exp_352 = 0;

  reg [31:0] exp_340_reg;
  always@(*) begin
    case (exp_296)
      0:exp_340_reg <= exp_324;
      1:exp_340_reg <= exp_338;
      default:exp_340_reg <= exp_339;
    endcase
  end
  assign exp_340 = exp_340_reg;
  assign exp_339 = 0;

  reg [31:0] exp_324_reg;
  always@(*) begin
    case (exp_294)
      0:exp_324_reg <= exp_318;
      1:exp_324_reg <= exp_322;
      default:exp_324_reg <= exp_323;
    endcase
  end
  assign exp_324 = exp_324_reg;
  assign exp_323 = 0;

  reg [31:0] exp_318_reg;
  always@(*) begin
    case (exp_314)
      0:exp_318_reg <= exp_306;
      1:exp_318_reg <= exp_316;
      default:exp_318_reg <= exp_317;
    endcase
  end
  assign exp_318 = exp_318_reg;
  assign exp_314 = exp_289 == exp_313;
  assign exp_289 = exp_96[24:20];
  assign exp_313 = 0;
  assign exp_317 = 0;

  reg [31:0] exp_306_reg;
  always@(*) begin
    case (exp_286)
      0:exp_306_reg <= exp_282;
      1:exp_306_reg <= exp_287;
      default:exp_306_reg <= exp_305;
    endcase
  end
  assign exp_306 = exp_306_reg;
  assign exp_286 = exp_862;
  assign exp_862 = exp_861 & exp_254;
  assign exp_861 = exp_860 & exp_262;
  assign exp_860 = exp_859 & exp_849;
  assign exp_859 = exp_268 == exp_850;
  assign exp_268 = exp_96[24:20];
  assign exp_305 = 0;

  //Create RAM
  reg [31:0] exp_282_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_280) begin
      exp_282_ram[exp_276] <= exp_278;
    end
  end
  assign exp_282 = exp_282_ram[exp_277];
  assign exp_281 = exp_284;
  assign exp_284 = 1;
  assign exp_277 = exp_268;
  assign exp_280 = exp_854;
  assign exp_854 = exp_853 & exp_254;
  assign exp_853 = exp_849 & exp_262;
  assign exp_276 = exp_850;
  assign exp_278 = exp_848;
  assign exp_287 = exp_848;
  assign exp_316 = $signed(exp_315);
  assign exp_315 = 0;
  assign exp_322 = exp_319 + exp_321;
  assign exp_319 = 0;
  assign exp_321 = $signed(exp_320);
  assign exp_320 = exp_96[31:20];
  assign exp_338 = 0;

      reg [31:0] exp_266_reg = 0;
      always@(posedge clk) begin
        if (exp_265) begin
          exp_266_reg <= exp_264;
        end
      end
      assign exp_266 = exp_266_reg;
      assign exp_265 = exp_256 & exp_254;
  assign exp_412 = exp_376 - exp_377;
  assign exp_416 = exp_376 << exp_415;
  assign exp_415 = $signed(exp_410);
  assign exp_410 = exp_409 + exp_408;
  assign exp_409 = 0;
  assign exp_408 = exp_379;

      reg [4:0] exp_379_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_379_reg <= exp_328;
        end
      end
      assign exp_379 = exp_379_reg;
    
  reg [4:0] exp_328_reg;
  always@(*) begin
    case (exp_294)
      0:exp_328_reg <= exp_326;
      1:exp_328_reg <= exp_291;
      default:exp_328_reg <= exp_327;
    endcase
  end
  assign exp_328 = exp_328_reg;
  assign exp_327 = 0;
  assign exp_326 = exp_324[4:0];
  assign exp_291 = exp_96[24:20];
  assign exp_432 = $signed(exp_418);
  assign exp_418 = exp_417;
  assign exp_417 = $signed(exp_376) < $signed(exp_377);
  assign exp_433 = $signed(exp_424);
  assign exp_424 = exp_423;
  assign exp_423 = exp_420 < exp_422;
  assign exp_420 = exp_419 + exp_376;
  assign exp_419 = 0;
  assign exp_422 = exp_421 + exp_377;
  assign exp_421 = 0;
  assign exp_425 = exp_376 ^ exp_377;
  assign exp_429 = exp_428[31:0];
  assign exp_428 = $signed(exp_426) >>> $signed(exp_427);
  assign exp_426 = {exp_407, exp_376};
  reg [0:0] exp_407_reg;
  always@(*) begin
    case (exp_381)
      0:exp_407_reg <= exp_405;
      1:exp_407_reg <= exp_404;
      default:exp_407_reg <= exp_406;
    endcase
  end
  assign exp_407 = exp_407_reg;

      reg [0:0] exp_381_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_381_reg <= exp_325;
        end
      end
      assign exp_381 = exp_381_reg;
      assign exp_325 = exp_96[30:30];
  assign exp_406 = 0;
  assign exp_405 = 0;
  assign exp_404 = exp_376[31:31];
  assign exp_427 = $signed(exp_410);
  assign exp_430 = exp_376 | exp_377;
  assign exp_431 = exp_376 & exp_377;

  reg [31:0] exp_482_reg;
  always@(*) begin
    case (exp_385)
      0:exp_482_reg <= exp_472;
      1:exp_482_reg <= exp_475;
      2:exp_482_reg <= exp_248;
      3:exp_482_reg <= exp_476;
      4:exp_482_reg <= exp_477;
      5:exp_482_reg <= exp_478;
      6:exp_482_reg <= exp_479;
      7:exp_482_reg <= exp_480;
      default:exp_482_reg <= exp_481;
    endcase
  end
  assign exp_482 = exp_482_reg;
  assign exp_481 = 0;
  assign exp_472 = $signed(exp_471);
  assign exp_471 = exp_470 + exp_465;
  assign exp_470 = 0;

  reg [7:0] exp_465_reg;
  always@(*) begin
    case (exp_456)
      0:exp_465_reg <= exp_460;
      1:exp_465_reg <= exp_461;
      2:exp_465_reg <= exp_462;
      3:exp_465_reg <= exp_463;
      default:exp_465_reg <= exp_464;
    endcase
  end
  assign exp_465 = exp_465_reg;
  assign exp_456 = exp_455 + exp_454;
  assign exp_455 = 0;
  assign exp_454 = exp_453[1:0];
  assign exp_464 = 0;
  assign exp_460 = exp_248[7:0];
  assign exp_248 = exp_238;

  reg [31:0] exp_238_reg;
  always@(*) begin
    case (exp_235)
      0:exp_238_reg <= exp_216;
      1:exp_238_reg <= exp_226;
      default:exp_238_reg <= exp_237;
    endcase
  end
  assign exp_238 = exp_238_reg;
  assign exp_237 = 0;

  reg [31:0] exp_216_reg;
  always@(*) begin
    case (exp_213)
      0:exp_216_reg <= exp_194;
      1:exp_216_reg <= exp_204;
      default:exp_216_reg <= exp_215;
    endcase
  end
  assign exp_216 = exp_216_reg;
  assign exp_215 = 0;

  reg [31:0] exp_194_reg;
  always@(*) begin
    case (exp_191)
      0:exp_194_reg <= exp_153;
      1:exp_194_reg <= exp_182;
      default:exp_194_reg <= exp_193;
    endcase
  end
  assign exp_194 = exp_194_reg;
  assign exp_193 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 0;
    exp_54_ram[32] = 255;
    exp_54_ram[33] = 125;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 0;
    exp_54_ram[36] = 0;
    exp_54_ram[37] = 0;
    exp_54_ram[38] = 0;
    exp_54_ram[39] = 0;
    exp_54_ram[40] = 40;
    exp_54_ram[41] = 0;
    exp_54_ram[42] = 188;
    exp_54_ram[43] = 14;
    exp_54_ram[44] = 0;
    exp_54_ram[45] = 12;
    exp_54_ram[46] = 15;
    exp_54_ram[47] = 0;
    exp_54_ram[48] = 0;
    exp_54_ram[49] = 0;
    exp_54_ram[50] = 0;
    exp_54_ram[51] = 0;
    exp_54_ram[52] = 2;
    exp_54_ram[53] = 0;
    exp_54_ram[54] = 64;
    exp_54_ram[55] = 0;
    exp_54_ram[56] = 0;
    exp_54_ram[57] = 0;
    exp_54_ram[58] = 0;
    exp_54_ram[59] = 0;
    exp_54_ram[60] = 0;
    exp_54_ram[61] = 1;
    exp_54_ram[62] = 3;
    exp_54_ram[63] = 1;
    exp_54_ram[64] = 1;
    exp_54_ram[65] = 1;
    exp_54_ram[66] = 3;
    exp_54_ram[67] = 0;
    exp_54_ram[68] = 2;
    exp_54_ram[69] = 1;
    exp_54_ram[70] = 0;
    exp_54_ram[71] = 0;
    exp_54_ram[72] = 1;
    exp_54_ram[73] = 255;
    exp_54_ram[74] = 1;
    exp_54_ram[75] = 0;
    exp_54_ram[76] = 255;
    exp_54_ram[77] = 1;
    exp_54_ram[78] = 64;
    exp_54_ram[79] = 3;
    exp_54_ram[80] = 1;
    exp_54_ram[81] = 1;
    exp_54_ram[82] = 3;
    exp_54_ram[83] = 1;
    exp_54_ram[84] = 0;
    exp_54_ram[85] = 2;
    exp_54_ram[86] = 0;
    exp_54_ram[87] = 0;
    exp_54_ram[88] = 0;
    exp_54_ram[89] = 255;
    exp_54_ram[90] = 1;
    exp_54_ram[91] = 0;
    exp_54_ram[92] = 255;
    exp_54_ram[93] = 1;
    exp_54_ram[94] = 0;
    exp_54_ram[95] = 0;
    exp_54_ram[96] = 14;
    exp_54_ram[97] = 1;
    exp_54_ram[98] = 1;
    exp_54_ram[99] = 242;
    exp_54_ram[100] = 1;
    exp_54_ram[101] = 243;
    exp_54_ram[102] = 0;
    exp_54_ram[103] = 0;
    exp_54_ram[104] = 2;
    exp_54_ram[105] = 0;
    exp_54_ram[106] = 12;
    exp_54_ram[107] = 15;
    exp_54_ram[108] = 1;
    exp_54_ram[109] = 0;
    exp_54_ram[110] = 0;
    exp_54_ram[111] = 0;
    exp_54_ram[112] = 0;
    exp_54_ram[113] = 2;
    exp_54_ram[114] = 0;
    exp_54_ram[115] = 64;
    exp_54_ram[116] = 10;
    exp_54_ram[117] = 65;
    exp_54_ram[118] = 0;
    exp_54_ram[119] = 1;
    exp_54_ram[120] = 1;
    exp_54_ram[121] = 1;
    exp_54_ram[122] = 1;
    exp_54_ram[123] = 3;
    exp_54_ram[124] = 3;
    exp_54_ram[125] = 1;
    exp_54_ram[126] = 0;
    exp_54_ram[127] = 2;
    exp_54_ram[128] = 0;
    exp_54_ram[129] = 1;
    exp_54_ram[130] = 1;
    exp_54_ram[131] = 255;
    exp_54_ram[132] = 1;
    exp_54_ram[133] = 1;
    exp_54_ram[134] = 255;
    exp_54_ram[135] = 1;
    exp_54_ram[136] = 65;
    exp_54_ram[137] = 3;
    exp_54_ram[138] = 1;
    exp_54_ram[139] = 1;
    exp_54_ram[140] = 3;
    exp_54_ram[141] = 1;
    exp_54_ram[142] = 0;
    exp_54_ram[143] = 2;
    exp_54_ram[144] = 0;
    exp_54_ram[145] = 0;
    exp_54_ram[146] = 0;
    exp_54_ram[147] = 255;
    exp_54_ram[148] = 1;
    exp_54_ram[149] = 0;
    exp_54_ram[150] = 255;
    exp_54_ram[151] = 1;
    exp_54_ram[152] = 0;
    exp_54_ram[153] = 0;
    exp_54_ram[154] = 1;
    exp_54_ram[155] = 1;
    exp_54_ram[156] = 244;
    exp_54_ram[157] = 1;
    exp_54_ram[158] = 244;
    exp_54_ram[159] = 0;
    exp_54_ram[160] = 0;
    exp_54_ram[161] = 0;
    exp_54_ram[162] = 0;
    exp_54_ram[163] = 0;
    exp_54_ram[164] = 1;
    exp_54_ram[165] = 0;
    exp_54_ram[166] = 3;
    exp_54_ram[167] = 1;
    exp_54_ram[168] = 1;
    exp_54_ram[169] = 1;
    exp_54_ram[170] = 3;
    exp_54_ram[171] = 1;
    exp_54_ram[172] = 0;
    exp_54_ram[173] = 2;
    exp_54_ram[174] = 0;
    exp_54_ram[175] = 0;
    exp_54_ram[176] = 1;
    exp_54_ram[177] = 255;
    exp_54_ram[178] = 1;
    exp_54_ram[179] = 0;
    exp_54_ram[180] = 255;
    exp_54_ram[181] = 1;
    exp_54_ram[182] = 64;
    exp_54_ram[183] = 3;
    exp_54_ram[184] = 1;
    exp_54_ram[185] = 1;
    exp_54_ram[186] = 3;
    exp_54_ram[187] = 1;
    exp_54_ram[188] = 2;
    exp_54_ram[189] = 0;
    exp_54_ram[190] = 0;
    exp_54_ram[191] = 0;
    exp_54_ram[192] = 1;
    exp_54_ram[193] = 255;
    exp_54_ram[194] = 1;
    exp_54_ram[195] = 0;
    exp_54_ram[196] = 255;
    exp_54_ram[197] = 1;
    exp_54_ram[198] = 1;
    exp_54_ram[199] = 64;
    exp_54_ram[200] = 0;
    exp_54_ram[201] = 235;
    exp_54_ram[202] = 24;
    exp_54_ram[203] = 0;
    exp_54_ram[204] = 4;
    exp_54_ram[205] = 15;
    exp_54_ram[206] = 0;
    exp_54_ram[207] = 0;
    exp_54_ram[208] = 0;
    exp_54_ram[209] = 0;
    exp_54_ram[210] = 188;
    exp_54_ram[211] = 0;
    exp_54_ram[212] = 0;
    exp_54_ram[213] = 2;
    exp_54_ram[214] = 0;
    exp_54_ram[215] = 64;
    exp_54_ram[216] = 2;
    exp_54_ram[217] = 0;
    exp_54_ram[218] = 238;
    exp_54_ram[219] = 0;
    exp_54_ram[220] = 0;
    exp_54_ram[221] = 239;
    exp_54_ram[222] = 1;
    exp_54_ram[223] = 1;
    exp_54_ram[224] = 252;
    exp_54_ram[225] = 1;
    exp_54_ram[226] = 251;
    exp_54_ram[227] = 0;
    exp_54_ram[228] = 0;
    exp_54_ram[229] = 0;
    exp_54_ram[230] = 0;
    exp_54_ram[231] = 1;
    exp_54_ram[232] = 3;
    exp_54_ram[233] = 0;
    exp_54_ram[234] = 0;
    exp_54_ram[235] = 0;
    exp_54_ram[236] = 0;
    exp_54_ram[237] = 1;
    exp_54_ram[238] = 1;
    exp_54_ram[239] = 1;
    exp_54_ram[240] = 3;
    exp_54_ram[241] = 1;
    exp_54_ram[242] = 0;
    exp_54_ram[243] = 3;
    exp_54_ram[244] = 0;
    exp_54_ram[245] = 1;
    exp_54_ram[246] = 1;
    exp_54_ram[247] = 255;
    exp_54_ram[248] = 1;
    exp_54_ram[249] = 1;
    exp_54_ram[250] = 255;
    exp_54_ram[251] = 1;
    exp_54_ram[252] = 65;
    exp_54_ram[253] = 3;
    exp_54_ram[254] = 3;
    exp_54_ram[255] = 1;
    exp_54_ram[256] = 2;
    exp_54_ram[257] = 1;
    exp_54_ram[258] = 1;
    exp_54_ram[259] = 0;
    exp_54_ram[260] = 0;
    exp_54_ram[261] = 1;
    exp_54_ram[262] = 1;
    exp_54_ram[263] = 255;
    exp_54_ram[264] = 1;
    exp_54_ram[265] = 1;
    exp_54_ram[266] = 255;
    exp_54_ram[267] = 1;
    exp_54_ram[268] = 1;
    exp_54_ram[269] = 0;
    exp_54_ram[270] = 0;
    exp_54_ram[271] = 255;
    exp_54_ram[272] = 0;
    exp_54_ram[273] = 1;
    exp_54_ram[274] = 0;
    exp_54_ram[275] = 1;
    exp_54_ram[276] = 65;
    exp_54_ram[277] = 2;
    exp_54_ram[278] = 2;
    exp_54_ram[279] = 1;
    exp_54_ram[280] = 2;
    exp_54_ram[281] = 0;
    exp_54_ram[282] = 1;
    exp_54_ram[283] = 2;
    exp_54_ram[284] = 0;
    exp_54_ram[285] = 1;
    exp_54_ram[286] = 1;
    exp_54_ram[287] = 0;
    exp_54_ram[288] = 2;
    exp_54_ram[289] = 206;
    exp_54_ram[290] = 0;
    exp_54_ram[291] = 255;
    exp_54_ram[292] = 0;
    exp_54_ram[293] = 1;
    exp_54_ram[294] = 0;
    exp_54_ram[295] = 0;
    exp_54_ram[296] = 1;
    exp_54_ram[297] = 0;
    exp_54_ram[298] = 218;
    exp_54_ram[299] = 255;
    exp_54_ram[300] = 204;
    exp_54_ram[301] = 0;
    exp_54_ram[302] = 0;
    exp_54_ram[303] = 218;
    exp_54_ram[304] = 0;
    exp_54_ram[305] = 255;
    exp_54_ram[306] = 1;
    exp_54_ram[307] = 0;
    exp_54_ram[308] = 0;
    exp_54_ram[309] = 0;
    exp_54_ram[310] = 127;
    exp_54_ram[311] = 1;
    exp_54_ram[312] = 127;
    exp_54_ram[313] = 1;
    exp_54_ram[314] = 0;
    exp_54_ram[315] = 0;
    exp_54_ram[316] = 127;
    exp_54_ram[317] = 1;
    exp_54_ram[318] = 1;
    exp_54_ram[319] = 0;
    exp_54_ram[320] = 8;
    exp_54_ram[321] = 0;
    exp_54_ram[322] = 0;
    exp_54_ram[323] = 1;
    exp_54_ram[324] = 0;
    exp_54_ram[325] = 254;
    exp_54_ram[326] = 8;
    exp_54_ram[327] = 0;
    exp_54_ram[328] = 0;
    exp_54_ram[329] = 0;
    exp_54_ram[330] = 0;
    exp_54_ram[331] = 4;
    exp_54_ram[332] = 0;
    exp_54_ram[333] = 0;
    exp_54_ram[334] = 3;
    exp_54_ram[335] = 4;
    exp_54_ram[336] = 255;
    exp_54_ram[337] = 0;
    exp_54_ram[338] = 255;
    exp_54_ram[339] = 0;
    exp_54_ram[340] = 0;
    exp_54_ram[341] = 0;
    exp_54_ram[342] = 0;
    exp_54_ram[343] = 254;
    exp_54_ram[344] = 0;
    exp_54_ram[345] = 253;
    exp_54_ram[346] = 2;
    exp_54_ram[347] = 252;
    exp_54_ram[348] = 255;
    exp_54_ram[349] = 0;
    exp_54_ram[350] = 0;
    exp_54_ram[351] = 0;
    exp_54_ram[352] = 0;
    exp_54_ram[353] = 254;
    exp_54_ram[354] = 251;
    exp_54_ram[355] = 252;
    exp_54_ram[356] = 254;
    exp_54_ram[357] = 247;
    exp_54_ram[358] = 248;
    exp_54_ram[359] = 0;
    exp_54_ram[360] = 248;
    exp_54_ram[361] = 255;
    exp_54_ram[362] = 0;
    exp_54_ram[363] = 0;
    exp_54_ram[364] = 0;
    exp_54_ram[365] = 6;
    exp_54_ram[366] = 55;
    exp_54_ram[367] = 65;
    exp_54_ram[368] = 0;
    exp_54_ram[369] = 64;
    exp_54_ram[370] = 4;
    exp_54_ram[371] = 0;
    exp_54_ram[372] = 64;
    exp_54_ram[373] = 1;
    exp_54_ram[374] = 0;
    exp_54_ram[375] = 0;
    exp_54_ram[376] = 0;
    exp_54_ram[377] = 0;
    exp_54_ram[378] = 0;
    exp_54_ram[379] = 0;
    exp_54_ram[380] = 1;
    exp_54_ram[381] = 0;
    exp_54_ram[382] = 0;
    exp_54_ram[383] = 0;
    exp_54_ram[384] = 1;
    exp_54_ram[385] = 0;
    exp_54_ram[386] = 255;
    exp_54_ram[387] = 0;
    exp_54_ram[388] = 0;
    exp_54_ram[389] = 252;
    exp_54_ram[390] = 0;
    exp_54_ram[391] = 0;
    exp_54_ram[392] = 252;
    exp_54_ram[393] = 254;
    exp_54_ram[394] = 0;
    exp_54_ram[395] = 0;
    exp_54_ram[396] = 0;
    exp_54_ram[397] = 1;
    exp_54_ram[398] = 1;
    exp_54_ram[399] = 1;
    exp_54_ram[400] = 0;
    exp_54_ram[401] = 24;
    exp_54_ram[402] = 0;
    exp_54_ram[403] = 0;
    exp_54_ram[404] = 0;
    exp_54_ram[405] = 8;
    exp_54_ram[406] = 0;
    exp_54_ram[407] = 45;
    exp_54_ram[408] = 0;
    exp_54_ram[409] = 67;
    exp_54_ram[410] = 65;
    exp_54_ram[411] = 67;
    exp_54_ram[412] = 9;
    exp_54_ram[413] = 0;
    exp_54_ram[414] = 0;
    exp_54_ram[415] = 3;
    exp_54_ram[416] = 2;
    exp_54_ram[417] = 7;
    exp_54_ram[418] = 2;
    exp_54_ram[419] = 255;
    exp_54_ram[420] = 65;
    exp_54_ram[421] = 0;
    exp_54_ram[422] = 0;
    exp_54_ram[423] = 0;
    exp_54_ram[424] = 0;
    exp_54_ram[425] = 1;
    exp_54_ram[426] = 1;
    exp_54_ram[427] = 0;
    exp_54_ram[428] = 1;
    exp_54_ram[429] = 0;
    exp_54_ram[430] = 0;
    exp_54_ram[431] = 1;
    exp_54_ram[432] = 1;
    exp_54_ram[433] = 0;
    exp_54_ram[434] = 0;
    exp_54_ram[435] = 0;
    exp_54_ram[436] = 0;
    exp_54_ram[437] = 2;
    exp_54_ram[438] = 0;
    exp_54_ram[439] = 37;
    exp_54_ram[440] = 2;
    exp_54_ram[441] = 248;
    exp_54_ram[442] = 253;
    exp_54_ram[443] = 0;
    exp_54_ram[444] = 0;
    exp_54_ram[445] = 251;
    exp_54_ram[446] = 67;
    exp_54_ram[447] = 3;
    exp_54_ram[448] = 3;
    exp_54_ram[449] = 0;
    exp_54_ram[450] = 0;
    exp_54_ram[451] = 31;
    exp_54_ram[452] = 0;
    exp_54_ram[453] = 0;
    exp_54_ram[454] = 0;
    exp_54_ram[455] = 0;
    exp_54_ram[456] = 0;
    exp_54_ram[457] = 65;
    exp_54_ram[458] = 25;
    exp_54_ram[459] = 0;
    exp_54_ram[460] = 0;
    exp_54_ram[461] = 0;
    exp_54_ram[462] = 0;
    exp_54_ram[463] = 0;
    exp_54_ram[464] = 3;
    exp_54_ram[465] = 2;
    exp_54_ram[466] = 9;
    exp_54_ram[467] = 255;
    exp_54_ram[468] = 0;
    exp_54_ram[469] = 2;
    exp_54_ram[470] = 65;
    exp_54_ram[471] = 1;
    exp_54_ram[472] = 0;
    exp_54_ram[473] = 0;
    exp_54_ram[474] = 255;
    exp_54_ram[475] = 255;
    exp_54_ram[476] = 0;
    exp_54_ram[477] = 0;
    exp_54_ram[478] = 2;
    exp_54_ram[479] = 0;
    exp_54_ram[480] = 0;
    exp_54_ram[481] = 0;
    exp_54_ram[482] = 0;
    exp_54_ram[483] = 0;
    exp_54_ram[484] = 0;
    exp_54_ram[485] = 0;
    exp_54_ram[486] = 0;
    exp_54_ram[487] = 0;
    exp_54_ram[488] = 0;
    exp_54_ram[489] = 255;
    exp_54_ram[490] = 255;
    exp_54_ram[491] = 67;
    exp_54_ram[492] = 0;
    exp_54_ram[493] = 65;
    exp_54_ram[494] = 0;
    exp_54_ram[495] = 1;
    exp_54_ram[496] = 0;
    exp_54_ram[497] = 0;
    exp_54_ram[498] = 237;
    exp_54_ram[499] = 253;
    exp_54_ram[500] = 0;
    exp_54_ram[501] = 0;
    exp_54_ram[502] = 249;
    exp_54_ram[503] = 0;
    exp_54_ram[504] = 0;
    exp_54_ram[505] = 0;
    exp_54_ram[506] = 235;
    exp_54_ram[507] = 0;
    exp_54_ram[508] = 0;
    exp_54_ram[509] = 0;
    exp_54_ram[510] = 0;
    exp_54_ram[511] = 0;
    exp_54_ram[512] = 0;
    exp_54_ram[513] = 0;
    exp_54_ram[514] = 254;
    exp_54_ram[515] = 0;
    exp_54_ram[516] = 6;
    exp_54_ram[517] = 6;
    exp_54_ram[518] = 0;
    exp_54_ram[519] = 0;
    exp_54_ram[520] = 255;
    exp_54_ram[521] = 2;
    exp_54_ram[522] = 0;
    exp_54_ram[523] = 0;
    exp_54_ram[524] = 0;
    exp_54_ram[525] = 0;
    exp_54_ram[526] = 0;
    exp_54_ram[527] = 254;
    exp_54_ram[528] = 0;
    exp_54_ram[529] = 0;
    exp_54_ram[530] = 64;
    exp_54_ram[531] = 0;
    exp_54_ram[532] = 0;
    exp_54_ram[533] = 0;
    exp_54_ram[534] = 254;
    exp_54_ram[535] = 0;
    exp_54_ram[536] = 0;
    exp_54_ram[537] = 251;
    exp_54_ram[538] = 0;
    exp_54_ram[539] = 0;
    exp_54_ram[540] = 64;
    exp_54_ram[541] = 0;
    exp_54_ram[542] = 64;
    exp_54_ram[543] = 249;
    exp_54_ram[544] = 64;
    exp_54_ram[545] = 0;
    exp_54_ram[546] = 249;
    exp_54_ram[547] = 64;
    exp_54_ram[548] = 0;
    exp_54_ram[549] = 0;
    exp_54_ram[550] = 0;
    exp_54_ram[551] = 0;
    exp_54_ram[552] = 247;
    exp_54_ram[553] = 0;
    exp_54_ram[554] = 0;
    exp_54_ram[555] = 64;
    exp_54_ram[556] = 254;
    exp_54_ram[557] = 64;
    exp_54_ram[558] = 246;
    exp_54_ram[559] = 64;
    exp_54_ram[560] = 0;
    exp_54_ram[561] = 2;
    exp_54_ram[562] = 2;
    exp_54_ram[563] = 64;
    exp_54_ram[564] = 0;
    exp_54_ram[565] = 254;
    exp_54_ram[566] = 0;
    exp_54_ram[567] = 0;
    exp_54_ram[568] = 0;
    exp_54_ram[569] = 0;
    exp_54_ram[570] = 0;
    exp_54_ram[571] = 0;
    exp_54_ram[572] = 0;
    exp_54_ram[573] = 0;
    exp_54_ram[574] = 254;
    exp_54_ram[575] = 2;
    exp_54_ram[576] = 2;
    exp_54_ram[577] = 64;
    exp_54_ram[578] = 0;
    exp_54_ram[579] = 254;
    exp_54_ram[580] = 0;
    exp_54_ram[581] = 0;
    exp_54_ram[582] = 0;
    exp_54_ram[583] = 0;
    exp_54_ram[584] = 0;
    exp_54_ram[585] = 0;
    exp_54_ram[586] = 0;
    exp_54_ram[587] = 0;
    exp_54_ram[588] = 254;
    exp_54_ram[589] = 0;
    exp_54_ram[590] = 2;
    exp_54_ram[591] = 15;
    exp_54_ram[592] = 0;
    exp_54_ram[593] = 0;
    exp_54_ram[594] = 0;
    exp_54_ram[595] = 2;
    exp_54_ram[596] = 64;
    exp_54_ram[597] = 0;
    exp_54_ram[598] = 188;
    exp_54_ram[599] = 0;
    exp_54_ram[600] = 0;
    exp_54_ram[601] = 64;
    exp_54_ram[602] = 0;
    exp_54_ram[603] = 1;
    exp_54_ram[604] = 1;
    exp_54_ram[605] = 252;
    exp_54_ram[606] = 1;
    exp_54_ram[607] = 252;
    exp_54_ram[608] = 99;
    exp_54_ram[609] = 46;
    exp_54_ram[610] = 0;
    exp_54_ram[611] = 0;
    exp_54_ram[612] = 108;
    exp_54_ram[613] = 0;
    exp_54_ram[614] = 97;
    exp_54_ram[615] = 0;
    exp_54_ram[616] = 97;
    exp_54_ram[617] = 0;
    exp_54_ram[618] = 0;
    exp_54_ram[619] = 97;
    exp_54_ram[620] = 0;
    exp_54_ram[621] = 97;
    exp_54_ram[622] = 0;
    exp_54_ram[623] = 115;
    exp_54_ram[624] = 0;
    exp_54_ram[625] = 110;
    exp_54_ram[626] = 46;
    exp_54_ram[627] = 0;
    exp_54_ram[628] = 120;
    exp_54_ram[629] = 0;
    exp_54_ram[630] = 99;
    exp_54_ram[631] = 46;
    exp_54_ram[632] = 0;
    exp_54_ram[633] = 99;
    exp_54_ram[634] = 46;
    exp_54_ram[635] = 0;
    exp_54_ram[636] = 110;
    exp_54_ram[637] = 46;
    exp_54_ram[638] = 0;
    exp_54_ram[639] = 99;
    exp_54_ram[640] = 46;
    exp_54_ram[641] = 0;
    exp_54_ram[642] = 97;
    exp_54_ram[643] = 0;
    exp_54_ram[644] = 99;
    exp_54_ram[645] = 46;
    exp_54_ram[646] = 0;
    exp_54_ram[647] = 97;
    exp_54_ram[648] = 0;
    exp_54_ram[649] = 99;
    exp_54_ram[650] = 46;
    exp_54_ram[651] = 0;
    exp_54_ram[652] = 102;
    exp_54_ram[653] = 0;
    exp_54_ram[654] = 102;
    exp_54_ram[655] = 102;
    exp_54_ram[656] = 0;
    exp_54_ram[657] = 102;
    exp_54_ram[658] = 102;
    exp_54_ram[659] = 0;
    exp_54_ram[660] = 97;
    exp_54_ram[661] = 52;
    exp_54_ram[662] = 0;
    exp_54_ram[663] = 102;
    exp_54_ram[664] = 102;
    exp_54_ram[665] = 0;
    exp_54_ram[666] = 112;
    exp_54_ram[667] = 46;
    exp_54_ram[668] = 0;
    exp_54_ram[669] = 102;
    exp_54_ram[670] = 49;
    exp_54_ram[671] = 0;
    exp_54_ram[672] = 50;
    exp_54_ram[673] = 0;
    exp_54_ram[674] = 51;
    exp_54_ram[675] = 0;
    exp_54_ram[676] = 100;
    exp_54_ram[677] = 0;
    exp_54_ram[678] = 102;
    exp_54_ram[679] = 102;
    exp_54_ram[680] = 0;
    exp_54_ram[681] = 114;
    exp_54_ram[682] = 46;
    exp_54_ram[683] = 0;
    exp_54_ram[684] = 115;
    exp_54_ram[685] = 46;
    exp_54_ram[686] = 0;
    exp_54_ram[687] = 100;
    exp_54_ram[688] = 0;
    exp_54_ram[689] = 100;
    exp_54_ram[690] = 115;
    exp_54_ram[691] = 0;
    exp_54_ram[692] = 102;
    exp_54_ram[693] = 50;
    exp_54_ram[694] = 0;
    exp_54_ram[695] = 100;
    exp_54_ram[696] = 52;
    exp_54_ram[697] = 102;
    exp_54_ram[698] = 0;
    exp_54_ram[699] = 115;
    exp_54_ram[700] = 46;
    exp_54_ram[701] = 0;
    exp_54_ram[702] = 52;
    exp_54_ram[703] = 0;
    exp_54_ram[704] = 0;
    exp_54_ram[705] = 0;
    exp_54_ram[706] = 115;
    exp_54_ram[707] = 46;
    exp_54_ram[708] = 0;
    exp_54_ram[709] = 52;
    exp_54_ram[710] = 0;
    exp_54_ram[711] = 52;
    exp_54_ram[712] = 0;
    exp_54_ram[713] = 52;
    exp_54_ram[714] = 0;
    exp_54_ram[715] = 100;
    exp_54_ram[716] = 0;
    exp_54_ram[717] = 108;
    exp_54_ram[718] = 46;
    exp_54_ram[719] = 0;
    exp_54_ram[720] = 101;
    exp_54_ram[721] = 0;
    exp_54_ram[722] = 32;
    exp_54_ram[723] = 32;
    exp_54_ram[724] = 48;
    exp_54_ram[725] = 49;
    exp_54_ram[726] = 32;
    exp_54_ram[727] = 48;
    exp_54_ram[728] = 0;
    exp_54_ram[729] = 32;
    exp_54_ram[730] = 32;
    exp_54_ram[731] = 48;
    exp_54_ram[732] = 49;
    exp_54_ram[733] = 32;
    exp_54_ram[734] = 48;
    exp_54_ram[735] = 0;
    exp_54_ram[736] = 97;
    exp_54_ram[737] = 0;
    exp_54_ram[738] = 97;
    exp_54_ram[739] = 0;
    exp_54_ram[740] = 97;
    exp_54_ram[741] = 0;
    exp_54_ram[742] = 32;
    exp_54_ram[743] = 32;
    exp_54_ram[744] = 48;
    exp_54_ram[745] = 49;
    exp_54_ram[746] = 32;
    exp_54_ram[747] = 48;
    exp_54_ram[748] = 0;
    exp_54_ram[749] = 102;
    exp_54_ram[750] = 0;
    exp_54_ram[751] = 102;
    exp_54_ram[752] = 0;
    exp_54_ram[753] = 102;
    exp_54_ram[754] = 0;
    exp_54_ram[755] = 2;
    exp_54_ram[756] = 3;
    exp_54_ram[757] = 4;
    exp_54_ram[758] = 4;
    exp_54_ram[759] = 5;
    exp_54_ram[760] = 5;
    exp_54_ram[761] = 5;
    exp_54_ram[762] = 5;
    exp_54_ram[763] = 6;
    exp_54_ram[764] = 6;
    exp_54_ram[765] = 6;
    exp_54_ram[766] = 6;
    exp_54_ram[767] = 6;
    exp_54_ram[768] = 6;
    exp_54_ram[769] = 6;
    exp_54_ram[770] = 6;
    exp_54_ram[771] = 7;
    exp_54_ram[772] = 7;
    exp_54_ram[773] = 7;
    exp_54_ram[774] = 7;
    exp_54_ram[775] = 7;
    exp_54_ram[776] = 7;
    exp_54_ram[777] = 7;
    exp_54_ram[778] = 7;
    exp_54_ram[779] = 7;
    exp_54_ram[780] = 7;
    exp_54_ram[781] = 7;
    exp_54_ram[782] = 7;
    exp_54_ram[783] = 7;
    exp_54_ram[784] = 7;
    exp_54_ram[785] = 7;
    exp_54_ram[786] = 7;
    exp_54_ram[787] = 8;
    exp_54_ram[788] = 8;
    exp_54_ram[789] = 8;
    exp_54_ram[790] = 8;
    exp_54_ram[791] = 8;
    exp_54_ram[792] = 8;
    exp_54_ram[793] = 8;
    exp_54_ram[794] = 8;
    exp_54_ram[795] = 8;
    exp_54_ram[796] = 8;
    exp_54_ram[797] = 8;
    exp_54_ram[798] = 8;
    exp_54_ram[799] = 8;
    exp_54_ram[800] = 8;
    exp_54_ram[801] = 8;
    exp_54_ram[802] = 8;
    exp_54_ram[803] = 8;
    exp_54_ram[804] = 8;
    exp_54_ram[805] = 8;
    exp_54_ram[806] = 8;
    exp_54_ram[807] = 8;
    exp_54_ram[808] = 8;
    exp_54_ram[809] = 8;
    exp_54_ram[810] = 8;
    exp_54_ram[811] = 8;
    exp_54_ram[812] = 8;
    exp_54_ram[813] = 8;
    exp_54_ram[814] = 8;
    exp_54_ram[815] = 8;
    exp_54_ram[816] = 8;
    exp_54_ram[817] = 8;
    exp_54_ram[818] = 8;
    exp_54_ram[819] = 0;
    exp_54_ram[820] = 0;
    exp_54_ram[821] = 0;
    exp_54_ram[822] = 0;
    exp_54_ram[823] = 0;
    exp_54_ram[824] = 0;
    exp_54_ram[825] = 0;
    exp_54_ram[826] = 0;
    exp_54_ram[827] = 254;
    exp_54_ram[828] = 255;
    exp_54_ram[829] = 0;
    exp_54_ram[830] = 0;
    exp_54_ram[831] = 12;
    exp_54_ram[832] = 0;
    exp_54_ram[833] = 0;
    exp_54_ram[834] = 252;
    exp_54_ram[835] = 0;
    exp_54_ram[836] = 0;
    exp_54_ram[837] = 0;
    exp_54_ram[838] = 0;
    exp_54_ram[839] = 0;
    exp_54_ram[840] = 1;
    exp_54_ram[841] = 0;
    exp_54_ram[842] = 0;
    exp_54_ram[843] = 0;
    exp_54_ram[844] = 0;
    exp_54_ram[845] = 6;
    exp_54_ram[846] = 0;
    exp_54_ram[847] = 0;
    exp_54_ram[848] = 0;
    exp_54_ram[849] = 2;
    exp_54_ram[850] = 0;
    exp_54_ram[851] = 1;
    exp_54_ram[852] = 1;
    exp_54_ram[853] = 255;
    exp_54_ram[854] = 255;
    exp_54_ram[855] = 255;
    exp_54_ram[856] = 255;
    exp_54_ram[857] = 255;
    exp_54_ram[858] = 255;
    exp_54_ram[859] = 255;
    exp_54_ram[860] = 64;
    exp_54_ram[861] = 253;
    exp_54_ram[862] = 0;
    exp_54_ram[863] = 255;
    exp_54_ram[864] = 0;
    exp_54_ram[865] = 0;
    exp_54_ram[866] = 0;
    exp_54_ram[867] = 64;
    exp_54_ram[868] = 3;
    exp_54_ram[869] = 0;
    exp_54_ram[870] = 0;
    exp_54_ram[871] = 0;
    exp_54_ram[872] = 0;
    exp_54_ram[873] = 0;
    exp_54_ram[874] = 2;
    exp_54_ram[875] = 0;
    exp_54_ram[876] = 0;
    exp_54_ram[877] = 0;
    exp_54_ram[878] = 0;
    exp_54_ram[879] = 0;
    exp_54_ram[880] = 1;
    exp_54_ram[881] = 252;
    exp_54_ram[882] = 0;
    exp_54_ram[883] = 0;
    exp_54_ram[884] = 0;
    exp_54_ram[885] = 0;
    exp_54_ram[886] = 1;
    exp_54_ram[887] = 252;
    exp_54_ram[888] = 0;
    exp_54_ram[889] = 0;
    exp_54_ram[890] = 0;
    exp_54_ram[891] = 0;
    exp_54_ram[892] = 0;
    exp_54_ram[893] = 0;
    exp_54_ram[894] = 255;
    exp_54_ram[895] = 2;
    exp_54_ram[896] = 0;
    exp_54_ram[897] = 0;
    exp_54_ram[898] = 253;
    exp_54_ram[899] = 254;
    exp_54_ram[900] = 0;
    exp_54_ram[901] = 0;
    exp_54_ram[902] = 254;
    exp_54_ram[903] = 253;
    exp_54_ram[904] = 0;
    exp_54_ram[905] = 0;
    exp_54_ram[906] = 0;
    exp_54_ram[907] = 0;
    exp_54_ram[908] = 2;
    exp_54_ram[909] = 254;
    exp_54_ram[910] = 128;
    exp_54_ram[911] = 239;
    exp_54_ram[912] = 8;
    exp_54_ram[913] = 0;
    exp_54_ram[914] = 0;
    exp_54_ram[915] = 0;
    exp_54_ram[916] = 0;
    exp_54_ram[917] = 0;
    exp_54_ram[918] = 0;
    exp_54_ram[919] = 2;
    exp_54_ram[920] = 64;
    exp_54_ram[921] = 0;
    exp_54_ram[922] = 0;
    exp_54_ram[923] = 255;
    exp_54_ram[924] = 0;
    exp_54_ram[925] = 0;
    exp_54_ram[926] = 0;
    exp_54_ram[927] = 0;
    exp_54_ram[928] = 0;
    exp_54_ram[929] = 252;
    exp_54_ram[930] = 0;
    exp_54_ram[931] = 0;
    exp_54_ram[932] = 252;
    exp_54_ram[933] = 0;
    exp_54_ram[934] = 0;
    exp_54_ram[935] = 0;
    exp_54_ram[936] = 0;
    exp_54_ram[937] = 0;
    exp_54_ram[938] = 0;
    exp_54_ram[939] = 0;
    exp_54_ram[940] = 0;
    exp_54_ram[941] = 0;
    exp_54_ram[942] = 254;
    exp_54_ram[943] = 0;
    exp_54_ram[944] = 0;
    exp_54_ram[945] = 0;
    exp_54_ram[946] = 0;
    exp_54_ram[947] = 0;
    exp_54_ram[948] = 0;
    exp_54_ram[949] = 254;
    exp_54_ram[950] = 0;
    exp_54_ram[951] = 0;
    exp_54_ram[952] = 0;
    exp_54_ram[953] = 0;
    exp_54_ram[954] = 1;
    exp_54_ram[955] = 0;
    exp_54_ram[956] = 0;
    exp_54_ram[957] = 0;
    exp_54_ram[958] = 254;
    exp_54_ram[959] = 0;
    exp_54_ram[960] = 255;
    exp_54_ram[961] = 0;
    exp_54_ram[962] = 0;
    exp_54_ram[963] = 0;
    exp_54_ram[964] = 0;
    exp_54_ram[965] = 0;
    exp_54_ram[966] = 248;
    exp_54_ram[967] = 0;
    exp_54_ram[968] = 0;
    exp_54_ram[969] = 0;
    exp_54_ram[970] = 0;
    exp_54_ram[971] = 1;
    exp_54_ram[972] = 0;
    exp_54_ram[973] = 0;
    exp_54_ram[974] = 0;
    exp_54_ram[975] = 254;
    exp_54_ram[976] = 0;
    exp_54_ram[977] = 0;
    exp_54_ram[978] = 0;
    exp_54_ram[979] = 1;
    exp_54_ram[980] = 0;
    exp_54_ram[981] = 255;
    exp_54_ram[982] = 0;
    exp_54_ram[983] = 0;
    exp_54_ram[984] = 0;
    exp_54_ram[985] = 0;
    exp_54_ram[986] = 0;
    exp_54_ram[987] = 243;
    exp_54_ram[988] = 255;
    exp_54_ram[989] = 0;
    exp_54_ram[990] = 0;
    exp_54_ram[991] = 0;
    exp_54_ram[992] = 1;
    exp_54_ram[993] = 0;
    exp_54_ram[994] = 0;
    exp_54_ram[995] = 255;
    exp_54_ram[996] = 254;
    exp_54_ram[997] = 0;
    exp_54_ram[998] = 0;
    exp_54_ram[999] = 0;
    exp_54_ram[1000] = 1;
    exp_54_ram[1001] = 0;
    exp_54_ram[1002] = 254;
    exp_54_ram[1003] = 0;
    exp_54_ram[1004] = 0;
    exp_54_ram[1005] = 1;
    exp_54_ram[1006] = 1;
    exp_54_ram[1007] = 0;
    exp_54_ram[1008] = 0;
    exp_54_ram[1009] = 0;
    exp_54_ram[1010] = 237;
    exp_54_ram[1011] = 0;
    exp_54_ram[1012] = 0;
    exp_54_ram[1013] = 2;
    exp_54_ram[1014] = 0;
    exp_54_ram[1015] = 236;
    exp_54_ram[1016] = 0;
    exp_54_ram[1017] = 0;
    exp_54_ram[1018] = 1;
    exp_54_ram[1019] = 0;
    exp_54_ram[1020] = 0;
    exp_54_ram[1021] = 0;
    exp_54_ram[1022] = 2;
    exp_54_ram[1023] = 0;
    exp_54_ram[1024] = 254;
    exp_54_ram[1025] = 1;
    exp_54_ram[1026] = 0;
    exp_54_ram[1027] = 1;
    exp_54_ram[1028] = 1;
    exp_54_ram[1029] = 1;
    exp_54_ram[1030] = 0;
    exp_54_ram[1031] = 2;
    exp_54_ram[1032] = 0;
    exp_54_ram[1033] = 0;
    exp_54_ram[1034] = 250;
    exp_54_ram[1035] = 254;
    exp_54_ram[1036] = 0;
    exp_54_ram[1037] = 0;
    exp_54_ram[1038] = 1;
    exp_54_ram[1039] = 1;
    exp_54_ram[1040] = 0;
    exp_54_ram[1041] = 0;
    exp_54_ram[1042] = 0;
    exp_54_ram[1043] = 229;
    exp_54_ram[1044] = 0;
    exp_54_ram[1045] = 0;
    exp_54_ram[1046] = 2;
    exp_54_ram[1047] = 0;
    exp_54_ram[1048] = 227;
    exp_54_ram[1049] = 0;
    exp_54_ram[1050] = 0;
    exp_54_ram[1051] = 1;
    exp_54_ram[1052] = 0;
    exp_54_ram[1053] = 0;
    exp_54_ram[1054] = 0;
    exp_54_ram[1055] = 0;
    exp_54_ram[1056] = 0;
    exp_54_ram[1057] = 254;
    exp_54_ram[1058] = 0;
    exp_54_ram[1059] = 252;
    exp_54_ram[1060] = 1;
    exp_54_ram[1061] = 0;
    exp_54_ram[1062] = 1;
    exp_54_ram[1063] = 1;
    exp_54_ram[1064] = 1;
    exp_54_ram[1065] = 0;
    exp_54_ram[1066] = 2;
    exp_54_ram[1067] = 0;
    exp_54_ram[1068] = 255;
    exp_54_ram[1069] = 0;
    exp_54_ram[1070] = 0;
    exp_54_ram[1071] = 1;
    exp_54_ram[1072] = 0;
    exp_54_ram[1073] = 0;
    exp_54_ram[1074] = 0;
    exp_54_ram[1075] = 221;
    exp_54_ram[1076] = 0;
    exp_54_ram[1077] = 3;
    exp_54_ram[1078] = 0;
    exp_54_ram[1079] = 220;
    exp_54_ram[1080] = 0;
    exp_54_ram[1081] = 0;
    exp_54_ram[1082] = 1;
    exp_54_ram[1083] = 0;
    exp_54_ram[1084] = 0;
    exp_54_ram[1085] = 0;
    exp_54_ram[1086] = 0;
    exp_54_ram[1087] = 0;
    exp_54_ram[1088] = 0;
    exp_54_ram[1089] = 254;
    exp_54_ram[1090] = 0;
    exp_54_ram[1091] = 252;
    exp_54_ram[1092] = 0;
    exp_54_ram[1093] = 0;
    exp_54_ram[1094] = 0;
    exp_54_ram[1095] = 0;
    exp_54_ram[1096] = 0;
    exp_54_ram[1097] = 1;
    exp_54_ram[1098] = 0;
    exp_54_ram[1099] = 254;
    exp_54_ram[1100] = 0;
    exp_54_ram[1101] = 0;
    exp_54_ram[1102] = 1;
    exp_54_ram[1103] = 1;
    exp_54_ram[1104] = 0;
    exp_54_ram[1105] = 0;
    exp_54_ram[1106] = 0;
    exp_54_ram[1107] = 213;
    exp_54_ram[1108] = 0;
    exp_54_ram[1109] = 0;
    exp_54_ram[1110] = 4;
    exp_54_ram[1111] = 0;
    exp_54_ram[1112] = 211;
    exp_54_ram[1113] = 0;
    exp_54_ram[1114] = 0;
    exp_54_ram[1115] = 0;
    exp_54_ram[1116] = 1;
    exp_54_ram[1117] = 0;
    exp_54_ram[1118] = 0;
    exp_54_ram[1119] = 0;
    exp_54_ram[1120] = 0;
    exp_54_ram[1121] = 2;
    exp_54_ram[1122] = 0;
    exp_54_ram[1123] = 254;
    exp_54_ram[1124] = 1;
    exp_54_ram[1125] = 1;
    exp_54_ram[1126] = 1;
    exp_54_ram[1127] = 1;
    exp_54_ram[1128] = 0;
    exp_54_ram[1129] = 2;
    exp_54_ram[1130] = 0;
    exp_54_ram[1131] = 0;
    exp_54_ram[1132] = 254;
    exp_54_ram[1133] = 0;
    exp_54_ram[1134] = 250;
    exp_54_ram[1135] = 0;
    exp_54_ram[1136] = 4;
    exp_54_ram[1137] = 255;
    exp_54_ram[1138] = 6;
    exp_54_ram[1139] = 0;
    exp_54_ram[1140] = 0;
    exp_54_ram[1141] = 0;
    exp_54_ram[1142] = 232;
    exp_54_ram[1143] = 0;
    exp_54_ram[1144] = 0;
    exp_54_ram[1145] = 25;
    exp_54_ram[1146] = 0;
    exp_54_ram[1147] = 231;
    exp_54_ram[1148] = 0;
    exp_54_ram[1149] = 0;
    exp_54_ram[1150] = 0;
    exp_54_ram[1151] = 0;
    exp_54_ram[1152] = 1;
    exp_54_ram[1153] = 0;
    exp_54_ram[1154] = 0;
    exp_54_ram[1155] = 0;
    exp_54_ram[1156] = 0;
    exp_54_ram[1157] = 255;
    exp_54_ram[1158] = 255;
    exp_54_ram[1159] = 4;
    exp_54_ram[1160] = 255;
    exp_54_ram[1161] = 0;
    exp_54_ram[1162] = 1;
    exp_54_ram[1163] = 2;
    exp_54_ram[1164] = 0;
    exp_54_ram[1165] = 1;
    exp_54_ram[1166] = 2;
    exp_54_ram[1167] = 255;
    exp_54_ram[1168] = 0;
    exp_54_ram[1169] = 247;
    exp_54_ram[1170] = 0;
    exp_54_ram[1171] = 0;
    exp_54_ram[1172] = 1;
    exp_54_ram[1173] = 0;
    exp_54_ram[1174] = 1;
    exp_54_ram[1175] = 0;
    exp_54_ram[1176] = 1;
    exp_54_ram[1177] = 0;
    exp_54_ram[1178] = 0;
    exp_54_ram[1179] = 128;
    exp_54_ram[1180] = 0;
    exp_54_ram[1181] = 0;
    exp_54_ram[1182] = 0;
    exp_54_ram[1183] = 0;
    exp_54_ram[1184] = 0;
    exp_54_ram[1185] = 0;
    exp_54_ram[1186] = 0;
    exp_54_ram[1187] = 0;
    exp_54_ram[1188] = 64;
    exp_54_ram[1189] = 0;
    exp_54_ram[1190] = 64;
    exp_54_ram[1191] = 255;
    exp_54_ram[1192] = 64;
    exp_54_ram[1193] = 0;
    exp_54_ram[1194] = 183;
    exp_54_ram[1195] = 0;
    exp_54_ram[1196] = 1;
    exp_54_ram[1197] = 0;
    exp_54_ram[1198] = 254;
    exp_54_ram[1199] = 1;
    exp_54_ram[1200] = 1;
    exp_54_ram[1201] = 0;
    exp_54_ram[1202] = 0;
    exp_54_ram[1203] = 0;
    exp_54_ram[1204] = 1;
    exp_54_ram[1205] = 1;
    exp_54_ram[1206] = 1;
    exp_54_ram[1207] = 0;
    exp_54_ram[1208] = 1;
    exp_54_ram[1209] = 0;
    exp_54_ram[1210] = 123;
    exp_54_ram[1211] = 0;
    exp_54_ram[1212] = 0;
    exp_54_ram[1213] = 118;
    exp_54_ram[1214] = 24;
    exp_54_ram[1215] = 4;
    exp_54_ram[1216] = 1;
    exp_54_ram[1217] = 0;
    exp_54_ram[1218] = 0;
    exp_54_ram[1219] = 24;
    exp_54_ram[1220] = 6;
    exp_54_ram[1221] = 0;
    exp_54_ram[1222] = 0;
    exp_54_ram[1223] = 239;
    exp_54_ram[1224] = 0;
    exp_54_ram[1225] = 204;
    exp_54_ram[1226] = 0;
    exp_54_ram[1227] = 1;
    exp_54_ram[1228] = 1;
    exp_54_ram[1229] = 0;
    exp_54_ram[1230] = 0;
    exp_54_ram[1231] = 253;
    exp_54_ram[1232] = 0;
    exp_54_ram[1233] = 231;
    exp_54_ram[1234] = 0;
    exp_54_ram[1235] = 0;
    exp_54_ram[1236] = 22;
    exp_54_ram[1237] = 201;
    exp_54_ram[1238] = 0;
    exp_54_ram[1239] = 1;
    exp_54_ram[1240] = 1;
    exp_54_ram[1241] = 0;
    exp_54_ram[1242] = 0;
    exp_54_ram[1243] = 249;
    exp_54_ram[1244] = 0;
    exp_54_ram[1245] = 0;
    exp_54_ram[1246] = 0;
    exp_54_ram[1247] = 0;
    exp_54_ram[1248] = 64;
    exp_54_ram[1249] = 0;
    exp_54_ram[1250] = 0;
    exp_54_ram[1251] = 0;
    exp_54_ram[1252] = 64;
    exp_54_ram[1253] = 0;
    exp_54_ram[1254] = 0;
    exp_54_ram[1255] = 0;
    exp_54_ram[1256] = 65;
    exp_54_ram[1257] = 65;
    exp_54_ram[1258] = 0;
    exp_54_ram[1259] = 0;
    exp_54_ram[1260] = 0;
    exp_54_ram[1261] = 0;
    exp_54_ram[1262] = 0;
    exp_54_ram[1263] = 65;
    exp_54_ram[1264] = 0;
    exp_54_ram[1265] = 0;
    exp_54_ram[1266] = 0;
    exp_54_ram[1267] = 24;
    exp_54_ram[1268] = 255;
    exp_54_ram[1269] = 0;
    exp_54_ram[1270] = 193;
    exp_54_ram[1271] = 0;
    exp_54_ram[1272] = 65;
    exp_54_ram[1273] = 0;
    exp_54_ram[1274] = 0;
    exp_54_ram[1275] = 1;
    exp_54_ram[1276] = 0;
    exp_54_ram[1277] = 1;
    exp_54_ram[1278] = 0;
    exp_54_ram[1279] = 1;
    exp_54_ram[1280] = 0;
    exp_54_ram[1281] = 1;
    exp_54_ram[1282] = 1;
    exp_54_ram[1283] = 1;
    exp_54_ram[1284] = 0;
    exp_54_ram[1285] = 0;
    exp_54_ram[1286] = 0;
    exp_54_ram[1287] = 0;
    exp_54_ram[1288] = 2;
    exp_54_ram[1289] = 0;
    exp_54_ram[1290] = 255;
    exp_54_ram[1291] = 0;
    exp_54_ram[1292] = 0;
    exp_54_ram[1293] = 0;
    exp_54_ram[1294] = 227;
    exp_54_ram[1295] = 0;
    exp_54_ram[1296] = 12;
    exp_54_ram[1297] = 0;
    exp_54_ram[1298] = 196;
    exp_54_ram[1299] = 0;
    exp_54_ram[1300] = 20;
    exp_54_ram[1301] = 0;
    exp_54_ram[1302] = 0;
    exp_54_ram[1303] = 0;
    exp_54_ram[1304] = 0;
    exp_54_ram[1305] = 0;
    exp_54_ram[1306] = 0;
    exp_54_ram[1307] = 0;
    exp_54_ram[1308] = 1;
    exp_54_ram[1309] = 0;
    exp_54_ram[1310] = 255;
    exp_54_ram[1311] = 0;
    exp_54_ram[1312] = 0;
    exp_54_ram[1313] = 0;
    exp_54_ram[1314] = 1;
    exp_54_ram[1315] = 0;
    exp_54_ram[1316] = 0;
    exp_54_ram[1317] = 221;
    exp_54_ram[1318] = 0;
    exp_54_ram[1319] = 12;
    exp_54_ram[1320] = 0;
    exp_54_ram[1321] = 0;
    exp_54_ram[1322] = 190;
    exp_54_ram[1323] = 64;
    exp_54_ram[1324] = 0;
    exp_54_ram[1325] = 64;
    exp_54_ram[1326] = 20;
    exp_54_ram[1327] = 64;
    exp_54_ram[1328] = 0;
    exp_54_ram[1329] = 0;
    exp_54_ram[1330] = 0;
    exp_54_ram[1331] = 0;
    exp_54_ram[1332] = 0;
    exp_54_ram[1333] = 0;
    exp_54_ram[1334] = 1;
    exp_54_ram[1335] = 0;
    exp_54_ram[1336] = 249;
    exp_54_ram[1337] = 0;
    exp_54_ram[1338] = 6;
    exp_54_ram[1339] = 1;
    exp_54_ram[1340] = 0;
    exp_54_ram[1341] = 12;
    exp_54_ram[1342] = 1;
    exp_54_ram[1343] = 6;
    exp_54_ram[1344] = 6;
    exp_54_ram[1345] = 7;
    exp_54_ram[1346] = 5;
    exp_54_ram[1347] = 5;
    exp_54_ram[1348] = 129;
    exp_54_ram[1349] = 0;
    exp_54_ram[1350] = 2;
    exp_54_ram[1351] = 14;
    exp_54_ram[1352] = 2;
    exp_54_ram[1353] = 128;
    exp_54_ram[1354] = 1;
    exp_54_ram[1355] = 0;
    exp_54_ram[1356] = 16;
    exp_54_ram[1357] = 0;
    exp_54_ram[1358] = 0;
    exp_54_ram[1359] = 1;
    exp_54_ram[1360] = 2;
    exp_54_ram[1361] = 0;
    exp_54_ram[1362] = 0;
    exp_54_ram[1363] = 16;
    exp_54_ram[1364] = 253;
    exp_54_ram[1365] = 1;
    exp_54_ram[1366] = 1;
    exp_54_ram[1367] = 0;
    exp_54_ram[1368] = 0;
    exp_54_ram[1369] = 0;
    exp_54_ram[1370] = 0;
    exp_54_ram[1371] = 2;
    exp_54_ram[1372] = 0;
    exp_54_ram[1373] = 251;
    exp_54_ram[1374] = 1;
    exp_54_ram[1375] = 0;
    exp_54_ram[1376] = 0;
    exp_54_ram[1377] = 3;
    exp_54_ram[1378] = 47;
    exp_54_ram[1379] = 0;
    exp_54_ram[1380] = 0;
    exp_54_ram[1381] = 0;
    exp_54_ram[1382] = 1;
    exp_54_ram[1383] = 3;
    exp_54_ram[1384] = 0;
    exp_54_ram[1385] = 0;
    exp_54_ram[1386] = 0;
    exp_54_ram[1387] = 3;
    exp_54_ram[1388] = 0;
    exp_54_ram[1389] = 0;
    exp_54_ram[1390] = 44;
    exp_54_ram[1391] = 0;
    exp_54_ram[1392] = 0;
    exp_54_ram[1393] = 0;
    exp_54_ram[1394] = 1;
    exp_54_ram[1395] = 3;
    exp_54_ram[1396] = 0;
    exp_54_ram[1397] = 0;
    exp_54_ram[1398] = 0;
    exp_54_ram[1399] = 3;
    exp_54_ram[1400] = 0;
    exp_54_ram[1401] = 0;
    exp_54_ram[1402] = 41;
    exp_54_ram[1403] = 0;
    exp_54_ram[1404] = 0;
    exp_54_ram[1405] = 0;
    exp_54_ram[1406] = 1;
    exp_54_ram[1407] = 3;
    exp_54_ram[1408] = 0;
    exp_54_ram[1409] = 0;
    exp_54_ram[1410] = 0;
    exp_54_ram[1411] = 3;
    exp_54_ram[1412] = 0;
    exp_54_ram[1413] = 0;
    exp_54_ram[1414] = 38;
    exp_54_ram[1415] = 0;
    exp_54_ram[1416] = 0;
    exp_54_ram[1417] = 0;
    exp_54_ram[1418] = 1;
    exp_54_ram[1419] = 3;
    exp_54_ram[1420] = 0;
    exp_54_ram[1421] = 0;
    exp_54_ram[1422] = 62;
    exp_54_ram[1423] = 3;
    exp_54_ram[1424] = 0;
    exp_54_ram[1425] = 1;
    exp_54_ram[1426] = 118;
    exp_54_ram[1427] = 35;
    exp_54_ram[1428] = 0;
    exp_54_ram[1429] = 0;
    exp_54_ram[1430] = 0;
    exp_54_ram[1431] = 0;
    exp_54_ram[1432] = 6;
    exp_54_ram[1433] = 3;
    exp_54_ram[1434] = 0;
    exp_54_ram[1435] = 33;
    exp_54_ram[1436] = 0;
    exp_54_ram[1437] = 0;
    exp_54_ram[1438] = 0;
    exp_54_ram[1439] = 0;
    exp_54_ram[1440] = 0;
    exp_54_ram[1441] = 3;
    exp_54_ram[1442] = 0;
    exp_54_ram[1443] = 31;
    exp_54_ram[1444] = 0;
    exp_54_ram[1445] = 0;
    exp_54_ram[1446] = 0;
    exp_54_ram[1447] = 6;
    exp_54_ram[1448] = 3;
    exp_54_ram[1449] = 0;
    exp_54_ram[1450] = 0;
    exp_54_ram[1451] = 6;
    exp_54_ram[1452] = 6;
    exp_54_ram[1453] = 3;
    exp_54_ram[1454] = 0;
    exp_54_ram[1455] = 0;
    exp_54_ram[1456] = 0;
    exp_54_ram[1457] = 6;
    exp_54_ram[1458] = 5;
    exp_54_ram[1459] = 16;
    exp_54_ram[1460] = 5;
    exp_54_ram[1461] = 7;
    exp_54_ram[1462] = 0;
    exp_54_ram[1463] = 252;
    exp_54_ram[1464] = 3;
    exp_54_ram[1465] = 0;
    exp_54_ram[1466] = 2;
    exp_54_ram[1467] = 2;
    exp_54_ram[1468] = 3;
    exp_54_ram[1469] = 3;
    exp_54_ram[1470] = 3;
    exp_54_ram[1471] = 2;
    exp_54_ram[1472] = 3;
    exp_54_ram[1473] = 1;
    exp_54_ram[1474] = 1;
    exp_54_ram[1475] = 1;
    exp_54_ram[1476] = 0;
    exp_54_ram[1477] = 0;
    exp_54_ram[1478] = 0;
    exp_54_ram[1479] = 123;
    exp_54_ram[1480] = 0;
    exp_54_ram[1481] = 24;
    exp_54_ram[1482] = 0;
    exp_54_ram[1483] = 169;
    exp_54_ram[1484] = 0;
    exp_54_ram[1485] = 22;
    exp_54_ram[1486] = 0;
    exp_54_ram[1487] = 0;
    exp_54_ram[1488] = 138;
    exp_54_ram[1489] = 0;
    exp_54_ram[1490] = 0;
    exp_54_ram[1491] = 2;
    exp_54_ram[1492] = 64;
    exp_54_ram[1493] = 0;
    exp_54_ram[1494] = 1;
    exp_54_ram[1495] = 0;
    exp_54_ram[1496] = 64;
    exp_54_ram[1497] = 0;
    exp_54_ram[1498] = 252;
    exp_54_ram[1499] = 0;
    exp_54_ram[1500] = 0;
    exp_54_ram[1501] = 0;
    exp_54_ram[1502] = 24;
    exp_54_ram[1503] = 0;
    exp_54_ram[1504] = 0;
    exp_54_ram[1505] = 169;
    exp_54_ram[1506] = 0;
    exp_54_ram[1507] = 0;
    exp_54_ram[1508] = 0;
    exp_54_ram[1509] = 0;
    exp_54_ram[1510] = 133;
    exp_54_ram[1511] = 0;
    exp_54_ram[1512] = 2;
    exp_54_ram[1513] = 64;
    exp_54_ram[1514] = 0;
    exp_54_ram[1515] = 1;
    exp_54_ram[1516] = 1;
    exp_54_ram[1517] = 0;
    exp_54_ram[1518] = 64;
    exp_54_ram[1519] = 252;
    exp_54_ram[1520] = 0;
    exp_54_ram[1521] = 0;
    exp_54_ram[1522] = 24;
    exp_54_ram[1523] = 11;
    exp_54_ram[1524] = 0;
    exp_54_ram[1525] = 0;
    exp_54_ram[1526] = 0;
    exp_54_ram[1527] = 0;
    exp_54_ram[1528] = 0;
    exp_54_ram[1529] = 0;
    exp_54_ram[1530] = 225;
    exp_54_ram[1531] = 9;
    exp_54_ram[1532] = 0;
    exp_54_ram[1533] = 0;
    exp_54_ram[1534] = 0;
    exp_54_ram[1535] = 0;
    exp_54_ram[1536] = 3;
    exp_54_ram[1537] = 137;
    exp_54_ram[1538] = 7;
    exp_54_ram[1539] = 0;
    exp_54_ram[1540] = 0;
    exp_54_ram[1541] = 0;
    exp_54_ram[1542] = 0;
    exp_54_ram[1543] = 0;
    exp_54_ram[1544] = 1;
    exp_54_ram[1545] = 1;
    exp_54_ram[1546] = 1;
    exp_54_ram[1547] = 0;
    exp_54_ram[1548] = 0;
    exp_54_ram[1549] = 0;
    exp_54_ram[1550] = 133;
    exp_54_ram[1551] = 0;
    exp_54_ram[1552] = 1;
    exp_54_ram[1553] = 3;
    exp_54_ram[1554] = 0;
    exp_54_ram[1555] = 3;
    exp_54_ram[1556] = 3;
    exp_54_ram[1557] = 3;
    exp_54_ram[1558] = 2;
    exp_54_ram[1559] = 2;
    exp_54_ram[1560] = 2;
    exp_54_ram[1561] = 2;
    exp_54_ram[1562] = 1;
    exp_54_ram[1563] = 1;
    exp_54_ram[1564] = 1;
    exp_54_ram[1565] = 4;
    exp_54_ram[1566] = 0;
    exp_54_ram[1567] = 246;
    exp_54_ram[1568] = 9;
    exp_54_ram[1569] = 1;
    exp_54_ram[1570] = 0;
    exp_54_ram[1571] = 8;
    exp_54_ram[1572] = 9;
    exp_54_ram[1573] = 9;
    exp_54_ram[1574] = 1;
    exp_54_ram[1575] = 0;
    exp_54_ram[1576] = 2;
    exp_54_ram[1577] = 0;
    exp_54_ram[1578] = 3;
    exp_54_ram[1579] = 0;
    exp_54_ram[1580] = 8;
    exp_54_ram[1581] = 4;
    exp_54_ram[1582] = 8;
    exp_54_ram[1583] = 9;
    exp_54_ram[1584] = 5;
    exp_54_ram[1585] = 4;
    exp_54_ram[1586] = 5;
    exp_54_ram[1587] = 2;
    exp_54_ram[1588] = 2;
    exp_54_ram[1589] = 4;
    exp_54_ram[1590] = 197;
    exp_54_ram[1591] = 0;
    exp_54_ram[1592] = 157;
    exp_54_ram[1593] = 0;
    exp_54_ram[1594] = 0;
    exp_54_ram[1595] = 3;
    exp_54_ram[1596] = 222;
    exp_54_ram[1597] = 5;
    exp_54_ram[1598] = 4;
    exp_54_ram[1599] = 2;
    exp_54_ram[1600] = 3;
    exp_54_ram[1601] = 64;
    exp_54_ram[1602] = 0;
    exp_54_ram[1603] = 4;
    exp_54_ram[1604] = 193;
    exp_54_ram[1605] = 0;
    exp_54_ram[1606] = 154;
    exp_54_ram[1607] = 0;
    exp_54_ram[1608] = 2;
    exp_54_ram[1609] = 0;
    exp_54_ram[1610] = 0;
    exp_54_ram[1611] = 0;
    exp_54_ram[1612] = 5;
    exp_54_ram[1613] = 6;
    exp_54_ram[1614] = 7;
    exp_54_ram[1615] = 6;
    exp_54_ram[1616] = 7;
    exp_54_ram[1617] = 6;
    exp_54_ram[1618] = 4;
    exp_54_ram[1619] = 189;
    exp_54_ram[1620] = 0;
    exp_54_ram[1621] = 150;
    exp_54_ram[1622] = 0;
    exp_54_ram[1623] = 0;
    exp_54_ram[1624] = 5;
    exp_54_ram[1625] = 215;
    exp_54_ram[1626] = 7;
    exp_54_ram[1627] = 6;
    exp_54_ram[1628] = 2;
    exp_54_ram[1629] = 5;
    exp_54_ram[1630] = 64;
    exp_54_ram[1631] = 0;
    exp_54_ram[1632] = 6;
    exp_54_ram[1633] = 186;
    exp_54_ram[1634] = 0;
    exp_54_ram[1635] = 146;
    exp_54_ram[1636] = 0;
    exp_54_ram[1637] = 0;
    exp_54_ram[1638] = 2;
    exp_54_ram[1639] = 0;
    exp_54_ram[1640] = 0;
    exp_54_ram[1641] = 184;
    exp_54_ram[1642] = 0;
    exp_54_ram[1643] = 144;
    exp_54_ram[1644] = 2;
    exp_54_ram[1645] = 0;
    exp_54_ram[1646] = 0;
    exp_54_ram[1647] = 0;
    exp_54_ram[1648] = 1;
    exp_54_ram[1649] = 0;
    exp_54_ram[1650] = 0;
    exp_54_ram[1651] = 0;
    exp_54_ram[1652] = 1;
    exp_54_ram[1653] = 0;
    exp_54_ram[1654] = 9;
    exp_54_ram[1655] = 9;
    exp_54_ram[1656] = 9;
    exp_54_ram[1657] = 9;
    exp_54_ram[1658] = 8;
    exp_54_ram[1659] = 8;
    exp_54_ram[1660] = 8;
    exp_54_ram[1661] = 10;
    exp_54_ram[1662] = 0;
    exp_54_ram[1663] = 248;
    exp_54_ram[1664] = 0;
    exp_54_ram[1665] = 7;
    exp_54_ram[1666] = 2;
    exp_54_ram[1667] = 0;
    exp_54_ram[1668] = 3;
    exp_54_ram[1669] = 6;
    exp_54_ram[1670] = 6;
    exp_54_ram[1671] = 6;
    exp_54_ram[1672] = 7;
    exp_54_ram[1673] = 176;
    exp_54_ram[1674] = 2;
    exp_54_ram[1675] = 3;
    exp_54_ram[1676] = 0;
    exp_54_ram[1677] = 2;
    exp_54_ram[1678] = 175;
    exp_54_ram[1679] = 0;
    exp_54_ram[1680] = 135;
    exp_54_ram[1681] = 0;
    exp_54_ram[1682] = 0;
    exp_54_ram[1683] = 7;
    exp_54_ram[1684] = 255;
    exp_54_ram[1685] = 31;
    exp_54_ram[1686] = 0;
    exp_54_ram[1687] = 0;
    exp_54_ram[1688] = 255;
    exp_54_ram[1689] = 0;
    exp_54_ram[1690] = 0;
    exp_54_ram[1691] = 0;
    exp_54_ram[1692] = 0;
    exp_54_ram[1693] = 0;
    exp_54_ram[1694] = 198;
    exp_54_ram[1695] = 2;
    exp_54_ram[1696] = 0;
    exp_54_ram[1697] = 0;
    exp_54_ram[1698] = 170;
    exp_54_ram[1699] = 7;
    exp_54_ram[1700] = 0;
    exp_54_ram[1701] = 2;
    exp_54_ram[1702] = 7;
    exp_54_ram[1703] = 0;
    exp_54_ram[1704] = 7;
    exp_54_ram[1705] = 7;
    exp_54_ram[1706] = 6;
    exp_54_ram[1707] = 0;
    exp_54_ram[1708] = 7;
    exp_54_ram[1709] = 8;
    exp_54_ram[1710] = 0;
    exp_54_ram[1711] = 250;
    exp_54_ram[1712] = 2;
    exp_54_ram[1713] = 3;
    exp_54_ram[1714] = 0;
    exp_54_ram[1715] = 165;
    exp_54_ram[1716] = 0;
    exp_54_ram[1717] = 218;
    exp_54_ram[1718] = 0;
    exp_54_ram[1719] = 0;
    exp_54_ram[1720] = 0;
    exp_54_ram[1721] = 225;
    exp_54_ram[1722] = 64;
    exp_54_ram[1723] = 0;
    exp_54_ram[1724] = 64;
    exp_54_ram[1725] = 0;
    exp_54_ram[1726] = 247;
    exp_54_ram[1727] = 2;
    exp_54_ram[1728] = 2;
    exp_54_ram[1729] = 3;
    exp_54_ram[1730] = 0;
    exp_54_ram[1731] = 161;
    exp_54_ram[1732] = 0;
    exp_54_ram[1733] = 214;
    exp_54_ram[1734] = 2;
    exp_54_ram[1735] = 247;
    exp_54_ram[1736] = 2;
    exp_54_ram[1737] = 247;
    exp_54_ram[1738] = 249;
    exp_54_ram[1739] = 0;
    exp_54_ram[1740] = 0;
    exp_54_ram[1741] = 3;
    exp_54_ram[1742] = 6;
    exp_54_ram[1743] = 186;
    exp_54_ram[1744] = 3;
    exp_54_ram[1745] = 2;
    exp_54_ram[1746] = 0;
    exp_54_ram[1747] = 157;
    exp_54_ram[1748] = 0;
    exp_54_ram[1749] = 210;
    exp_54_ram[1750] = 6;
    exp_54_ram[1751] = 7;
    exp_54_ram[1752] = 0;
    exp_54_ram[1753] = 0;
    exp_54_ram[1754] = 0;
    exp_54_ram[1755] = 252;
    exp_54_ram[1756] = 0;
    exp_54_ram[1757] = 2;
    exp_54_ram[1758] = 2;
    exp_54_ram[1759] = 182;
    exp_54_ram[1760] = 0;
    exp_54_ram[1761] = 0;
    exp_54_ram[1762] = 18;
    exp_54_ram[1763] = 2;
    exp_54_ram[1764] = 153;
    exp_54_ram[1765] = 3;
    exp_54_ram[1766] = 18;
    exp_54_ram[1767] = 3;
    exp_54_ram[1768] = 4;
    exp_54_ram[1769] = 0;
    exp_54_ram[1770] = 251;
    exp_54_ram[1771] = 4;
    exp_54_ram[1772] = 5;
    exp_54_ram[1773] = 0;
    exp_54_ram[1774] = 0;
    exp_54_ram[1775] = 4;
    exp_54_ram[1776] = 0;
    exp_54_ram[1777] = 0;
    exp_54_ram[1778] = 4;
    exp_54_ram[1779] = 3;
    exp_54_ram[1780] = 245;
    exp_54_ram[1781] = 0;
    exp_54_ram[1782] = 0;
    exp_54_ram[1783] = 0;
    exp_54_ram[1784] = 225;
    exp_54_ram[1785] = 1;
    exp_54_ram[1786] = 0;
    exp_54_ram[1787] = 0;
    exp_54_ram[1788] = 0;
    exp_54_ram[1789] = 174;
    exp_54_ram[1790] = 0;
    exp_54_ram[1791] = 0;
    exp_54_ram[1792] = 2;
    exp_54_ram[1793] = 18;
    exp_54_ram[1794] = 146;
    exp_54_ram[1795] = 0;
    exp_54_ram[1796] = 0;
    exp_54_ram[1797] = 241;
    exp_54_ram[1798] = 18;
    exp_54_ram[1799] = 2;
    exp_54_ram[1800] = 4;
    exp_54_ram[1801] = 18;
    exp_54_ram[1802] = 4;
    exp_54_ram[1803] = 4;
    exp_54_ram[1804] = 4;
    exp_54_ram[1805] = 3;
    exp_54_ram[1806] = 5;
    exp_54_ram[1807] = 0;
    exp_54_ram[1808] = 255;
    exp_54_ram[1809] = 0;
    exp_54_ram[1810] = 246;
    exp_54_ram[1811] = 0;
    exp_54_ram[1812] = 1;
    exp_54_ram[1813] = 136;
    exp_54_ram[1814] = 254;
    exp_54_ram[1815] = 0;
    exp_54_ram[1816] = 0;
    exp_54_ram[1817] = 2;
    exp_54_ram[1818] = 0;
    exp_54_ram[1819] = 152;
    exp_54_ram[1820] = 136;
    exp_54_ram[1821] = 254;
    exp_54_ram[1822] = 0;
    exp_54_ram[1823] = 84;
    exp_54_ram[1824] = 0;
    exp_54_ram[1825] = 0;
    exp_54_ram[1826] = 254;
    exp_54_ram[1827] = 0;
    exp_54_ram[1828] = 160;
    exp_54_ram[1829] = 0;
    exp_54_ram[1830] = 0;
    exp_54_ram[1831] = 254;
    exp_54_ram[1832] = 0;
    exp_54_ram[1833] = 0;
    exp_54_ram[1834] = 152;
    exp_54_ram[1835] = 152;
    exp_54_ram[1836] = 0;
    exp_54_ram[1837] = 152;
    exp_54_ram[1838] = 0;
    exp_54_ram[1839] = 152;
    exp_54_ram[1840] = 0;
    exp_54_ram[1841] = 0;
    exp_54_ram[1842] = 0;
    exp_54_ram[1843] = 0;
    exp_54_ram[1844] = 0;
    exp_54_ram[1845] = 254;
    exp_54_ram[1846] = 0;
    exp_54_ram[1847] = 153;
    exp_54_ram[1848] = 0;
    exp_54_ram[1849] = 148;
    exp_54_ram[1850] = 0;
    exp_54_ram[1851] = 0;
    exp_54_ram[1852] = 0;
    exp_54_ram[1853] = 153;
    exp_54_ram[1854] = 255;
    exp_54_ram[1855] = 63;
    exp_54_ram[1856] = 254;
    exp_54_ram[1857] = 254;
    exp_54_ram[1858] = 0;
    exp_54_ram[1859] = 153;
    exp_54_ram[1860] = 0;
    exp_54_ram[1861] = 0;
    exp_54_ram[1862] = 254;
    exp_54_ram[1863] = 0;
    exp_54_ram[1864] = 0;
    exp_54_ram[1865] = 152;
    exp_54_ram[1866] = 152;
    exp_54_ram[1867] = 0;
    exp_54_ram[1868] = 152;
    exp_54_ram[1869] = 0;
    exp_54_ram[1870] = 152;
    exp_54_ram[1871] = 0;
    exp_54_ram[1872] = 0;
    exp_54_ram[1873] = 0;
    exp_54_ram[1874] = 0;
    exp_54_ram[1875] = 0;
    exp_54_ram[1876] = 254;
    exp_54_ram[1877] = 0;
    exp_54_ram[1878] = 152;
    exp_54_ram[1879] = 0;
    exp_54_ram[1880] = 140;
    exp_54_ram[1881] = 0;
    exp_54_ram[1882] = 0;
    exp_54_ram[1883] = 0;
    exp_54_ram[1884] = 154;
    exp_54_ram[1885] = 247;
    exp_54_ram[1886] = 56;
    exp_54_ram[1887] = 254;
    exp_54_ram[1888] = 0;
    exp_54_ram[1889] = 84;
    exp_54_ram[1890] = 0;
    exp_54_ram[1891] = 0;
    exp_54_ram[1892] = 254;
    exp_54_ram[1893] = 0;
    exp_54_ram[1894] = 154;
    exp_54_ram[1895] = 0;
    exp_54_ram[1896] = 136;
    exp_54_ram[1897] = 0;
    exp_54_ram[1898] = 0;
    exp_54_ram[1899] = 0;
    exp_54_ram[1900] = 154;
    exp_54_ram[1901] = 243;
    exp_54_ram[1902] = 52;
    exp_54_ram[1903] = 254;
    exp_54_ram[1904] = 254;
    exp_54_ram[1905] = 0;
    exp_54_ram[1906] = 0;
    exp_54_ram[1907] = 0;
    exp_54_ram[1908] = 155;
    exp_54_ram[1909] = 241;
    exp_54_ram[1910] = 50;
    exp_54_ram[1911] = 0;
    exp_54_ram[1912] = 155;
    exp_54_ram[1913] = 240;
    exp_54_ram[1914] = 0;
    exp_54_ram[1915] = 156;
    exp_54_ram[1916] = 240;
    exp_54_ram[1917] = 254;
    exp_54_ram[1918] = 0;
    exp_54_ram[1919] = 84;
    exp_54_ram[1920] = 0;
    exp_54_ram[1921] = 0;
    exp_54_ram[1922] = 254;
    exp_54_ram[1923] = 0;
    exp_54_ram[1924] = 0;
    exp_54_ram[1925] = 157;
    exp_54_ram[1926] = 0;
    exp_54_ram[1927] = 252;
    exp_54_ram[1928] = 0;
    exp_54_ram[1929] = 0;
    exp_54_ram[1930] = 153;
    exp_54_ram[1931] = 0;
    exp_54_ram[1932] = 255;
    exp_54_ram[1933] = 0;
    exp_54_ram[1934] = 0;
    exp_54_ram[1935] = 0;
    exp_54_ram[1936] = 153;
    exp_54_ram[1937] = 234;
    exp_54_ram[1938] = 43;
    exp_54_ram[1939] = 254;
    exp_54_ram[1940] = 254;
    exp_54_ram[1941] = 0;
    exp_54_ram[1942] = 0;
    exp_54_ram[1943] = 157;
    exp_54_ram[1944] = 0;
    exp_54_ram[1945] = 247;
    exp_54_ram[1946] = 0;
    exp_54_ram[1947] = 0;
    exp_54_ram[1948] = 152;
    exp_54_ram[1949] = 0;
    exp_54_ram[1950] = 251;
    exp_54_ram[1951] = 0;
    exp_54_ram[1952] = 0;
    exp_54_ram[1953] = 0;
    exp_54_ram[1954] = 154;
    exp_54_ram[1955] = 230;
    exp_54_ram[1956] = 38;
    exp_54_ram[1957] = 254;
    exp_54_ram[1958] = 0;
    exp_54_ram[1959] = 84;
    exp_54_ram[1960] = 0;
    exp_54_ram[1961] = 0;
    exp_54_ram[1962] = 254;
    exp_54_ram[1963] = 0;
    exp_54_ram[1964] = 154;
    exp_54_ram[1965] = 0;
    exp_54_ram[1966] = 247;
    exp_54_ram[1967] = 0;
    exp_54_ram[1968] = 0;
    exp_54_ram[1969] = 0;
    exp_54_ram[1970] = 154;
    exp_54_ram[1971] = 226;
    exp_54_ram[1972] = 34;
    exp_54_ram[1973] = 254;
    exp_54_ram[1974] = 254;
    exp_54_ram[1975] = 0;
    exp_54_ram[1976] = 0;
    exp_54_ram[1977] = 0;
    exp_54_ram[1978] = 155;
    exp_54_ram[1979] = 224;
    exp_54_ram[1980] = 32;
    exp_54_ram[1981] = 0;
    exp_54_ram[1982] = 155;
    exp_54_ram[1983] = 223;
    exp_54_ram[1984] = 0;
    exp_54_ram[1985] = 157;
    exp_54_ram[1986] = 222;
    exp_54_ram[1987] = 0;
    exp_54_ram[1988] = 155;
    exp_54_ram[1989] = 221;
    exp_54_ram[1990] = 0;
    exp_54_ram[1991] = 158;
    exp_54_ram[1992] = 221;
    exp_54_ram[1993] = 0;
    exp_54_ram[1994] = 155;
    exp_54_ram[1995] = 220;
    exp_54_ram[1996] = 0;
    exp_54_ram[1997] = 159;
    exp_54_ram[1998] = 219;
    exp_54_ram[1999] = 0;
    exp_54_ram[2000] = 155;
    exp_54_ram[2001] = 218;
    exp_54_ram[2002] = 0;
    exp_54_ram[2003] = 159;
    exp_54_ram[2004] = 218;
    exp_54_ram[2005] = 254;
    exp_54_ram[2006] = 52;
    exp_54_ram[2007] = 35;
    exp_54_ram[2008] = 0;
    exp_54_ram[2009] = 0;
    exp_54_ram[2010] = 254;
    exp_54_ram[2011] = 0;
    exp_54_ram[2012] = 3;
    exp_54_ram[2013] = 0;
    exp_54_ram[2014] = 246;
    exp_54_ram[2015] = 0;
    exp_54_ram[2016] = 254;
    exp_54_ram[2017] = 0;
    exp_54_ram[2018] = 0;
    exp_54_ram[2019] = 153;
    exp_54_ram[2020] = 214;
    exp_54_ram[2021] = 22;
    exp_54_ram[2022] = 254;
    exp_54_ram[2023] = 0;
    exp_54_ram[2024] = 3;
    exp_54_ram[2025] = 0;
    exp_54_ram[2026] = 243;
    exp_54_ram[2027] = 0;
    exp_54_ram[2028] = 254;
    exp_54_ram[2029] = 64;
    exp_54_ram[2030] = 0;
    exp_54_ram[2031] = 0;
    exp_54_ram[2032] = 0;
    exp_54_ram[2033] = 154;
    exp_54_ram[2034] = 210;
    exp_54_ram[2035] = 18;
    exp_54_ram[2036] = 254;
    exp_54_ram[2037] = 0;
    exp_54_ram[2038] = 3;
    exp_54_ram[2039] = 0;
    exp_54_ram[2040] = 239;
    exp_54_ram[2041] = 0;
    exp_54_ram[2042] = 254;
    exp_54_ram[2043] = 64;
    exp_54_ram[2044] = 0;
    exp_54_ram[2045] = 0;
    exp_54_ram[2046] = 0;
    exp_54_ram[2047] = 154;
    exp_54_ram[2048] = 207;
    exp_54_ram[2049] = 15;
    exp_54_ram[2050] = 254;
    exp_54_ram[2051] = 0;
    exp_54_ram[2052] = 3;
    exp_54_ram[2053] = 0;
    exp_54_ram[2054] = 236;
    exp_54_ram[2055] = 0;
    exp_54_ram[2056] = 254;
    exp_54_ram[2057] = 64;
    exp_54_ram[2058] = 0;
    exp_54_ram[2059] = 0;
    exp_54_ram[2060] = 0;
    exp_54_ram[2061] = 155;
    exp_54_ram[2062] = 203;
    exp_54_ram[2063] = 11;
    exp_54_ram[2064] = 254;
    exp_54_ram[2065] = 0;
    exp_54_ram[2066] = 3;
    exp_54_ram[2067] = 0;
    exp_54_ram[2068] = 232;
    exp_54_ram[2069] = 0;
    exp_54_ram[2070] = 0;
    exp_54_ram[2071] = 0;
    exp_54_ram[2072] = 160;
    exp_54_ram[2073] = 200;
    exp_54_ram[2074] = 9;
    exp_54_ram[2075] = 0;
    exp_54_ram[2076] = 155;
    exp_54_ram[2077] = 199;
    exp_54_ram[2078] = 0;
    exp_54_ram[2079] = 161;
    exp_54_ram[2080] = 199;
    exp_54_ram[2081] = 254;
    exp_54_ram[2082] = 52;
    exp_54_ram[2083] = 35;
    exp_54_ram[2084] = 0;
    exp_54_ram[2085] = 52;
    exp_54_ram[2086] = 35;
    exp_54_ram[2087] = 0;
    exp_54_ram[2088] = 0;
    exp_54_ram[2089] = 254;
    exp_54_ram[2090] = 3;
    exp_54_ram[2091] = 0;
    exp_54_ram[2092] = 229;
    exp_54_ram[2093] = 0;
    exp_54_ram[2094] = 254;
    exp_54_ram[2095] = 0;
    exp_54_ram[2096] = 0;
    exp_54_ram[2097] = 153;
    exp_54_ram[2098] = 194;
    exp_54_ram[2099] = 2;
    exp_54_ram[2100] = 254;
    exp_54_ram[2101] = 3;
    exp_54_ram[2102] = 0;
    exp_54_ram[2103] = 226;
    exp_54_ram[2104] = 0;
    exp_54_ram[2105] = 254;
    exp_54_ram[2106] = 64;
    exp_54_ram[2107] = 0;
    exp_54_ram[2108] = 0;
    exp_54_ram[2109] = 0;
    exp_54_ram[2110] = 154;
    exp_54_ram[2111] = 191;
    exp_54_ram[2112] = 127;
    exp_54_ram[2113] = 254;
    exp_54_ram[2114] = 3;
    exp_54_ram[2115] = 0;
    exp_54_ram[2116] = 223;
    exp_54_ram[2117] = 0;
    exp_54_ram[2118] = 254;
    exp_54_ram[2119] = 64;
    exp_54_ram[2120] = 0;
    exp_54_ram[2121] = 0;
    exp_54_ram[2122] = 0;
    exp_54_ram[2123] = 154;
    exp_54_ram[2124] = 188;
    exp_54_ram[2125] = 124;
    exp_54_ram[2126] = 254;
    exp_54_ram[2127] = 3;
    exp_54_ram[2128] = 0;
    exp_54_ram[2129] = 219;
    exp_54_ram[2130] = 0;
    exp_54_ram[2131] = 254;
    exp_54_ram[2132] = 64;
    exp_54_ram[2133] = 0;
    exp_54_ram[2134] = 0;
    exp_54_ram[2135] = 0;
    exp_54_ram[2136] = 155;
    exp_54_ram[2137] = 184;
    exp_54_ram[2138] = 121;
    exp_54_ram[2139] = 254;
    exp_54_ram[2140] = 0;
    exp_54_ram[2141] = 210;
    exp_54_ram[2142] = 0;
    exp_54_ram[2143] = 0;
    exp_54_ram[2144] = 254;
    exp_54_ram[2145] = 0;
    exp_54_ram[2146] = 254;
    exp_54_ram[2147] = 64;
    exp_54_ram[2148] = 0;
    exp_54_ram[2149] = 0;
    exp_54_ram[2150] = 0;
    exp_54_ram[2151] = 160;
    exp_54_ram[2152] = 181;
    exp_54_ram[2153] = 117;
    exp_54_ram[2154] = 254;
    exp_54_ram[2155] = 3;
    exp_54_ram[2156] = 0;
    exp_54_ram[2157] = 212;
    exp_54_ram[2158] = 0;
    exp_54_ram[2159] = 0;
    exp_54_ram[2160] = 0;
    exp_54_ram[2161] = 161;
    exp_54_ram[2162] = 178;
    exp_54_ram[2163] = 114;
    exp_54_ram[2164] = 0;
    exp_54_ram[2165] = 155;
    exp_54_ram[2166] = 177;
    exp_54_ram[2167] = 0;
    exp_54_ram[2168] = 162;
    exp_54_ram[2169] = 176;
    exp_54_ram[2170] = 254;
    exp_54_ram[2171] = 52;
    exp_54_ram[2172] = 35;
    exp_54_ram[2173] = 0;
    exp_54_ram[2174] = 0;
    exp_54_ram[2175] = 254;
    exp_54_ram[2176] = 0;
    exp_54_ram[2177] = 163;
    exp_54_ram[2178] = 0;
    exp_54_ram[2179] = 226;
    exp_54_ram[2180] = 0;
    exp_54_ram[2181] = 0;
    exp_54_ram[2182] = 0;
    exp_54_ram[2183] = 153;
    exp_54_ram[2184] = 173;
    exp_54_ram[2185] = 109;
    exp_54_ram[2186] = 254;
    exp_54_ram[2187] = 0;
    exp_54_ram[2188] = 163;
    exp_54_ram[2189] = 0;
    exp_54_ram[2190] = 223;
    exp_54_ram[2191] = 0;
    exp_54_ram[2192] = 0;
    exp_54_ram[2193] = 0;
    exp_54_ram[2194] = 0;
    exp_54_ram[2195] = 154;
    exp_54_ram[2196] = 170;
    exp_54_ram[2197] = 106;
    exp_54_ram[2198] = 254;
    exp_54_ram[2199] = 0;
    exp_54_ram[2200] = 164;
    exp_54_ram[2201] = 0;
    exp_54_ram[2202] = 220;
    exp_54_ram[2203] = 0;
    exp_54_ram[2204] = 0;
    exp_54_ram[2205] = 0;
    exp_54_ram[2206] = 0;
    exp_54_ram[2207] = 154;
    exp_54_ram[2208] = 167;
    exp_54_ram[2209] = 103;
    exp_54_ram[2210] = 254;
    exp_54_ram[2211] = 0;
    exp_54_ram[2212] = 165;
    exp_54_ram[2213] = 0;
    exp_54_ram[2214] = 217;
    exp_54_ram[2215] = 0;
    exp_54_ram[2216] = 0;
    exp_54_ram[2217] = 0;
    exp_54_ram[2218] = 0;
    exp_54_ram[2219] = 155;
    exp_54_ram[2220] = 164;
    exp_54_ram[2221] = 100;
    exp_54_ram[2222] = 254;
    exp_54_ram[2223] = 0;
    exp_54_ram[2224] = 165;
    exp_54_ram[2225] = 0;
    exp_54_ram[2226] = 214;
    exp_54_ram[2227] = 0;
    exp_54_ram[2228] = 0;
    exp_54_ram[2229] = 0;
    exp_54_ram[2230] = 0;
    exp_54_ram[2231] = 161;
    exp_54_ram[2232] = 161;
    exp_54_ram[2233] = 97;
    exp_54_ram[2234] = 0;
    exp_54_ram[2235] = 155;
    exp_54_ram[2236] = 160;
    exp_54_ram[2237] = 0;
    exp_54_ram[2238] = 166;
    exp_54_ram[2239] = 159;
    exp_54_ram[2240] = 254;
    exp_54_ram[2241] = 52;
    exp_54_ram[2242] = 35;
    exp_54_ram[2243] = 0;
    exp_54_ram[2244] = 0;
    exp_54_ram[2245] = 254;
    exp_54_ram[2246] = 0;
    exp_54_ram[2247] = 167;
    exp_54_ram[2248] = 0;
    exp_54_ram[2249] = 216;
    exp_54_ram[2250] = 0;
    exp_54_ram[2251] = 254;
    exp_54_ram[2252] = 0;
    exp_54_ram[2253] = 0;
    exp_54_ram[2254] = 153;
    exp_54_ram[2255] = 155;
    exp_54_ram[2256] = 91;
    exp_54_ram[2257] = 254;
    exp_54_ram[2258] = 0;
    exp_54_ram[2259] = 168;
    exp_54_ram[2260] = 0;
    exp_54_ram[2261] = 213;
    exp_54_ram[2262] = 0;
    exp_54_ram[2263] = 254;
    exp_54_ram[2264] = 64;
    exp_54_ram[2265] = 0;
    exp_54_ram[2266] = 0;
    exp_54_ram[2267] = 0;
    exp_54_ram[2268] = 154;
    exp_54_ram[2269] = 151;
    exp_54_ram[2270] = 88;
    exp_54_ram[2271] = 254;
    exp_54_ram[2272] = 0;
    exp_54_ram[2273] = 168;
    exp_54_ram[2274] = 0;
    exp_54_ram[2275] = 210;
    exp_54_ram[2276] = 0;
    exp_54_ram[2277] = 254;
    exp_54_ram[2278] = 64;
    exp_54_ram[2279] = 0;
    exp_54_ram[2280] = 0;
    exp_54_ram[2281] = 0;
    exp_54_ram[2282] = 154;
    exp_54_ram[2283] = 148;
    exp_54_ram[2284] = 84;
    exp_54_ram[2285] = 254;
    exp_54_ram[2286] = 0;
    exp_54_ram[2287] = 169;
    exp_54_ram[2288] = 0;
    exp_54_ram[2289] = 206;
    exp_54_ram[2290] = 0;
    exp_54_ram[2291] = 254;
    exp_54_ram[2292] = 64;
    exp_54_ram[2293] = 0;
    exp_54_ram[2294] = 0;
    exp_54_ram[2295] = 0;
    exp_54_ram[2296] = 155;
    exp_54_ram[2297] = 144;
    exp_54_ram[2298] = 81;
    exp_54_ram[2299] = 254;
    exp_54_ram[2300] = 0;
    exp_54_ram[2301] = 169;
    exp_54_ram[2302] = 0;
    exp_54_ram[2303] = 203;
    exp_54_ram[2304] = 0;
    exp_54_ram[2305] = 0;
    exp_54_ram[2306] = 0;
    exp_54_ram[2307] = 160;
    exp_54_ram[2308] = 142;
    exp_54_ram[2309] = 78;
    exp_54_ram[2310] = 0;
    exp_54_ram[2311] = 155;
    exp_54_ram[2312] = 141;
    exp_54_ram[2313] = 0;
    exp_54_ram[2314] = 170;
    exp_54_ram[2315] = 140;
    exp_54_ram[2316] = 254;
    exp_54_ram[2317] = 52;
    exp_54_ram[2318] = 35;
    exp_54_ram[2319] = 0;
    exp_54_ram[2320] = 52;
    exp_54_ram[2321] = 35;
    exp_54_ram[2322] = 0;
    exp_54_ram[2323] = 0;
    exp_54_ram[2324] = 254;
    exp_54_ram[2325] = 3;
    exp_54_ram[2326] = 0;
    exp_54_ram[2327] = 175;
    exp_54_ram[2328] = 0;
    exp_54_ram[2329] = 254;
    exp_54_ram[2330] = 64;
    exp_54_ram[2331] = 0;
    exp_54_ram[2332] = 0;
    exp_54_ram[2333] = 0;
    exp_54_ram[2334] = 153;
    exp_54_ram[2335] = 135;
    exp_54_ram[2336] = 71;
    exp_54_ram[2337] = 254;
    exp_54_ram[2338] = 3;
    exp_54_ram[2339] = 0;
    exp_54_ram[2340] = 172;
    exp_54_ram[2341] = 0;
    exp_54_ram[2342] = 254;
    exp_54_ram[2343] = 64;
    exp_54_ram[2344] = 0;
    exp_54_ram[2345] = 0;
    exp_54_ram[2346] = 0;
    exp_54_ram[2347] = 154;
    exp_54_ram[2348] = 132;
    exp_54_ram[2349] = 68;
    exp_54_ram[2350] = 254;
    exp_54_ram[2351] = 3;
    exp_54_ram[2352] = 0;
    exp_54_ram[2353] = 169;
    exp_54_ram[2354] = 0;
    exp_54_ram[2355] = 254;
    exp_54_ram[2356] = 64;
    exp_54_ram[2357] = 0;
    exp_54_ram[2358] = 0;
    exp_54_ram[2359] = 0;
    exp_54_ram[2360] = 154;
    exp_54_ram[2361] = 128;
    exp_54_ram[2362] = 65;
    exp_54_ram[2363] = 254;
    exp_54_ram[2364] = 3;
    exp_54_ram[2365] = 0;
    exp_54_ram[2366] = 165;
    exp_54_ram[2367] = 0;
    exp_54_ram[2368] = 254;
    exp_54_ram[2369] = 64;
    exp_54_ram[2370] = 0;
    exp_54_ram[2371] = 0;
    exp_54_ram[2372] = 0;
    exp_54_ram[2373] = 155;
    exp_54_ram[2374] = 253;
    exp_54_ram[2375] = 61;
    exp_54_ram[2376] = 254;
    exp_54_ram[2377] = 0;
    exp_54_ram[2378] = 151;
    exp_54_ram[2379] = 0;
    exp_54_ram[2380] = 0;
    exp_54_ram[2381] = 254;
    exp_54_ram[2382] = 0;
    exp_54_ram[2383] = 254;
    exp_54_ram[2384] = 64;
    exp_54_ram[2385] = 0;
    exp_54_ram[2386] = 0;
    exp_54_ram[2387] = 0;
    exp_54_ram[2388] = 160;
    exp_54_ram[2389] = 249;
    exp_54_ram[2390] = 58;
    exp_54_ram[2391] = 254;
    exp_54_ram[2392] = 3;
    exp_54_ram[2393] = 0;
    exp_54_ram[2394] = 158;
    exp_54_ram[2395] = 0;
    exp_54_ram[2396] = 0;
    exp_54_ram[2397] = 0;
    exp_54_ram[2398] = 161;
    exp_54_ram[2399] = 247;
    exp_54_ram[2400] = 55;
    exp_54_ram[2401] = 0;
    exp_54_ram[2402] = 155;
    exp_54_ram[2403] = 246;
    exp_54_ram[2404] = 0;
    exp_54_ram[2405] = 171;
    exp_54_ram[2406] = 245;
    exp_54_ram[2407] = 254;
    exp_54_ram[2408] = 52;
    exp_54_ram[2409] = 35;
    exp_54_ram[2410] = 0;
    exp_54_ram[2411] = 0;
    exp_54_ram[2412] = 254;
    exp_54_ram[2413] = 0;
    exp_54_ram[2414] = 171;
    exp_54_ram[2415] = 0;
    exp_54_ram[2416] = 158;
    exp_54_ram[2417] = 0;
    exp_54_ram[2418] = 0;
    exp_54_ram[2419] = 0;
    exp_54_ram[2420] = 0;
    exp_54_ram[2421] = 153;
    exp_54_ram[2422] = 241;
    exp_54_ram[2423] = 49;
    exp_54_ram[2424] = 254;
    exp_54_ram[2425] = 0;
    exp_54_ram[2426] = 172;
    exp_54_ram[2427] = 0;
    exp_54_ram[2428] = 155;
    exp_54_ram[2429] = 0;
    exp_54_ram[2430] = 0;
    exp_54_ram[2431] = 0;
    exp_54_ram[2432] = 0;
    exp_54_ram[2433] = 154;
    exp_54_ram[2434] = 238;
    exp_54_ram[2435] = 46;
    exp_54_ram[2436] = 254;
    exp_54_ram[2437] = 0;
    exp_54_ram[2438] = 173;
    exp_54_ram[2439] = 0;
    exp_54_ram[2440] = 152;
    exp_54_ram[2441] = 0;
    exp_54_ram[2442] = 0;
    exp_54_ram[2443] = 0;
    exp_54_ram[2444] = 0;
    exp_54_ram[2445] = 154;
    exp_54_ram[2446] = 235;
    exp_54_ram[2447] = 43;
    exp_54_ram[2448] = 254;
    exp_54_ram[2449] = 0;
    exp_54_ram[2450] = 165;
    exp_54_ram[2451] = 0;
    exp_54_ram[2452] = 149;
    exp_54_ram[2453] = 0;
    exp_54_ram[2454] = 0;
    exp_54_ram[2455] = 0;
    exp_54_ram[2456] = 155;
    exp_54_ram[2457] = 232;
    exp_54_ram[2458] = 41;
    exp_54_ram[2459] = 254;
    exp_54_ram[2460] = 0;
    exp_54_ram[2461] = 173;
    exp_54_ram[2462] = 0;
    exp_54_ram[2463] = 146;
    exp_54_ram[2464] = 0;
    exp_54_ram[2465] = 0;
    exp_54_ram[2466] = 0;
    exp_54_ram[2467] = 0;
    exp_54_ram[2468] = 161;
    exp_54_ram[2469] = 229;
    exp_54_ram[2470] = 38;
    exp_54_ram[2471] = 0;
    exp_54_ram[2472] = 155;
    exp_54_ram[2473] = 228;
    exp_54_ram[2474] = 0;
    exp_54_ram[2475] = 174;
    exp_54_ram[2476] = 228;
    exp_54_ram[2477] = 254;
    exp_54_ram[2478] = 52;
    exp_54_ram[2479] = 35;
    exp_54_ram[2480] = 0;
    exp_54_ram[2481] = 0;
    exp_54_ram[2482] = 254;
    exp_54_ram[2483] = 0;
    exp_54_ram[2484] = 175;
    exp_54_ram[2485] = 0;
    exp_54_ram[2486] = 165;
    exp_54_ram[2487] = 0;
    exp_54_ram[2488] = 254;
    exp_54_ram[2489] = 0;
    exp_54_ram[2490] = 0;
    exp_54_ram[2491] = 153;
    exp_54_ram[2492] = 224;
    exp_54_ram[2493] = 32;
    exp_54_ram[2494] = 254;
    exp_54_ram[2495] = 0;
    exp_54_ram[2496] = 176;
    exp_54_ram[2497] = 0;
    exp_54_ram[2498] = 162;
    exp_54_ram[2499] = 0;
    exp_54_ram[2500] = 254;
    exp_54_ram[2501] = 64;
    exp_54_ram[2502] = 0;
    exp_54_ram[2503] = 0;
    exp_54_ram[2504] = 0;
    exp_54_ram[2505] = 154;
    exp_54_ram[2506] = 220;
    exp_54_ram[2507] = 28;
    exp_54_ram[2508] = 254;
    exp_54_ram[2509] = 0;
    exp_54_ram[2510] = 176;
    exp_54_ram[2511] = 0;
    exp_54_ram[2512] = 158;
    exp_54_ram[2513] = 0;
    exp_54_ram[2514] = 254;
    exp_54_ram[2515] = 64;
    exp_54_ram[2516] = 0;
    exp_54_ram[2517] = 0;
    exp_54_ram[2518] = 0;
    exp_54_ram[2519] = 154;
    exp_54_ram[2520] = 217;
    exp_54_ram[2521] = 25;
    exp_54_ram[2522] = 254;
    exp_54_ram[2523] = 3;
    exp_54_ram[2524] = 0;
    exp_54_ram[2525] = 248;
    exp_54_ram[2526] = 0;
    exp_54_ram[2527] = 254;
    exp_54_ram[2528] = 64;
    exp_54_ram[2529] = 0;
    exp_54_ram[2530] = 0;
    exp_54_ram[2531] = 0;
    exp_54_ram[2532] = 155;
    exp_54_ram[2533] = 213;
    exp_54_ram[2534] = 22;
    exp_54_ram[2535] = 254;
    exp_54_ram[2536] = 0;
    exp_54_ram[2537] = 173;
    exp_54_ram[2538] = 0;
    exp_54_ram[2539] = 152;
    exp_54_ram[2540] = 0;
    exp_54_ram[2541] = 0;
    exp_54_ram[2542] = 0;
    exp_54_ram[2543] = 161;
    exp_54_ram[2544] = 211;
    exp_54_ram[2545] = 19;
    exp_54_ram[2546] = 0;
    exp_54_ram[2547] = 155;
    exp_54_ram[2548] = 210;
    exp_54_ram[2549] = 0;
    exp_54_ram[2550] = 176;
    exp_54_ram[2551] = 209;
    exp_54_ram[2552] = 6;
    exp_54_ram[2553] = 254;
    exp_54_ram[2554] = 254;
    exp_54_ram[2555] = 0;
    exp_54_ram[2556] = 177;
    exp_54_ram[2557] = 0;
    exp_54_ram[2558] = 227;
    exp_54_ram[2559] = 0;
    exp_54_ram[2560] = 0;
    exp_54_ram[2561] = 0;
    exp_54_ram[2562] = 153;
    exp_54_ram[2563] = 206;
    exp_54_ram[2564] = 14;
    exp_54_ram[2565] = 254;
    exp_54_ram[2566] = 0;
    exp_54_ram[2567] = 6;
    exp_54_ram[2568] = 0;
    exp_54_ram[2569] = 233;
    exp_54_ram[2570] = 0;
    exp_54_ram[2571] = 0;
    exp_54_ram[2572] = 177;
    exp_54_ram[2573] = 0;
    exp_54_ram[2574] = 223;
    exp_54_ram[2575] = 0;
    exp_54_ram[2576] = 0;
    exp_54_ram[2577] = 0;
    exp_54_ram[2578] = 154;
    exp_54_ram[2579] = 202;
    exp_54_ram[2580] = 10;
    exp_54_ram[2581] = 254;
    exp_54_ram[2582] = 0;
    exp_54_ram[2583] = 6;
    exp_54_ram[2584] = 0;
    exp_54_ram[2585] = 229;
    exp_54_ram[2586] = 0;
    exp_54_ram[2587] = 0;
    exp_54_ram[2588] = 178;
    exp_54_ram[2589] = 0;
    exp_54_ram[2590] = 219;
    exp_54_ram[2591] = 0;
    exp_54_ram[2592] = 0;
    exp_54_ram[2593] = 0;
    exp_54_ram[2594] = 154;
    exp_54_ram[2595] = 198;
    exp_54_ram[2596] = 6;
    exp_54_ram[2597] = 254;
    exp_54_ram[2598] = 0;
    exp_54_ram[2599] = 6;
    exp_54_ram[2600] = 0;
    exp_54_ram[2601] = 225;
    exp_54_ram[2602] = 0;
    exp_54_ram[2603] = 0;
    exp_54_ram[2604] = 178;
    exp_54_ram[2605] = 0;
    exp_54_ram[2606] = 215;
    exp_54_ram[2607] = 0;
    exp_54_ram[2608] = 0;
    exp_54_ram[2609] = 0;
    exp_54_ram[2610] = 155;
    exp_54_ram[2611] = 194;
    exp_54_ram[2612] = 2;
    exp_54_ram[2613] = 0;
    exp_54_ram[2614] = 155;
    exp_54_ram[2615] = 193;
    exp_54_ram[2616] = 0;
    exp_54_ram[2617] = 179;
    exp_54_ram[2618] = 192;
    exp_54_ram[2619] = 0;
    exp_54_ram[2620] = 155;
    exp_54_ram[2621] = 191;
    exp_54_ram[2622] = 1;
    exp_54_ram[2623] = 1;
    exp_54_ram[2624] = 2;
    exp_54_ram[2625] = 0;
    exp_54_ram[2626] = 250;
    exp_54_ram[2627] = 4;
    exp_54_ram[2628] = 4;
    exp_54_ram[2629] = 5;
    exp_54_ram[2630] = 5;
    exp_54_ram[2631] = 5;
    exp_54_ram[2632] = 5;
    exp_54_ram[2633] = 5;
    exp_54_ram[2634] = 5;
    exp_54_ram[2635] = 6;
    exp_54_ram[2636] = 0;
    exp_54_ram[2637] = 180;
    exp_54_ram[2638] = 187;
    exp_54_ram[2639] = 7;
    exp_54_ram[2640] = 252;
    exp_54_ram[2641] = 0;
    exp_54_ram[2642] = 250;
    exp_54_ram[2643] = 1;
    exp_54_ram[2644] = 250;
    exp_54_ram[2645] = 0;
    exp_54_ram[2646] = 250;
    exp_54_ram[2647] = 1;
    exp_54_ram[2648] = 250;
    exp_54_ram[2649] = 250;
    exp_54_ram[2650] = 255;
    exp_54_ram[2651] = 252;
    exp_54_ram[2652] = 250;
    exp_54_ram[2653] = 0;
    exp_54_ram[2654] = 136;
    exp_54_ram[2655] = 0;
    exp_54_ram[2656] = 0;
    exp_54_ram[2657] = 250;
    exp_54_ram[2658] = 250;
    exp_54_ram[2659] = 250;
    exp_54_ram[2660] = 0;
    exp_54_ram[2661] = 180;
    exp_54_ram[2662] = 0;
    exp_54_ram[2663] = 0;
    exp_54_ram[2664] = 180;
    exp_54_ram[2665] = 0;
    exp_54_ram[2666] = 200;
    exp_54_ram[2667] = 0;
    exp_54_ram[2668] = 0;
    exp_54_ram[2669] = 0;
    exp_54_ram[2670] = 153;
    exp_54_ram[2671] = 179;
    exp_54_ram[2672] = 103;
    exp_54_ram[2673] = 250;
    exp_54_ram[2674] = 0;
    exp_54_ram[2675] = 157;
    exp_54_ram[2676] = 0;
    exp_54_ram[2677] = 0;
    exp_54_ram[2678] = 176;
    exp_54_ram[2679] = 0;
    exp_54_ram[2680] = 0;
    exp_54_ram[2681] = 182;
    exp_54_ram[2682] = 0;
    exp_54_ram[2683] = 195;
    exp_54_ram[2684] = 0;
    exp_54_ram[2685] = 0;
    exp_54_ram[2686] = 0;
    exp_54_ram[2687] = 154;
    exp_54_ram[2688] = 175;
    exp_54_ram[2689] = 98;
    exp_54_ram[2690] = 250;
    exp_54_ram[2691] = 0;
    exp_54_ram[2692] = 149;
    exp_54_ram[2693] = 0;
    exp_54_ram[2694] = 0;
    exp_54_ram[2695] = 172;
    exp_54_ram[2696] = 0;
    exp_54_ram[2697] = 0;
    exp_54_ram[2698] = 180;
    exp_54_ram[2699] = 0;
    exp_54_ram[2700] = 191;
    exp_54_ram[2701] = 0;
    exp_54_ram[2702] = 0;
    exp_54_ram[2703] = 0;
    exp_54_ram[2704] = 154;
    exp_54_ram[2705] = 170;
    exp_54_ram[2706] = 94;
    exp_54_ram[2707] = 250;
    exp_54_ram[2708] = 0;
    exp_54_ram[2709] = 158;
    exp_54_ram[2710] = 0;
    exp_54_ram[2711] = 0;
    exp_54_ram[2712] = 182;
    exp_54_ram[2713] = 0;
    exp_54_ram[2714] = 188;
    exp_54_ram[2715] = 0;
    exp_54_ram[2716] = 0;
    exp_54_ram[2717] = 0;
    exp_54_ram[2718] = 155;
    exp_54_ram[2719] = 167;
    exp_54_ram[2720] = 91;
    exp_54_ram[2721] = 7;
    exp_54_ram[2722] = 252;
    exp_54_ram[2723] = 0;
    exp_54_ram[2724] = 250;
    exp_54_ram[2725] = 1;
    exp_54_ram[2726] = 250;
    exp_54_ram[2727] = 0;
    exp_54_ram[2728] = 250;
    exp_54_ram[2729] = 1;
    exp_54_ram[2730] = 250;
    exp_54_ram[2731] = 250;
    exp_54_ram[2732] = 0;
    exp_54_ram[2733] = 252;
    exp_54_ram[2734] = 250;
    exp_54_ram[2735] = 0;
    exp_54_ram[2736] = 243;
    exp_54_ram[2737] = 0;
    exp_54_ram[2738] = 0;
    exp_54_ram[2739] = 250;
    exp_54_ram[2740] = 250;
    exp_54_ram[2741] = 250;
    exp_54_ram[2742] = 0;
    exp_54_ram[2743] = 160;
    exp_54_ram[2744] = 0;
    exp_54_ram[2745] = 0;
    exp_54_ram[2746] = 180;
    exp_54_ram[2747] = 0;
    exp_54_ram[2748] = 179;
    exp_54_ram[2749] = 0;
    exp_54_ram[2750] = 0;
    exp_54_ram[2751] = 0;
    exp_54_ram[2752] = 160;
    exp_54_ram[2753] = 158;
    exp_54_ram[2754] = 82;
    exp_54_ram[2755] = 250;
    exp_54_ram[2756] = 0;
    exp_54_ram[2757] = 137;
    exp_54_ram[2758] = 0;
    exp_54_ram[2759] = 0;
    exp_54_ram[2760] = 156;
    exp_54_ram[2761] = 0;
    exp_54_ram[2762] = 0;
    exp_54_ram[2763] = 182;
    exp_54_ram[2764] = 0;
    exp_54_ram[2765] = 175;
    exp_54_ram[2766] = 0;
    exp_54_ram[2767] = 0;
    exp_54_ram[2768] = 0;
    exp_54_ram[2769] = 161;
    exp_54_ram[2770] = 154;
    exp_54_ram[2771] = 78;
    exp_54_ram[2772] = 250;
    exp_54_ram[2773] = 0;
    exp_54_ram[2774] = 128;
    exp_54_ram[2775] = 0;
    exp_54_ram[2776] = 0;
    exp_54_ram[2777] = 151;
    exp_54_ram[2778] = 0;
    exp_54_ram[2779] = 0;
    exp_54_ram[2780] = 180;
    exp_54_ram[2781] = 0;
    exp_54_ram[2782] = 171;
    exp_54_ram[2783] = 0;
    exp_54_ram[2784] = 0;
    exp_54_ram[2785] = 0;
    exp_54_ram[2786] = 184;
    exp_54_ram[2787] = 150;
    exp_54_ram[2788] = 74;
    exp_54_ram[2789] = 250;
    exp_54_ram[2790] = 0;
    exp_54_ram[2791] = 138;
    exp_54_ram[2792] = 0;
    exp_54_ram[2793] = 0;
    exp_54_ram[2794] = 182;
    exp_54_ram[2795] = 0;
    exp_54_ram[2796] = 167;
    exp_54_ram[2797] = 0;
    exp_54_ram[2798] = 0;
    exp_54_ram[2799] = 0;
    exp_54_ram[2800] = 184;
    exp_54_ram[2801] = 146;
    exp_54_ram[2802] = 70;
    exp_54_ram[2803] = 7;
    exp_54_ram[2804] = 252;
    exp_54_ram[2805] = 0;
    exp_54_ram[2806] = 250;
    exp_54_ram[2807] = 1;
    exp_54_ram[2808] = 250;
    exp_54_ram[2809] = 0;
    exp_54_ram[2810] = 250;
    exp_54_ram[2811] = 1;
    exp_54_ram[2812] = 250;
    exp_54_ram[2813] = 250;
    exp_54_ram[2814] = 252;
    exp_54_ram[2815] = 250;
    exp_54_ram[2816] = 0;
    exp_54_ram[2817] = 223;
    exp_54_ram[2818] = 0;
    exp_54_ram[2819] = 0;
    exp_54_ram[2820] = 250;
    exp_54_ram[2821] = 250;
    exp_54_ram[2822] = 250;
    exp_54_ram[2823] = 0;
    exp_54_ram[2824] = 140;
    exp_54_ram[2825] = 0;
    exp_54_ram[2826] = 0;
    exp_54_ram[2827] = 182;
    exp_54_ram[2828] = 0;
    exp_54_ram[2829] = 159;
    exp_54_ram[2830] = 0;
    exp_54_ram[2831] = 0;
    exp_54_ram[2832] = 0;
    exp_54_ram[2833] = 185;
    exp_54_ram[2834] = 138;
    exp_54_ram[2835] = 62;
    exp_54_ram[2836] = 250;
    exp_54_ram[2837] = 0;
    exp_54_ram[2838] = 245;
    exp_54_ram[2839] = 0;
    exp_54_ram[2840] = 0;
    exp_54_ram[2841] = 135;
    exp_54_ram[2842] = 0;
    exp_54_ram[2843] = 0;
    exp_54_ram[2844] = 185;
    exp_54_ram[2845] = 0;
    exp_54_ram[2846] = 155;
    exp_54_ram[2847] = 0;
    exp_54_ram[2848] = 0;
    exp_54_ram[2849] = 0;
    exp_54_ram[2850] = 187;
    exp_54_ram[2851] = 134;
    exp_54_ram[2852] = 58;
    exp_54_ram[2853] = 250;
    exp_54_ram[2854] = 0;
    exp_54_ram[2855] = 236;
    exp_54_ram[2856] = 0;
    exp_54_ram[2857] = 0;
    exp_54_ram[2858] = 131;
    exp_54_ram[2859] = 0;
    exp_54_ram[2860] = 0;
    exp_54_ram[2861] = 182;
    exp_54_ram[2862] = 0;
    exp_54_ram[2863] = 150;
    exp_54_ram[2864] = 0;
    exp_54_ram[2865] = 0;
    exp_54_ram[2866] = 0;
    exp_54_ram[2867] = 187;
    exp_54_ram[2868] = 130;
    exp_54_ram[2869] = 53;
    exp_54_ram[2870] = 250;
    exp_54_ram[2871] = 0;
    exp_54_ram[2872] = 246;
    exp_54_ram[2873] = 0;
    exp_54_ram[2874] = 0;
    exp_54_ram[2875] = 185;
    exp_54_ram[2876] = 0;
    exp_54_ram[2877] = 147;
    exp_54_ram[2878] = 0;
    exp_54_ram[2879] = 0;
    exp_54_ram[2880] = 0;
    exp_54_ram[2881] = 188;
    exp_54_ram[2882] = 254;
    exp_54_ram[2883] = 50;
    exp_54_ram[2884] = 0;
    exp_54_ram[2885] = 155;
    exp_54_ram[2886] = 253;
    exp_54_ram[2887] = 7;
    exp_54_ram[2888] = 252;
    exp_54_ram[2889] = 0;
    exp_54_ram[2890] = 250;
    exp_54_ram[2891] = 1;
    exp_54_ram[2892] = 250;
    exp_54_ram[2893] = 250;
    exp_54_ram[2894] = 3;
    exp_54_ram[2895] = 250;
    exp_54_ram[2896] = 3;
    exp_54_ram[2897] = 250;
    exp_54_ram[2898] = 255;
    exp_54_ram[2899] = 252;
    exp_54_ram[2900] = 250;
    exp_54_ram[2901] = 0;
    exp_54_ram[2902] = 202;
    exp_54_ram[2903] = 0;
    exp_54_ram[2904] = 0;
    exp_54_ram[2905] = 250;
    exp_54_ram[2906] = 250;
    exp_54_ram[2907] = 250;
    exp_54_ram[2908] = 250;
    exp_54_ram[2909] = 0;
    exp_54_ram[2910] = 0;
    exp_54_ram[2911] = 239;
    exp_54_ram[2912] = 206;
    exp_54_ram[2913] = 252;
    exp_54_ram[2914] = 252;
    exp_54_ram[2915] = 252;
    exp_54_ram[2916] = 13;
    exp_54_ram[2917] = 0;
    exp_54_ram[2918] = 205;
    exp_54_ram[2919] = 0;
    exp_54_ram[2920] = 0;
    exp_54_ram[2921] = 253;
    exp_54_ram[2922] = 253;
    exp_54_ram[2923] = 0;
    exp_54_ram[2924] = 0;
    exp_54_ram[2925] = 205;
    exp_54_ram[2926] = 0;
    exp_54_ram[2927] = 0;
    exp_54_ram[2928] = 0;
    exp_54_ram[2929] = 12;
    exp_54_ram[2930] = 0;
    exp_54_ram[2931] = 253;
    exp_54_ram[2932] = 0;
    exp_54_ram[2933] = 0;
    exp_54_ram[2934] = 0;
    exp_54_ram[2935] = 0;
    exp_54_ram[2936] = 0;
    exp_54_ram[2937] = 0;
    exp_54_ram[2938] = 237;
    exp_54_ram[2939] = 0;
    exp_54_ram[2940] = 250;
    exp_54_ram[2941] = 0;
    exp_54_ram[2942] = 12;
    exp_54_ram[2943] = 0;
    exp_54_ram[2944] = 0;
    exp_54_ram[2945] = 253;
    exp_54_ram[2946] = 253;
    exp_54_ram[2947] = 1;
    exp_54_ram[2948] = 0;
    exp_54_ram[2949] = 0;
    exp_54_ram[2950] = 1;
    exp_54_ram[2951] = 0;
    exp_54_ram[2952] = 0;
    exp_54_ram[2953] = 252;
    exp_54_ram[2954] = 252;
    exp_54_ram[2955] = 0;
    exp_54_ram[2956] = 223;
    exp_54_ram[2957] = 0;
    exp_54_ram[2958] = 0;
    exp_54_ram[2959] = 250;
    exp_54_ram[2960] = 250;
    exp_54_ram[2961] = 250;
    exp_54_ram[2962] = 0;
    exp_54_ram[2963] = 223;
    exp_54_ram[2964] = 0;
    exp_54_ram[2965] = 0;
    exp_54_ram[2966] = 233;
    exp_54_ram[2967] = 253;
    exp_54_ram[2968] = 0;
    exp_54_ram[2969] = 252;
    exp_54_ram[2970] = 253;
    exp_54_ram[2971] = 0;
    exp_54_ram[2972] = 242;
    exp_54_ram[2973] = 7;
    exp_54_ram[2974] = 252;
    exp_54_ram[2975] = 0;
    exp_54_ram[2976] = 250;
    exp_54_ram[2977] = 1;
    exp_54_ram[2978] = 250;
    exp_54_ram[2979] = 0;
    exp_54_ram[2980] = 250;
    exp_54_ram[2981] = 3;
    exp_54_ram[2982] = 250;
    exp_54_ram[2983] = 3;
    exp_54_ram[2984] = 250;
    exp_54_ram[2985] = 0;
    exp_54_ram[2986] = 252;
    exp_54_ram[2987] = 250;
    exp_54_ram[2988] = 0;
    exp_54_ram[2989] = 180;
    exp_54_ram[2990] = 0;
    exp_54_ram[2991] = 0;
    exp_54_ram[2992] = 250;
    exp_54_ram[2993] = 250;
    exp_54_ram[2994] = 250;
    exp_54_ram[2995] = 0;
    exp_54_ram[2996] = 225;
    exp_54_ram[2997] = 0;
    exp_54_ram[2998] = 0;
    exp_54_ram[2999] = 225;
    exp_54_ram[3000] = 250;
    exp_54_ram[3001] = 0;
    exp_54_ram[3002] = 213;
    exp_54_ram[3003] = 0;
    exp_54_ram[3004] = 0;
    exp_54_ram[3005] = 223;
    exp_54_ram[3006] = 250;
    exp_54_ram[3007] = 250;
    exp_54_ram[3008] = 0;
    exp_54_ram[3009] = 0;
    exp_54_ram[3010] = 215;
    exp_54_ram[3011] = 0;
    exp_54_ram[3012] = 209;
    exp_54_ram[3013] = 0;
    exp_54_ram[3014] = 0;
    exp_54_ram[3015] = 250;
    exp_54_ram[3016] = 250;
    exp_54_ram[3017] = 250;
    exp_54_ram[3018] = 0;
    exp_54_ram[3019] = 209;
    exp_54_ram[3020] = 0;
    exp_54_ram[3021] = 0;
    exp_54_ram[3022] = 219;
    exp_54_ram[3023] = 179;
    exp_54_ram[3024] = 252;
    exp_54_ram[3025] = 252;
    exp_54_ram[3026] = 252;
    exp_54_ram[3027] = 13;
    exp_54_ram[3028] = 0;
    exp_54_ram[3029] = 177;
    exp_54_ram[3030] = 0;
    exp_54_ram[3031] = 0;
    exp_54_ram[3032] = 253;
    exp_54_ram[3033] = 253;
    exp_54_ram[3034] = 0;
    exp_54_ram[3035] = 0;
    exp_54_ram[3036] = 177;
    exp_54_ram[3037] = 0;
    exp_54_ram[3038] = 0;
    exp_54_ram[3039] = 0;
    exp_54_ram[3040] = 12;
    exp_54_ram[3041] = 0;
    exp_54_ram[3042] = 225;
    exp_54_ram[3043] = 0;
    exp_54_ram[3044] = 0;
    exp_54_ram[3045] = 0;
    exp_54_ram[3046] = 0;
    exp_54_ram[3047] = 0;
    exp_54_ram[3048] = 0;
    exp_54_ram[3049] = 209;
    exp_54_ram[3050] = 0;
    exp_54_ram[3051] = 250;
    exp_54_ram[3052] = 0;
    exp_54_ram[3053] = 12;
    exp_54_ram[3054] = 0;
    exp_54_ram[3055] = 0;
    exp_54_ram[3056] = 253;
    exp_54_ram[3057] = 253;
    exp_54_ram[3058] = 1;
    exp_54_ram[3059] = 0;
    exp_54_ram[3060] = 0;
    exp_54_ram[3061] = 1;
    exp_54_ram[3062] = 0;
    exp_54_ram[3063] = 0;
    exp_54_ram[3064] = 252;
    exp_54_ram[3065] = 252;
    exp_54_ram[3066] = 0;
    exp_54_ram[3067] = 195;
    exp_54_ram[3068] = 0;
    exp_54_ram[3069] = 0;
    exp_54_ram[3070] = 250;
    exp_54_ram[3071] = 250;
    exp_54_ram[3072] = 250;
    exp_54_ram[3073] = 0;
    exp_54_ram[3074] = 195;
    exp_54_ram[3075] = 0;
    exp_54_ram[3076] = 0;
    exp_54_ram[3077] = 205;
    exp_54_ram[3078] = 253;
    exp_54_ram[3079] = 0;
    exp_54_ram[3080] = 252;
    exp_54_ram[3081] = 253;
    exp_54_ram[3082] = 0;
    exp_54_ram[3083] = 242;
    exp_54_ram[3084] = 5;
    exp_54_ram[3085] = 5;
    exp_54_ram[3086] = 5;
    exp_54_ram[3087] = 5;
    exp_54_ram[3088] = 4;
    exp_54_ram[3089] = 4;
    exp_54_ram[3090] = 4;
    exp_54_ram[3091] = 4;
    exp_54_ram[3092] = 6;
    exp_54_ram[3093] = 0;
    exp_54_ram[3094] = 255;
    exp_54_ram[3095] = 0;
    exp_54_ram[3096] = 0;
    exp_54_ram[3097] = 1;
    exp_54_ram[3098] = 191;
    exp_54_ram[3099] = 137;
    exp_54_ram[3100] = 0;
    exp_54_ram[3101] = 0;
    exp_54_ram[3102] = 0;
    exp_54_ram[3103] = 1;
    exp_54_ram[3104] = 0;
    exp_54_ram[3105] = 0;
    exp_54_ram[3106] = 0;
    exp_54_ram[3107] = 2;
    exp_54_ram[3108] = 255;
    exp_54_ram[3109] = 2;
    exp_54_ram[3110] = 0;
    exp_54_ram[3111] = 0;
    exp_54_ram[3112] = 0;
    exp_54_ram[3113] = 64;
    exp_54_ram[3114] = 1;
    exp_54_ram[3115] = 0;
    exp_54_ram[3116] = 254;
    exp_54_ram[3117] = 255;
    exp_54_ram[3118] = 0;
    exp_54_ram[3119] = 254;
    exp_54_ram[3120] = 2;
    exp_54_ram[3121] = 128;
    exp_54_ram[3122] = 77;
    exp_54_ram[3123] = 117;
    exp_54_ram[3124] = 100;
    exp_54_ram[3125] = 70;
    exp_54_ram[3126] = 97;
    exp_54_ram[3127] = 0;
    exp_54_ram[3128] = 70;
    exp_54_ram[3129] = 97;
    exp_54_ram[3130] = 114;
    exp_54_ram[3131] = 74;
    exp_54_ram[3132] = 117;
    exp_54_ram[3133] = 103;
    exp_54_ram[3134] = 79;
    exp_54_ram[3135] = 111;
    exp_54_ram[3136] = 99;
    exp_54_ram[3137] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_252;
  assign exp_252 = exp_533;

  reg [3:0] exp_533_reg;
  always@(*) begin
    case (exp_385)
      0:exp_533_reg <= exp_520;
      1:exp_533_reg <= exp_525;
      2:exp_533_reg <= exp_526;
      3:exp_533_reg <= exp_527;
      4:exp_533_reg <= exp_528;
      5:exp_533_reg <= exp_529;
      6:exp_533_reg <= exp_530;
      7:exp_533_reg <= exp_531;
      default:exp_533_reg <= exp_532;
    endcase
  end
  assign exp_533 = exp_533_reg;
  assign exp_532 = 0;
  assign exp_520 = exp_516 << exp_519;
  assign exp_516 = 1;
  assign exp_519 = exp_518 + exp_517;
  assign exp_518 = 0;
  assign exp_517 = exp_453[1:0];
  assign exp_525 = exp_521 << exp_524;
  assign exp_521 = 3;
  assign exp_524 = exp_523 + exp_522;
  assign exp_523 = 0;
  assign exp_522 = exp_453[1:1];
  assign exp_526 = 15;
  assign exp_527 = 0;
  assign exp_528 = 0;
  assign exp_529 = 0;
  assign exp_530 = 0;
  assign exp_531 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_247;
  assign exp_247 = exp_515;

  reg [31:0] exp_515_reg;
  always@(*) begin
    case (exp_385)
      0:exp_515_reg <= exp_502;
      1:exp_515_reg <= exp_506;
      2:exp_515_reg <= exp_508;
      3:exp_515_reg <= exp_509;
      4:exp_515_reg <= exp_510;
      5:exp_515_reg <= exp_511;
      6:exp_515_reg <= exp_512;
      7:exp_515_reg <= exp_513;
      default:exp_515_reg <= exp_514;
    endcase
  end
  assign exp_515 = exp_515_reg;
  assign exp_514 = 0;

  reg [31:0] exp_502_reg;
  always@(*) begin
    case (exp_456)
      0:exp_502_reg <= exp_488;
      1:exp_502_reg <= exp_496;
      2:exp_502_reg <= exp_498;
      3:exp_502_reg <= exp_500;
      default:exp_502_reg <= exp_501;
    endcase
  end
  assign exp_502 = exp_502_reg;
  assign exp_501 = 0;
  assign exp_488 = exp_487;
  assign exp_487 = exp_486 + exp_485;
  assign exp_486 = 0;
  assign exp_485 = exp_375[7:0];

      reg [31:0] exp_375_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_375_reg <= exp_318;
        end
      end
      assign exp_375 = exp_375_reg;
      assign exp_496 = exp_488 << exp_495;
  assign exp_495 = 8;
  assign exp_498 = exp_488 << exp_497;
  assign exp_497 = 16;
  assign exp_500 = exp_488 << exp_499;
  assign exp_499 = 24;

  reg [31:0] exp_506_reg;
  always@(*) begin
    case (exp_459)
      0:exp_506_reg <= exp_492;
      1:exp_506_reg <= exp_504;
      default:exp_506_reg <= exp_505;
    endcase
  end
  assign exp_506 = exp_506_reg;
  assign exp_459 = exp_458 + exp_457;
  assign exp_458 = 0;
  assign exp_457 = exp_453[1:1];
  assign exp_505 = 0;
  assign exp_492 = exp_491;
  assign exp_491 = exp_490 + exp_489;
  assign exp_490 = 0;
  assign exp_489 = exp_375[15:0];
  assign exp_504 = exp_492 << exp_503;
  assign exp_503 = 16;
  assign exp_508 = exp_507 + exp_494;
  assign exp_507 = 0;
  assign exp_494 = exp_493 + exp_375;
  assign exp_493 = 0;
  assign exp_509 = 0;
  assign exp_510 = 0;
  assign exp_511 = 0;
  assign exp_512 = 0;
  assign exp_513 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 0;
    exp_47_ram[32] = 193;
    exp_47_ram[33] = 80;
    exp_47_ram[34] = 0;
    exp_47_ram[35] = 5;
    exp_47_ram[36] = 5;
    exp_47_ram[37] = 6;
    exp_47_ram[38] = 6;
    exp_47_ram[39] = 8;
    exp_47_ram[40] = 6;
    exp_47_ram[41] = 0;
    exp_47_ram[42] = 198;
    exp_47_ram[43] = 197;
    exp_47_ram[44] = 1;
    exp_47_ram[45] = 230;
    exp_47_ram[46] = 240;
    exp_47_ram[47] = 199;
    exp_47_ram[48] = 55;
    exp_47_ram[49] = 230;
    exp_47_ram[50] = 166;
    exp_47_ram[51] = 6;
    exp_47_ram[52] = 0;
    exp_47_ram[53] = 230;
    exp_47_ram[54] = 229;
    exp_47_ram[55] = 229;
    exp_47_ram[56] = 215;
    exp_47_ram[57] = 232;
    exp_47_ram[58] = 214;
    exp_47_ram[59] = 183;
    exp_47_ram[60] = 216;
    exp_47_ram[61] = 8;
    exp_47_ram[62] = 21;
    exp_47_ram[63] = 8;
    exp_47_ram[64] = 6;
    exp_47_ram[65] = 3;
    exp_47_ram[66] = 21;
    exp_47_ram[67] = 6;
    exp_47_ram[68] = 214;
    exp_47_ram[69] = 7;
    exp_47_ram[70] = 247;
    exp_47_ram[71] = 183;
    exp_47_ram[72] = 7;
    exp_47_ram[73] = 246;
    exp_47_ram[74] = 7;
    exp_47_ram[75] = 183;
    exp_47_ram[76] = 230;
    exp_47_ram[77] = 7;
    exp_47_ram[78] = 183;
    exp_47_ram[79] = 23;
    exp_47_ram[80] = 3;
    exp_47_ram[81] = 3;
    exp_47_ram[82] = 23;
    exp_47_ram[83] = 7;
    exp_47_ram[84] = 103;
    exp_47_ram[85] = 246;
    exp_47_ram[86] = 7;
    exp_47_ram[87] = 211;
    exp_47_ram[88] = 104;
    exp_47_ram[89] = 247;
    exp_47_ram[90] = 3;
    exp_47_ram[91] = 211;
    exp_47_ram[92] = 231;
    exp_47_ram[93] = 5;
    exp_47_ram[94] = 197;
    exp_47_ram[95] = 0;
    exp_47_ram[96] = 64;
    exp_47_ram[97] = 0;
    exp_47_ram[98] = 0;
    exp_47_ram[99] = 166;
    exp_47_ram[100] = 128;
    exp_47_ram[101] = 31;
    exp_47_ram[102] = 6;
    exp_47_ram[103] = 16;
    exp_47_ram[104] = 199;
    exp_47_ram[105] = 1;
    exp_47_ram[106] = 232;
    exp_47_ram[107] = 240;
    exp_47_ram[108] = 7;
    exp_47_ram[109] = 128;
    exp_47_ram[110] = 168;
    exp_47_ram[111] = 230;
    exp_47_ram[112] = 6;
    exp_47_ram[113] = 0;
    exp_47_ram[114] = 167;
    exp_47_ram[115] = 230;
    exp_47_ram[116] = 230;
    exp_47_ram[117] = 7;
    exp_47_ram[118] = 16;
    exp_47_ram[119] = 8;
    exp_47_ram[120] = 8;
    exp_47_ram[121] = 6;
    exp_47_ram[122] = 3;
    exp_47_ram[123] = 23;
    exp_47_ram[124] = 23;
    exp_47_ram[125] = 6;
    exp_47_ram[126] = 230;
    exp_47_ram[127] = 246;
    exp_47_ram[128] = 7;
    exp_47_ram[129] = 199;
    exp_47_ram[130] = 7;
    exp_47_ram[131] = 247;
    exp_47_ram[132] = 7;
    exp_47_ram[133] = 199;
    exp_47_ram[134] = 231;
    exp_47_ram[135] = 7;
    exp_47_ram[136] = 199;
    exp_47_ram[137] = 23;
    exp_47_ram[138] = 3;
    exp_47_ram[139] = 3;
    exp_47_ram[140] = 23;
    exp_47_ram[141] = 7;
    exp_47_ram[142] = 103;
    exp_47_ram[143] = 230;
    exp_47_ram[144] = 7;
    exp_47_ram[145] = 211;
    exp_47_ram[146] = 104;
    exp_47_ram[147] = 247;
    exp_47_ram[148] = 3;
    exp_47_ram[149] = 211;
    exp_47_ram[150] = 231;
    exp_47_ram[151] = 5;
    exp_47_ram[152] = 197;
    exp_47_ram[153] = 0;
    exp_47_ram[154] = 0;
    exp_47_ram[155] = 0;
    exp_47_ram[156] = 232;
    exp_47_ram[157] = 128;
    exp_47_ram[158] = 31;
    exp_47_ram[159] = 216;
    exp_47_ram[160] = 231;
    exp_47_ram[161] = 216;
    exp_47_ram[162] = 215;
    exp_47_ram[163] = 232;
    exp_47_ram[164] = 8;
    exp_47_ram[165] = 247;
    exp_47_ram[166] = 21;
    exp_47_ram[167] = 8;
    exp_47_ram[168] = 7;
    exp_47_ram[169] = 6;
    exp_47_ram[170] = 21;
    exp_47_ram[171] = 7;
    exp_47_ram[172] = 183;
    exp_47_ram[173] = 167;
    exp_47_ram[174] = 5;
    exp_47_ram[175] = 215;
    exp_47_ram[176] = 7;
    exp_47_ram[177] = 245;
    exp_47_ram[178] = 7;
    exp_47_ram[179] = 215;
    exp_47_ram[180] = 229;
    exp_47_ram[181] = 7;
    exp_47_ram[182] = 215;
    exp_47_ram[183] = 22;
    exp_47_ram[184] = 6;
    exp_47_ram[185] = 6;
    exp_47_ram[186] = 22;
    exp_47_ram[187] = 7;
    exp_47_ram[188] = 215;
    exp_47_ram[189] = 199;
    exp_47_ram[190] = 6;
    exp_47_ram[191] = 167;
    exp_47_ram[192] = 7;
    exp_47_ram[193] = 246;
    exp_47_ram[194] = 7;
    exp_47_ram[195] = 167;
    exp_47_ram[196] = 230;
    exp_47_ram[197] = 7;
    exp_47_ram[198] = 5;
    exp_47_ram[199] = 167;
    exp_47_ram[200] = 229;
    exp_47_ram[201] = 159;
    exp_47_ram[202] = 213;
    exp_47_ram[203] = 1;
    exp_47_ram[204] = 230;
    exp_47_ram[205] = 240;
    exp_47_ram[206] = 215;
    exp_47_ram[207] = 53;
    exp_47_ram[208] = 0;
    exp_47_ram[209] = 182;
    exp_47_ram[210] = 199;
    exp_47_ram[211] = 167;
    exp_47_ram[212] = 7;
    exp_47_ram[213] = 0;
    exp_47_ram[214] = 183;
    exp_47_ram[215] = 229;
    exp_47_ram[216] = 229;
    exp_47_ram[217] = 16;
    exp_47_ram[218] = 246;
    exp_47_ram[219] = 200;
    exp_47_ram[220] = 21;
    exp_47_ram[221] = 31;
    exp_47_ram[222] = 0;
    exp_47_ram[223] = 0;
    exp_47_ram[224] = 230;
    exp_47_ram[225] = 128;
    exp_47_ram[226] = 159;
    exp_47_ram[227] = 230;
    exp_47_ram[228] = 182;
    exp_47_ram[229] = 216;
    exp_47_ram[230] = 231;
    exp_47_ram[231] = 8;
    exp_47_ram[232] = 222;
    exp_47_ram[233] = 183;
    exp_47_ram[234] = 232;
    exp_47_ram[235] = 182;
    exp_47_ram[236] = 247;
    exp_47_ram[237] = 8;
    exp_47_ram[238] = 7;
    exp_47_ram[239] = 6;
    exp_47_ram[240] = 222;
    exp_47_ram[241] = 6;
    exp_47_ram[242] = 230;
    exp_47_ram[243] = 199;
    exp_47_ram[244] = 14;
    exp_47_ram[245] = 231;
    exp_47_ram[246] = 7;
    exp_47_ram[247] = 254;
    exp_47_ram[248] = 7;
    exp_47_ram[249] = 231;
    exp_47_ram[250] = 238;
    exp_47_ram[251] = 7;
    exp_47_ram[252] = 231;
    exp_47_ram[253] = 215;
    exp_47_ram[254] = 215;
    exp_47_ram[255] = 6;
    exp_47_ram[256] = 231;
    exp_47_ram[257] = 6;
    exp_47_ram[258] = 7;
    exp_47_ram[259] = 246;
    exp_47_ram[260] = 7;
    exp_47_ram[261] = 199;
    exp_47_ram[262] = 7;
    exp_47_ram[263] = 247;
    exp_47_ram[264] = 7;
    exp_47_ram[265] = 199;
    exp_47_ram[266] = 231;
    exp_47_ram[267] = 7;
    exp_47_ram[268] = 5;
    exp_47_ram[269] = 1;
    exp_47_ram[270] = 197;
    exp_47_ram[271] = 254;
    exp_47_ram[272] = 213;
    exp_47_ram[273] = 5;
    exp_47_ram[274] = 211;
    exp_47_ram[275] = 3;
    exp_47_ram[276] = 199;
    exp_47_ram[277] = 216;
    exp_47_ram[278] = 214;
    exp_47_ram[279] = 14;
    exp_47_ram[280] = 104;
    exp_47_ram[281] = 216;
    exp_47_ram[282] = 7;
    exp_47_ram[283] = 102;
    exp_47_ram[284] = 215;
    exp_47_ram[285] = 214;
    exp_47_ram[286] = 7;
    exp_47_ram[287] = 198;
    exp_47_ram[288] = 199;
    exp_47_ram[289] = 199;
    exp_47_ram[290] = 1;
    exp_47_ram[291] = 247;
    exp_47_ram[292] = 247;
    exp_47_ram[293] = 7;
    exp_47_ram[294] = 254;
    exp_47_ram[295] = 184;
    exp_47_ram[296] = 199;
    exp_47_ram[297] = 0;
    exp_47_ram[298] = 232;
    exp_47_ram[299] = 245;
    exp_47_ram[300] = 223;
    exp_47_ram[301] = 0;
    exp_47_ram[302] = 0;
    exp_47_ram[303] = 159;
    exp_47_ram[304] = 16;
    exp_47_ram[305] = 247;
    exp_47_ram[306] = 69;
    exp_47_ram[307] = 183;
    exp_47_ram[308] = 5;
    exp_47_ram[309] = 5;
    exp_47_ram[310] = 248;
    exp_47_ram[311] = 245;
    exp_47_ram[312] = 240;
    exp_47_ram[313] = 70;
    exp_47_ram[314] = 215;
    exp_47_ram[315] = 6;
    exp_47_ram[316] = 245;
    exp_47_ram[317] = 246;
    exp_47_ram[318] = 216;
    exp_47_ram[319] = 248;
    exp_47_ram[320] = 14;
    exp_47_ram[321] = 32;
    exp_47_ram[322] = 0;
    exp_47_ram[323] = 213;
    exp_47_ram[324] = 199;
    exp_47_ram[325] = 14;
    exp_47_ram[326] = 8;
    exp_47_ram[327] = 248;
    exp_47_ram[328] = 23;
    exp_47_ram[329] = 5;
    exp_47_ram[330] = 199;
    exp_47_ram[331] = 6;
    exp_47_ram[332] = 7;
    exp_47_ram[333] = 213;
    exp_47_ram[334] = 5;
    exp_47_ram[335] = 5;
    exp_47_ram[336] = 240;
    exp_47_ram[337] = 0;
    exp_47_ram[338] = 240;
    exp_47_ram[339] = 6;
    exp_47_ram[340] = 6;
    exp_47_ram[341] = 0;
    exp_47_ram[342] = 184;
    exp_47_ram[343] = 5;
    exp_47_ram[344] = 0;
    exp_47_ram[345] = 23;
    exp_47_ram[346] = 232;
    exp_47_ram[347] = 110;
    exp_47_ram[348] = 195;
    exp_47_ram[349] = 0;
    exp_47_ram[350] = 0;
    exp_47_ram[351] = 16;
    exp_47_ram[352] = 0;
    exp_47_ram[353] = 7;
    exp_47_ram[354] = 95;
    exp_47_ram[355] = 232;
    exp_47_ram[356] = 95;
    exp_47_ram[357] = 5;
    exp_47_ram[358] = 5;
    exp_47_ram[359] = 0;
    exp_47_ram[360] = 159;
    exp_47_ram[361] = 1;
    exp_47_ram[362] = 129;
    exp_47_ram[363] = 17;
    exp_47_ram[364] = 5;
    exp_47_ram[365] = 5;
    exp_47_ram[366] = 192;
    exp_47_ram[367] = 224;
    exp_47_ram[368] = 160;
    exp_47_ram[369] = 167;
    exp_47_ram[370] = 167;
    exp_47_ram[371] = 176;
    exp_47_ram[372] = 167;
    exp_47_ram[373] = 85;
    exp_47_ram[374] = 244;
    exp_47_ram[375] = 164;
    exp_47_ram[376] = 193;
    exp_47_ram[377] = 4;
    exp_47_ram[378] = 199;
    exp_47_ram[379] = 129;
    exp_47_ram[380] = 71;
    exp_47_ram[381] = 199;
    exp_47_ram[382] = 247;
    exp_47_ram[383] = 6;
    exp_47_ram[384] = 1;
    exp_47_ram[385] = 0;
    exp_47_ram[386] = 85;
    exp_47_ram[387] = 244;
    exp_47_ram[388] = 0;
    exp_47_ram[389] = 223;
    exp_47_ram[390] = 0;
    exp_47_ram[391] = 0;
    exp_47_ram[392] = 31;
    exp_47_ram[393] = 1;
    exp_47_ram[394] = 17;
    exp_47_ram[395] = 129;
    exp_47_ram[396] = 145;
    exp_47_ram[397] = 33;
    exp_47_ram[398] = 49;
    exp_47_ram[399] = 65;
    exp_47_ram[400] = 181;
    exp_47_ram[401] = 7;
    exp_47_ram[402] = 5;
    exp_47_ram[403] = 5;
    exp_47_ram[404] = 5;
    exp_47_ram[405] = 5;
    exp_47_ram[406] = 5;
    exp_47_ram[407] = 128;
    exp_47_ram[408] = 5;
    exp_47_ram[409] = 224;
    exp_47_ram[410] = 58;
    exp_47_ram[411] = 48;
    exp_47_ram[412] = 71;
    exp_47_ram[413] = 176;
    exp_47_ram[414] = 4;
    exp_47_ram[415] = 55;
    exp_47_ram[416] = 160;
    exp_47_ram[417] = 55;
    exp_47_ram[418] = 176;
    exp_47_ram[419] = 89;
    exp_47_ram[420] = 52;
    exp_47_ram[421] = 148;
    exp_47_ram[422] = 233;
    exp_47_ram[423] = 180;
    exp_47_ram[424] = 228;
    exp_47_ram[425] = 193;
    exp_47_ram[426] = 129;
    exp_47_ram[427] = 196;
    exp_47_ram[428] = 74;
    exp_47_ram[429] = 197;
    exp_47_ram[430] = 186;
    exp_47_ram[431] = 65;
    exp_47_ram[432] = 1;
    exp_47_ram[433] = 193;
    exp_47_ram[434] = 129;
    exp_47_ram[435] = 7;
    exp_47_ram[436] = 7;
    exp_47_ram[437] = 1;
    exp_47_ram[438] = 0;
    exp_47_ram[439] = 128;
    exp_47_ram[440] = 5;
    exp_47_ram[441] = 31;
    exp_47_ram[442] = 89;
    exp_47_ram[443] = 180;
    exp_47_ram[444] = 0;
    exp_47_ram[445] = 31;
    exp_47_ram[446] = 96;
    exp_47_ram[447] = 71;
    exp_47_ram[448] = 137;
    exp_47_ram[449] = 4;
    exp_47_ram[450] = 9;
    exp_47_ram[451] = 0;
    exp_47_ram[452] = 181;
    exp_47_ram[453] = 128;
    exp_47_ram[454] = 160;
    exp_47_ram[455] = 9;
    exp_47_ram[456] = 4;
    exp_47_ram[457] = 54;
    exp_47_ram[458] = 192;
    exp_47_ram[459] = 164;
    exp_47_ram[460] = 5;
    exp_47_ram[461] = 128;
    exp_47_ram[462] = 4;
    exp_47_ram[463] = 9;
    exp_47_ram[464] = 55;
    exp_47_ram[465] = 112;
    exp_47_ram[466] = 55;
    exp_47_ram[467] = 137;
    exp_47_ram[468] = 233;
    exp_47_ram[469] = 128;
    exp_47_ram[470] = 57;
    exp_47_ram[471] = 36;
    exp_47_ram[472] = 185;
    exp_47_ram[473] = 228;
    exp_47_ram[474] = 128;
    exp_47_ram[475] = 247;
    exp_47_ram[476] = 229;
    exp_47_ram[477] = 119;
    exp_47_ram[478] = 7;
    exp_47_ram[479] = 247;
    exp_47_ram[480] = 64;
    exp_47_ram[481] = 215;
    exp_47_ram[482] = 71;
    exp_47_ram[483] = 247;
    exp_47_ram[484] = 245;
    exp_47_ram[485] = 7;
    exp_47_ram[486] = 128;
    exp_47_ram[487] = 229;
    exp_47_ram[488] = 7;
    exp_47_ram[489] = 128;
    exp_47_ram[490] = 247;
    exp_47_ram[491] = 240;
    exp_47_ram[492] = 229;
    exp_47_ram[493] = 58;
    exp_47_ram[494] = 55;
    exp_47_ram[495] = 213;
    exp_47_ram[496] = 245;
    exp_47_ram[497] = 53;
    exp_47_ram[498] = 223;
    exp_47_ram[499] = 137;
    exp_47_ram[500] = 180;
    exp_47_ram[501] = 0;
    exp_47_ram[502] = 31;
    exp_47_ram[503] = 0;
    exp_47_ram[504] = 0;
    exp_47_ram[505] = 0;
    exp_47_ram[506] = 223;
    exp_47_ram[507] = 5;
    exp_47_ram[508] = 0;
    exp_47_ram[509] = 21;
    exp_47_ram[510] = 6;
    exp_47_ram[511] = 197;
    exp_47_ram[512] = 21;
    exp_47_ram[513] = 22;
    exp_47_ram[514] = 5;
    exp_47_ram[515] = 0;
    exp_47_ram[516] = 5;
    exp_47_ram[517] = 5;
    exp_47_ram[518] = 5;
    exp_47_ram[519] = 5;
    exp_47_ram[520] = 240;
    exp_47_ram[521] = 6;
    exp_47_ram[522] = 16;
    exp_47_ram[523] = 182;
    exp_47_ram[524] = 192;
    exp_47_ram[525] = 22;
    exp_47_ram[526] = 22;
    exp_47_ram[527] = 182;
    exp_47_ram[528] = 0;
    exp_47_ram[529] = 197;
    exp_47_ram[530] = 197;
    exp_47_ram[531] = 213;
    exp_47_ram[532] = 22;
    exp_47_ram[533] = 22;
    exp_47_ram[534] = 6;
    exp_47_ram[535] = 0;
    exp_47_ram[536] = 0;
    exp_47_ram[537] = 95;
    exp_47_ram[538] = 5;
    exp_47_ram[539] = 2;
    exp_47_ram[540] = 160;
    exp_47_ram[541] = 176;
    exp_47_ram[542] = 176;
    exp_47_ram[543] = 223;
    exp_47_ram[544] = 176;
    exp_47_ram[545] = 0;
    exp_47_ram[546] = 31;
    exp_47_ram[547] = 160;
    exp_47_ram[548] = 2;
    exp_47_ram[549] = 0;
    exp_47_ram[550] = 5;
    exp_47_ram[551] = 5;
    exp_47_ram[552] = 159;
    exp_47_ram[553] = 5;
    exp_47_ram[554] = 2;
    exp_47_ram[555] = 176;
    exp_47_ram[556] = 5;
    exp_47_ram[557] = 160;
    exp_47_ram[558] = 31;
    exp_47_ram[559] = 176;
    exp_47_ram[560] = 2;
    exp_47_ram[561] = 6;
    exp_47_ram[562] = 0;
    exp_47_ram[563] = 199;
    exp_47_ram[564] = 240;
    exp_47_ram[565] = 6;
    exp_47_ram[566] = 0;
    exp_47_ram[567] = 165;
    exp_47_ram[568] = 7;
    exp_47_ram[569] = 0;
    exp_47_ram[570] = 197;
    exp_47_ram[571] = 197;
    exp_47_ram[572] = 245;
    exp_47_ram[573] = 181;
    exp_47_ram[574] = 159;
    exp_47_ram[575] = 6;
    exp_47_ram[576] = 0;
    exp_47_ram[577] = 199;
    exp_47_ram[578] = 240;
    exp_47_ram[579] = 6;
    exp_47_ram[580] = 0;
    exp_47_ram[581] = 181;
    exp_47_ram[582] = 7;
    exp_47_ram[583] = 0;
    exp_47_ram[584] = 197;
    exp_47_ram[585] = 197;
    exp_47_ram[586] = 245;
    exp_47_ram[587] = 165;
    exp_47_ram[588] = 159;
    exp_47_ram[589] = 1;
    exp_47_ram[590] = 245;
    exp_47_ram[591] = 240;
    exp_47_ram[592] = 167;
    exp_47_ram[593] = 55;
    exp_47_ram[594] = 0;
    exp_47_ram[595] = 0;
    exp_47_ram[596] = 246;
    exp_47_ram[597] = 245;
    exp_47_ram[598] = 199;
    exp_47_ram[599] = 167;
    exp_47_ram[600] = 5;
    exp_47_ram[601] = 166;
    exp_47_ram[602] = 0;
    exp_47_ram[603] = 0;
    exp_47_ram[604] = 0;
    exp_47_ram[605] = 229;
    exp_47_ram[606] = 128;
    exp_47_ram[607] = 223;
    exp_47_ram[608] = 114;
    exp_47_ram[609] = 46;
    exp_47_ram[610] = 0;
    exp_47_ram[611] = 111;
    exp_47_ram[612] = 108;
    exp_47_ram[613] = 0;
    exp_47_ram[614] = 102;
    exp_47_ram[615] = 0;
    exp_47_ram[616] = 102;
    exp_47_ram[617] = 0;
    exp_47_ram[618] = 0;
    exp_47_ram[619] = 102;
    exp_47_ram[620] = 0;
    exp_47_ram[621] = 102;
    exp_47_ram[622] = 0;
    exp_47_ram[623] = 115;
    exp_47_ram[624] = 0;
    exp_47_ram[625] = 114;
    exp_47_ram[626] = 116;
    exp_47_ram[627] = 0;
    exp_47_ram[628] = 111;
    exp_47_ram[629] = 0;
    exp_47_ram[630] = 109;
    exp_47_ram[631] = 46;
    exp_47_ram[632] = 0;
    exp_47_ram[633] = 114;
    exp_47_ram[634] = 46;
    exp_47_ram[635] = 0;
    exp_47_ram[636] = 114;
    exp_47_ram[637] = 112;
    exp_47_ram[638] = 0;
    exp_47_ram[639] = 109;
    exp_47_ram[640] = 46;
    exp_47_ram[641] = 0;
    exp_47_ram[642] = 102;
    exp_47_ram[643] = 0;
    exp_47_ram[644] = 114;
    exp_47_ram[645] = 46;
    exp_47_ram[646] = 0;
    exp_47_ram[647] = 102;
    exp_47_ram[648] = 0;
    exp_47_ram[649] = 114;
    exp_47_ram[650] = 110;
    exp_47_ram[651] = 0;
    exp_47_ram[652] = 100;
    exp_47_ram[653] = 0;
    exp_47_ram[654] = 100;
    exp_47_ram[655] = 100;
    exp_47_ram[656] = 0;
    exp_47_ram[657] = 100;
    exp_47_ram[658] = 100;
    exp_47_ram[659] = 0;
    exp_47_ram[660] = 100;
    exp_47_ram[661] = 102;
    exp_47_ram[662] = 0;
    exp_47_ram[663] = 100;
    exp_47_ram[664] = 103;
    exp_47_ram[665] = 0;
    exp_47_ram[666] = 114;
    exp_47_ram[667] = 107;
    exp_47_ram[668] = 0;
    exp_47_ram[669] = 100;
    exp_47_ram[670] = 100;
    exp_47_ram[671] = 0;
    exp_47_ram[672] = 115;
    exp_47_ram[673] = 100;
    exp_47_ram[674] = 106;
    exp_47_ram[675] = 106;
    exp_47_ram[676] = 115;
    exp_47_ram[677] = 0;
    exp_47_ram[678] = 100;
    exp_47_ram[679] = 100;
    exp_47_ram[680] = 0;
    exp_47_ram[681] = 114;
    exp_47_ram[682] = 114;
    exp_47_ram[683] = 0;
    exp_47_ram[684] = 114;
    exp_47_ram[685] = 46;
    exp_47_ram[686] = 0;
    exp_47_ram[687] = 51;
    exp_47_ram[688] = 49;
    exp_47_ram[689] = 52;
    exp_47_ram[690] = 97;
    exp_47_ram[691] = 50;
    exp_47_ram[692] = 100;
    exp_47_ram[693] = 115;
    exp_47_ram[694] = 51;
    exp_47_ram[695] = 49;
    exp_47_ram[696] = 97;
    exp_47_ram[697] = 103;
    exp_47_ram[698] = 0;
    exp_47_ram[699] = 114;
    exp_47_ram[700] = 46;
    exp_47_ram[701] = 0;
    exp_47_ram[702] = 51;
    exp_47_ram[703] = 0;
    exp_47_ram[704] = 52;
    exp_47_ram[705] = 0;
    exp_47_ram[706] = 109;
    exp_47_ram[707] = 46;
    exp_47_ram[708] = 0;
    exp_47_ram[709] = 51;
    exp_47_ram[710] = 0;
    exp_47_ram[711] = 51;
    exp_47_ram[712] = 0;
    exp_47_ram[713] = 99;
    exp_47_ram[714] = 0;
    exp_47_ram[715] = 100;
    exp_47_ram[716] = 0;
    exp_47_ram[717] = 114;
    exp_47_ram[718] = 46;
    exp_47_ram[719] = 0;
    exp_47_ram[720] = 109;
    exp_47_ram[721] = 46;
    exp_47_ram[722] = 117;
    exp_47_ram[723] = 112;
    exp_47_ram[724] = 32;
    exp_47_ram[725] = 50;
    exp_47_ram[726] = 48;
    exp_47_ram[727] = 50;
    exp_47_ram[728] = 0;
    exp_47_ram[729] = 117;
    exp_47_ram[730] = 112;
    exp_47_ram[731] = 32;
    exp_47_ram[732] = 50;
    exp_47_ram[733] = 48;
    exp_47_ram[734] = 50;
    exp_47_ram[735] = 0;
    exp_47_ram[736] = 102;
    exp_47_ram[737] = 0;
    exp_47_ram[738] = 102;
    exp_47_ram[739] = 0;
    exp_47_ram[740] = 102;
    exp_47_ram[741] = 0;
    exp_47_ram[742] = 117;
    exp_47_ram[743] = 112;
    exp_47_ram[744] = 32;
    exp_47_ram[745] = 50;
    exp_47_ram[746] = 48;
    exp_47_ram[747] = 50;
    exp_47_ram[748] = 0;
    exp_47_ram[749] = 32;
    exp_47_ram[750] = 108;
    exp_47_ram[751] = 32;
    exp_47_ram[752] = 108;
    exp_47_ram[753] = 32;
    exp_47_ram[754] = 108;
    exp_47_ram[755] = 2;
    exp_47_ram[756] = 3;
    exp_47_ram[757] = 4;
    exp_47_ram[758] = 4;
    exp_47_ram[759] = 5;
    exp_47_ram[760] = 5;
    exp_47_ram[761] = 5;
    exp_47_ram[762] = 5;
    exp_47_ram[763] = 6;
    exp_47_ram[764] = 6;
    exp_47_ram[765] = 6;
    exp_47_ram[766] = 6;
    exp_47_ram[767] = 6;
    exp_47_ram[768] = 6;
    exp_47_ram[769] = 6;
    exp_47_ram[770] = 6;
    exp_47_ram[771] = 7;
    exp_47_ram[772] = 7;
    exp_47_ram[773] = 7;
    exp_47_ram[774] = 7;
    exp_47_ram[775] = 7;
    exp_47_ram[776] = 7;
    exp_47_ram[777] = 7;
    exp_47_ram[778] = 7;
    exp_47_ram[779] = 7;
    exp_47_ram[780] = 7;
    exp_47_ram[781] = 7;
    exp_47_ram[782] = 7;
    exp_47_ram[783] = 7;
    exp_47_ram[784] = 7;
    exp_47_ram[785] = 7;
    exp_47_ram[786] = 7;
    exp_47_ram[787] = 8;
    exp_47_ram[788] = 8;
    exp_47_ram[789] = 8;
    exp_47_ram[790] = 8;
    exp_47_ram[791] = 8;
    exp_47_ram[792] = 8;
    exp_47_ram[793] = 8;
    exp_47_ram[794] = 8;
    exp_47_ram[795] = 8;
    exp_47_ram[796] = 8;
    exp_47_ram[797] = 8;
    exp_47_ram[798] = 8;
    exp_47_ram[799] = 8;
    exp_47_ram[800] = 8;
    exp_47_ram[801] = 8;
    exp_47_ram[802] = 8;
    exp_47_ram[803] = 8;
    exp_47_ram[804] = 8;
    exp_47_ram[805] = 8;
    exp_47_ram[806] = 8;
    exp_47_ram[807] = 8;
    exp_47_ram[808] = 8;
    exp_47_ram[809] = 8;
    exp_47_ram[810] = 8;
    exp_47_ram[811] = 8;
    exp_47_ram[812] = 8;
    exp_47_ram[813] = 8;
    exp_47_ram[814] = 8;
    exp_47_ram[815] = 8;
    exp_47_ram[816] = 8;
    exp_47_ram[817] = 8;
    exp_47_ram[818] = 8;
    exp_47_ram[819] = 5;
    exp_47_ram[820] = 0;
    exp_47_ram[821] = 167;
    exp_47_ram[822] = 7;
    exp_47_ram[823] = 7;
    exp_47_ram[824] = 0;
    exp_47_ram[825] = 21;
    exp_47_ram[826] = 229;
    exp_47_ram[827] = 159;
    exp_47_ram[828] = 1;
    exp_47_ram[829] = 0;
    exp_47_ram[830] = 129;
    exp_47_ram[831] = 71;
    exp_47_ram[832] = 17;
    exp_47_ram[833] = 4;
    exp_47_ram[834] = 95;
    exp_47_ram[835] = 160;
    exp_47_ram[836] = 193;
    exp_47_ram[837] = 244;
    exp_47_ram[838] = 129;
    exp_47_ram[839] = 0;
    exp_47_ram[840] = 1;
    exp_47_ram[841] = 0;
    exp_47_ram[842] = 181;
    exp_47_ram[843] = 55;
    exp_47_ram[844] = 5;
    exp_47_ram[845] = 7;
    exp_47_ram[846] = 5;
    exp_47_ram[847] = 197;
    exp_47_ram[848] = 240;
    exp_47_ram[849] = 192;
    exp_47_ram[850] = 7;
    exp_47_ram[851] = 7;
    exp_47_ram[852] = 6;
    exp_47_ram[853] = 22;
    exp_47_ram[854] = 71;
    exp_47_ram[855] = 22;
    exp_47_ram[856] = 135;
    exp_47_ram[857] = 22;
    exp_47_ram[858] = 199;
    exp_47_ram[859] = 22;
    exp_47_ram[860] = 227;
    exp_47_ram[861] = 24;
    exp_47_ram[862] = 246;
    exp_47_ram[863] = 6;
    exp_47_ram[864] = 197;
    exp_47_ram[865] = 197;
    exp_47_ram[866] = 48;
    exp_47_ram[867] = 247;
    exp_47_ram[868] = 6;
    exp_47_ram[869] = 55;
    exp_47_ram[870] = 199;
    exp_47_ram[871] = 230;
    exp_47_ram[872] = 229;
    exp_47_ram[873] = 0;
    exp_47_ram[874] = 246;
    exp_47_ram[875] = 0;
    exp_47_ram[876] = 245;
    exp_47_ram[877] = 8;
    exp_47_ram[878] = 246;
    exp_47_ram[879] = 71;
    exp_47_ram[880] = 24;
    exp_47_ram[881] = 159;
    exp_47_ram[882] = 245;
    exp_47_ram[883] = 7;
    exp_47_ram[884] = 246;
    exp_47_ram[885] = 23;
    exp_47_ram[886] = 7;
    exp_47_ram[887] = 223;
    exp_47_ram[888] = 5;
    exp_47_ram[889] = 7;
    exp_47_ram[890] = 7;
    exp_47_ram[891] = 199;
    exp_47_ram[892] = 5;
    exp_47_ram[893] = 7;
    exp_47_ram[894] = 247;
    exp_47_ram[895] = 7;
    exp_47_ram[896] = 0;
    exp_47_ram[897] = 23;
    exp_47_ram[898] = 223;
    exp_47_ram[899] = 199;
    exp_47_ram[900] = 23;
    exp_47_ram[901] = 21;
    exp_47_ram[902] = 231;
    exp_47_ram[903] = 95;
    exp_47_ram[904] = 7;
    exp_47_ram[905] = 0;
    exp_47_ram[906] = 181;
    exp_47_ram[907] = 55;
    exp_47_ram[908] = 7;
    exp_47_ram[909] = 255;
    exp_47_ram[910] = 128;
    exp_47_ram[911] = 246;
    exp_47_ram[912] = 6;
    exp_47_ram[913] = 5;
    exp_47_ram[914] = 5;
    exp_47_ram[915] = 231;
    exp_47_ram[916] = 5;
    exp_47_ram[917] = 5;
    exp_47_ram[918] = 7;
    exp_47_ram[919] = 231;
    exp_47_ram[920] = 231;
    exp_47_ram[921] = 0;
    exp_47_ram[922] = 215;
    exp_47_ram[923] = 247;
    exp_47_ram[924] = 247;
    exp_47_ram[925] = 199;
    exp_47_ram[926] = 7;
    exp_47_ram[927] = 69;
    exp_47_ram[928] = 69;
    exp_47_ram[929] = 31;
    exp_47_ram[930] = 21;
    exp_47_ram[931] = 21;
    exp_47_ram[932] = 31;
    exp_47_ram[933] = 0;
    exp_47_ram[934] = 0;
    exp_47_ram[935] = 5;
    exp_47_ram[936] = 0;
    exp_47_ram[937] = 167;
    exp_47_ram[938] = 7;
    exp_47_ram[939] = 7;
    exp_47_ram[940] = 0;
    exp_47_ram[941] = 21;
    exp_47_ram[942] = 223;
    exp_47_ram[943] = 0;
    exp_47_ram[944] = 199;
    exp_47_ram[945] = 0;
    exp_47_ram[946] = 245;
    exp_47_ram[947] = 183;
    exp_47_ram[948] = 23;
    exp_47_ram[949] = 223;
    exp_47_ram[950] = 5;
    exp_47_ram[951] = 197;
    exp_47_ram[952] = 199;
    exp_47_ram[953] = 0;
    exp_47_ram[954] = 64;
    exp_47_ram[955] = 7;
    exp_47_ram[956] = 5;
    exp_47_ram[957] = 23;
    exp_47_ram[958] = 183;
    exp_47_ram[959] = 0;
    exp_47_ram[960] = 1;
    exp_47_ram[961] = 129;
    exp_47_ram[962] = 145;
    exp_47_ram[963] = 5;
    exp_47_ram[964] = 17;
    exp_47_ram[965] = 5;
    exp_47_ram[966] = 95;
    exp_47_ram[967] = 4;
    exp_47_ram[968] = 164;
    exp_47_ram[969] = 231;
    exp_47_ram[970] = 0;
    exp_47_ram[971] = 64;
    exp_47_ram[972] = 7;
    exp_47_ram[973] = 5;
    exp_47_ram[974] = 23;
    exp_47_ram[975] = 150;
    exp_47_ram[976] = 193;
    exp_47_ram[977] = 129;
    exp_47_ram[978] = 65;
    exp_47_ram[979] = 1;
    exp_47_ram[980] = 0;
    exp_47_ram[981] = 1;
    exp_47_ram[982] = 129;
    exp_47_ram[983] = 145;
    exp_47_ram[984] = 5;
    exp_47_ram[985] = 17;
    exp_47_ram[986] = 5;
    exp_47_ram[987] = 31;
    exp_47_ram[988] = 245;
    exp_47_ram[989] = 244;
    exp_47_ram[990] = 244;
    exp_47_ram[991] = 0;
    exp_47_ram[992] = 64;
    exp_47_ram[993] = 7;
    exp_47_ram[994] = 5;
    exp_47_ram[995] = 247;
    exp_47_ram[996] = 151;
    exp_47_ram[997] = 193;
    exp_47_ram[998] = 129;
    exp_47_ram[999] = 65;
    exp_47_ram[1000] = 1;
    exp_47_ram[1001] = 0;
    exp_47_ram[1002] = 1;
    exp_47_ram[1003] = 129;
    exp_47_ram[1004] = 145;
    exp_47_ram[1005] = 33;
    exp_47_ram[1006] = 49;
    exp_47_ram[1007] = 17;
    exp_47_ram[1008] = 5;
    exp_47_ram[1009] = 5;
    exp_47_ram[1010] = 95;
    exp_47_ram[1011] = 5;
    exp_47_ram[1012] = 0;
    exp_47_ram[1013] = 137;
    exp_47_ram[1014] = 4;
    exp_47_ram[1015] = 31;
    exp_47_ram[1016] = 0;
    exp_47_ram[1017] = 137;
    exp_47_ram[1018] = 128;
    exp_47_ram[1019] = 244;
    exp_47_ram[1020] = 6;
    exp_47_ram[1021] = 7;
    exp_47_ram[1022] = 230;
    exp_47_ram[1023] = 23;
    exp_47_ram[1024] = 245;
    exp_47_ram[1025] = 193;
    exp_47_ram[1026] = 4;
    exp_47_ram[1027] = 129;
    exp_47_ram[1028] = 65;
    exp_47_ram[1029] = 1;
    exp_47_ram[1030] = 193;
    exp_47_ram[1031] = 1;
    exp_47_ram[1032] = 0;
    exp_47_ram[1033] = 20;
    exp_47_ram[1034] = 223;
    exp_47_ram[1035] = 1;
    exp_47_ram[1036] = 129;
    exp_47_ram[1037] = 145;
    exp_47_ram[1038] = 33;
    exp_47_ram[1039] = 49;
    exp_47_ram[1040] = 17;
    exp_47_ram[1041] = 5;
    exp_47_ram[1042] = 5;
    exp_47_ram[1043] = 31;
    exp_47_ram[1044] = 5;
    exp_47_ram[1045] = 0;
    exp_47_ram[1046] = 137;
    exp_47_ram[1047] = 4;
    exp_47_ram[1048] = 223;
    exp_47_ram[1049] = 0;
    exp_47_ram[1050] = 137;
    exp_47_ram[1051] = 128;
    exp_47_ram[1052] = 244;
    exp_47_ram[1053] = 6;
    exp_47_ram[1054] = 7;
    exp_47_ram[1055] = 230;
    exp_47_ram[1056] = 23;
    exp_47_ram[1057] = 245;
    exp_47_ram[1058] = 20;
    exp_47_ram[1059] = 223;
    exp_47_ram[1060] = 193;
    exp_47_ram[1061] = 4;
    exp_47_ram[1062] = 129;
    exp_47_ram[1063] = 65;
    exp_47_ram[1064] = 1;
    exp_47_ram[1065] = 193;
    exp_47_ram[1066] = 1;
    exp_47_ram[1067] = 0;
    exp_47_ram[1068] = 1;
    exp_47_ram[1069] = 129;
    exp_47_ram[1070] = 145;
    exp_47_ram[1071] = 33;
    exp_47_ram[1072] = 5;
    exp_47_ram[1073] = 17;
    exp_47_ram[1074] = 5;
    exp_47_ram[1075] = 31;
    exp_47_ram[1076] = 164;
    exp_47_ram[1077] = 36;
    exp_47_ram[1078] = 4;
    exp_47_ram[1079] = 31;
    exp_47_ram[1080] = 5;
    exp_47_ram[1081] = 0;
    exp_47_ram[1082] = 192;
    exp_47_ram[1083] = 244;
    exp_47_ram[1084] = 4;
    exp_47_ram[1085] = 6;
    exp_47_ram[1086] = 4;
    exp_47_ram[1087] = 214;
    exp_47_ram[1088] = 23;
    exp_47_ram[1089] = 247;
    exp_47_ram[1090] = 20;
    exp_47_ram[1091] = 159;
    exp_47_ram[1092] = 0;
    exp_47_ram[1093] = 193;
    exp_47_ram[1094] = 129;
    exp_47_ram[1095] = 65;
    exp_47_ram[1096] = 1;
    exp_47_ram[1097] = 1;
    exp_47_ram[1098] = 0;
    exp_47_ram[1099] = 1;
    exp_47_ram[1100] = 129;
    exp_47_ram[1101] = 145;
    exp_47_ram[1102] = 33;
    exp_47_ram[1103] = 49;
    exp_47_ram[1104] = 17;
    exp_47_ram[1105] = 5;
    exp_47_ram[1106] = 5;
    exp_47_ram[1107] = 31;
    exp_47_ram[1108] = 5;
    exp_47_ram[1109] = 0;
    exp_47_ram[1110] = 137;
    exp_47_ram[1111] = 4;
    exp_47_ram[1112] = 223;
    exp_47_ram[1113] = 5;
    exp_47_ram[1114] = 0;
    exp_47_ram[1115] = 137;
    exp_47_ram[1116] = 192;
    exp_47_ram[1117] = 245;
    exp_47_ram[1118] = 244;
    exp_47_ram[1119] = 6;
    exp_47_ram[1120] = 6;
    exp_47_ram[1121] = 214;
    exp_47_ram[1122] = 23;
    exp_47_ram[1123] = 247;
    exp_47_ram[1124] = 193;
    exp_47_ram[1125] = 129;
    exp_47_ram[1126] = 65;
    exp_47_ram[1127] = 1;
    exp_47_ram[1128] = 193;
    exp_47_ram[1129] = 1;
    exp_47_ram[1130] = 0;
    exp_47_ram[1131] = 0;
    exp_47_ram[1132] = 31;
    exp_47_ram[1133] = 20;
    exp_47_ram[1134] = 31;
    exp_47_ram[1135] = 53;
    exp_47_ram[1136] = 7;
    exp_47_ram[1137] = 1;
    exp_47_ram[1138] = 64;
    exp_47_ram[1139] = 129;
    exp_47_ram[1140] = 17;
    exp_47_ram[1141] = 5;
    exp_47_ram[1142] = 143;
    exp_47_ram[1143] = 16;
    exp_47_ram[1144] = 5;
    exp_47_ram[1145] = 0;
    exp_47_ram[1146] = 4;
    exp_47_ram[1147] = 79;
    exp_47_ram[1148] = 21;
    exp_47_ram[1149] = 193;
    exp_47_ram[1150] = 129;
    exp_47_ram[1151] = 7;
    exp_47_ram[1152] = 1;
    exp_47_ram[1153] = 0;
    exp_47_ram[1154] = 0;
    exp_47_ram[1155] = 7;
    exp_47_ram[1156] = 0;
    exp_47_ram[1157] = 213;
    exp_47_ram[1158] = 215;
    exp_47_ram[1159] = 7;
    exp_47_ram[1160] = 213;
    exp_47_ram[1161] = 128;
    exp_47_ram[1162] = 224;
    exp_47_ram[1163] = 215;
    exp_47_ram[1164] = 16;
    exp_47_ram[1165] = 240;
    exp_47_ram[1166] = 229;
    exp_47_ram[1167] = 1;
    exp_47_ram[1168] = 17;
    exp_47_ram[1169] = 159;
    exp_47_ram[1170] = 193;
    exp_47_ram[1171] = 160;
    exp_47_ram[1172] = 199;
    exp_47_ram[1173] = 7;
    exp_47_ram[1174] = 1;
    exp_47_ram[1175] = 0;
    exp_47_ram[1176] = 224;
    exp_47_ram[1177] = 7;
    exp_47_ram[1178] = 0;
    exp_47_ram[1179] = 0;
    exp_47_ram[1180] = 7;
    exp_47_ram[1181] = 71;
    exp_47_ram[1182] = 71;
    exp_47_ram[1183] = 6;
    exp_47_ram[1184] = 135;
    exp_47_ram[1185] = 213;
    exp_47_ram[1186] = 0;
    exp_47_ram[1187] = 5;
    exp_47_ram[1188] = 197;
    exp_47_ram[1189] = 167;
    exp_47_ram[1190] = 213;
    exp_47_ram[1191] = 1;
    exp_47_ram[1192] = 245;
    exp_47_ram[1193] = 17;
    exp_47_ram[1194] = 207;
    exp_47_ram[1195] = 193;
    exp_47_ram[1196] = 1;
    exp_47_ram[1197] = 0;
    exp_47_ram[1198] = 1;
    exp_47_ram[1199] = 81;
    exp_47_ram[1200] = 69;
    exp_47_ram[1201] = 145;
    exp_47_ram[1202] = 1;
    exp_47_ram[1203] = 129;
    exp_47_ram[1204] = 33;
    exp_47_ram[1205] = 49;
    exp_47_ram[1206] = 65;
    exp_47_ram[1207] = 17;
    exp_47_ram[1208] = 97;
    exp_47_ram[1209] = 5;
    exp_47_ram[1210] = 32;
    exp_47_ram[1211] = 0;
    exp_47_ram[1212] = 0;
    exp_47_ram[1213] = 202;
    exp_47_ram[1214] = 4;
    exp_47_ram[1215] = 138;
    exp_47_ram[1216] = 10;
    exp_47_ram[1217] = 1;
    exp_47_ram[1218] = 0;
    exp_47_ram[1219] = 10;
    exp_47_ram[1220] = 155;
    exp_47_ram[1221] = 4;
    exp_47_ram[1222] = 4;
    exp_47_ram[1223] = 159;
    exp_47_ram[1224] = 10;
    exp_47_ram[1225] = 143;
    exp_47_ram[1226] = 169;
    exp_47_ram[1227] = 37;
    exp_47_ram[1228] = 55;
    exp_47_ram[1229] = 5;
    exp_47_ram[1230] = 20;
    exp_47_ram[1231] = 95;
    exp_47_ram[1232] = 4;
    exp_47_ram[1233] = 159;
    exp_47_ram[1234] = 160;
    exp_47_ram[1235] = 4;
    exp_47_ram[1236] = 213;
    exp_47_ram[1237] = 143;
    exp_47_ram[1238] = 169;
    exp_47_ram[1239] = 37;
    exp_47_ram[1240] = 55;
    exp_47_ram[1241] = 5;
    exp_47_ram[1242] = 20;
    exp_47_ram[1243] = 31;
    exp_47_ram[1244] = 138;
    exp_47_ram[1245] = 74;
    exp_47_ram[1246] = 10;
    exp_47_ram[1247] = 55;
    exp_47_ram[1248] = 231;
    exp_47_ram[1249] = 87;
    exp_47_ram[1250] = 231;
    exp_47_ram[1251] = 70;
    exp_47_ram[1252] = 199;
    exp_47_ram[1253] = 71;
    exp_47_ram[1254] = 39;
    exp_47_ram[1255] = 202;
    exp_47_ram[1256] = 247;
    exp_47_ram[1257] = 247;
    exp_47_ram[1258] = 231;
    exp_47_ram[1259] = 198;
    exp_47_ram[1260] = 247;
    exp_47_ram[1261] = 215;
    exp_47_ram[1262] = 1;
    exp_47_ram[1263] = 244;
    exp_47_ram[1264] = 151;
    exp_47_ram[1265] = 228;
    exp_47_ram[1266] = 215;
    exp_47_ram[1267] = 5;
    exp_47_ram[1268] = 245;
    exp_47_ram[1269] = 247;
    exp_47_ram[1270] = 79;
    exp_47_ram[1271] = 164;
    exp_47_ram[1272] = 245;
    exp_47_ram[1273] = 149;
    exp_47_ram[1274] = 244;
    exp_47_ram[1275] = 37;
    exp_47_ram[1276] = 244;
    exp_47_ram[1277] = 52;
    exp_47_ram[1278] = 181;
    exp_47_ram[1279] = 193;
    exp_47_ram[1280] = 133;
    exp_47_ram[1281] = 129;
    exp_47_ram[1282] = 65;
    exp_47_ram[1283] = 1;
    exp_47_ram[1284] = 193;
    exp_47_ram[1285] = 129;
    exp_47_ram[1286] = 65;
    exp_47_ram[1287] = 1;
    exp_47_ram[1288] = 1;
    exp_47_ram[1289] = 0;
    exp_47_ram[1290] = 1;
    exp_47_ram[1291] = 17;
    exp_47_ram[1292] = 129;
    exp_47_ram[1293] = 5;
    exp_47_ram[1294] = 95;
    exp_47_ram[1295] = 0;
    exp_47_ram[1296] = 7;
    exp_47_ram[1297] = 0;
    exp_47_ram[1298] = 95;
    exp_47_ram[1299] = 0;
    exp_47_ram[1300] = 135;
    exp_47_ram[1301] = 245;
    exp_47_ram[1302] = 4;
    exp_47_ram[1303] = 164;
    exp_47_ram[1304] = 4;
    exp_47_ram[1305] = 193;
    exp_47_ram[1306] = 129;
    exp_47_ram[1307] = 0;
    exp_47_ram[1308] = 1;
    exp_47_ram[1309] = 0;
    exp_47_ram[1310] = 1;
    exp_47_ram[1311] = 17;
    exp_47_ram[1312] = 129;
    exp_47_ram[1313] = 145;
    exp_47_ram[1314] = 33;
    exp_47_ram[1315] = 5;
    exp_47_ram[1316] = 5;
    exp_47_ram[1317] = 159;
    exp_47_ram[1318] = 0;
    exp_47_ram[1319] = 7;
    exp_47_ram[1320] = 0;
    exp_47_ram[1321] = 0;
    exp_47_ram[1322] = 95;
    exp_47_ram[1323] = 164;
    exp_47_ram[1324] = 164;
    exp_47_ram[1325] = 180;
    exp_47_ram[1326] = 137;
    exp_47_ram[1327] = 148;
    exp_47_ram[1328] = 137;
    exp_47_ram[1329] = 193;
    exp_47_ram[1330] = 129;
    exp_47_ram[1331] = 169;
    exp_47_ram[1332] = 65;
    exp_47_ram[1333] = 1;
    exp_47_ram[1334] = 1;
    exp_47_ram[1335] = 0;
    exp_47_ram[1336] = 1;
    exp_47_ram[1337] = 0;
    exp_47_ram[1338] = 145;
    exp_47_ram[1339] = 96;
    exp_47_ram[1340] = 5;
    exp_47_ram[1341] = 133;
    exp_47_ram[1342] = 1;
    exp_47_ram[1343] = 17;
    exp_47_ram[1344] = 129;
    exp_47_ram[1345] = 33;
    exp_47_ram[1346] = 49;
    exp_47_ram[1347] = 65;
    exp_47_ram[1348] = 159;
    exp_47_ram[1349] = 0;
    exp_47_ram[1350] = 80;
    exp_47_ram[1351] = 5;
    exp_47_ram[1352] = 129;
    exp_47_ram[1353] = 95;
    exp_47_ram[1354] = 132;
    exp_47_ram[1355] = 0;
    exp_47_ram[1356] = 137;
    exp_47_ram[1357] = 23;
    exp_47_ram[1358] = 245;
    exp_47_ram[1359] = 1;
    exp_47_ram[1360] = 0;
    exp_47_ram[1361] = 183;
    exp_47_ram[1362] = 48;
    exp_47_ram[1363] = 137;
    exp_47_ram[1364] = 143;
    exp_47_ram[1365] = 36;
    exp_47_ram[1366] = 4;
    exp_47_ram[1367] = 48;
    exp_47_ram[1368] = 68;
    exp_47_ram[1369] = 23;
    exp_47_ram[1370] = 245;
    exp_47_ram[1371] = 129;
    exp_47_ram[1372] = 183;
    exp_47_ram[1373] = 79;
    exp_47_ram[1374] = 36;
    exp_47_ram[1375] = 196;
    exp_47_ram[1376] = 160;
    exp_47_ram[1377] = 160;
    exp_47_ram[1378] = 208;
    exp_47_ram[1379] = 161;
    exp_47_ram[1380] = 129;
    exp_47_ram[1381] = 177;
    exp_47_ram[1382] = 36;
    exp_47_ram[1383] = 7;
    exp_47_ram[1384] = 244;
    exp_47_ram[1385] = 193;
    exp_47_ram[1386] = 160;
    exp_47_ram[1387] = 7;
    exp_47_ram[1388] = 244;
    exp_47_ram[1389] = 132;
    exp_47_ram[1390] = 208;
    exp_47_ram[1391] = 161;
    exp_47_ram[1392] = 129;
    exp_47_ram[1393] = 177;
    exp_47_ram[1394] = 68;
    exp_47_ram[1395] = 7;
    exp_47_ram[1396] = 244;
    exp_47_ram[1397] = 193;
    exp_47_ram[1398] = 160;
    exp_47_ram[1399] = 7;
    exp_47_ram[1400] = 244;
    exp_47_ram[1401] = 68;
    exp_47_ram[1402] = 208;
    exp_47_ram[1403] = 161;
    exp_47_ram[1404] = 129;
    exp_47_ram[1405] = 177;
    exp_47_ram[1406] = 68;
    exp_47_ram[1407] = 7;
    exp_47_ram[1408] = 244;
    exp_47_ram[1409] = 193;
    exp_47_ram[1410] = 160;
    exp_47_ram[1411] = 7;
    exp_47_ram[1412] = 244;
    exp_47_ram[1413] = 4;
    exp_47_ram[1414] = 208;
    exp_47_ram[1415] = 161;
    exp_47_ram[1416] = 129;
    exp_47_ram[1417] = 177;
    exp_47_ram[1418] = 36;
    exp_47_ram[1419] = 7;
    exp_47_ram[1420] = 244;
    exp_47_ram[1421] = 193;
    exp_47_ram[1422] = 128;
    exp_47_ram[1423] = 7;
    exp_47_ram[1424] = 244;
    exp_47_ram[1425] = 68;
    exp_47_ram[1426] = 197;
    exp_47_ram[1427] = 144;
    exp_47_ram[1428] = 161;
    exp_47_ram[1429] = 177;
    exp_47_ram[1430] = 129;
    exp_47_ram[1431] = 193;
    exp_47_ram[1432] = 64;
    exp_47_ram[1433] = 7;
    exp_47_ram[1434] = 244;
    exp_47_ram[1435] = 144;
    exp_47_ram[1436] = 161;
    exp_47_ram[1437] = 177;
    exp_47_ram[1438] = 129;
    exp_47_ram[1439] = 193;
    exp_47_ram[1440] = 160;
    exp_47_ram[1441] = 7;
    exp_47_ram[1442] = 244;
    exp_47_ram[1443] = 144;
    exp_47_ram[1444] = 161;
    exp_47_ram[1445] = 129;
    exp_47_ram[1446] = 177;
    exp_47_ram[1447] = 193;
    exp_47_ram[1448] = 7;
    exp_47_ram[1449] = 244;
    exp_47_ram[1450] = 193;
    exp_47_ram[1451] = 65;
    exp_47_ram[1452] = 1;
    exp_47_ram[1453] = 7;
    exp_47_ram[1454] = 244;
    exp_47_ram[1455] = 160;
    exp_47_ram[1456] = 244;
    exp_47_ram[1457] = 129;
    exp_47_ram[1458] = 129;
    exp_47_ram[1459] = 137;
    exp_47_ram[1460] = 193;
    exp_47_ram[1461] = 1;
    exp_47_ram[1462] = 0;
    exp_47_ram[1463] = 1;
    exp_47_ram[1464] = 97;
    exp_47_ram[1465] = 1;
    exp_47_ram[1466] = 129;
    exp_47_ram[1467] = 145;
    exp_47_ram[1468] = 33;
    exp_47_ram[1469] = 49;
    exp_47_ram[1470] = 81;
    exp_47_ram[1471] = 17;
    exp_47_ram[1472] = 65;
    exp_47_ram[1473] = 113;
    exp_47_ram[1474] = 129;
    exp_47_ram[1475] = 145;
    exp_47_ram[1476] = 5;
    exp_47_ram[1477] = 5;
    exp_47_ram[1478] = 6;
    exp_47_ram[1479] = 32;
    exp_47_ram[1480] = 64;
    exp_47_ram[1481] = 11;
    exp_47_ram[1482] = 9;
    exp_47_ram[1483] = 31;
    exp_47_ram[1484] = 160;
    exp_47_ram[1485] = 218;
    exp_47_ram[1486] = 11;
    exp_47_ram[1487] = 10;
    exp_47_ram[1488] = 207;
    exp_47_ram[1489] = 25;
    exp_47_ram[1490] = 9;
    exp_47_ram[1491] = 164;
    exp_47_ram[1492] = 164;
    exp_47_ram[1493] = 164;
    exp_47_ram[1494] = 74;
    exp_47_ram[1495] = 5;
    exp_47_ram[1496] = 233;
    exp_47_ram[1497] = 7;
    exp_47_ram[1498] = 31;
    exp_47_ram[1499] = 1;
    exp_47_ram[1500] = 0;
    exp_47_ram[1501] = 0;
    exp_47_ram[1502] = 12;
    exp_47_ram[1503] = 12;
    exp_47_ram[1504] = 9;
    exp_47_ram[1505] = 31;
    exp_47_ram[1506] = 12;
    exp_47_ram[1507] = 12;
    exp_47_ram[1508] = 5;
    exp_47_ram[1509] = 28;
    exp_47_ram[1510] = 79;
    exp_47_ram[1511] = 9;
    exp_47_ram[1512] = 164;
    exp_47_ram[1513] = 164;
    exp_47_ram[1514] = 164;
    exp_47_ram[1515] = 122;
    exp_47_ram[1516] = 122;
    exp_47_ram[1517] = 5;
    exp_47_ram[1518] = 249;
    exp_47_ram[1519] = 31;
    exp_47_ram[1520] = 1;
    exp_47_ram[1521] = 4;
    exp_47_ram[1522] = 5;
    exp_47_ram[1523] = 144;
    exp_47_ram[1524] = 177;
    exp_47_ram[1525] = 5;
    exp_47_ram[1526] = 161;
    exp_47_ram[1527] = 170;
    exp_47_ram[1528] = 193;
    exp_47_ram[1529] = 0;
    exp_47_ram[1530] = 5;
    exp_47_ram[1531] = 144;
    exp_47_ram[1532] = 177;
    exp_47_ram[1533] = 5;
    exp_47_ram[1534] = 161;
    exp_47_ram[1535] = 193;
    exp_47_ram[1536] = 192;
    exp_47_ram[1537] = 73;
    exp_47_ram[1538] = 208;
    exp_47_ram[1539] = 20;
    exp_47_ram[1540] = 161;
    exp_47_ram[1541] = 177;
    exp_47_ram[1542] = 180;
    exp_47_ram[1543] = 164;
    exp_47_ram[1544] = 36;
    exp_47_ram[1545] = 100;
    exp_47_ram[1546] = 52;
    exp_47_ram[1547] = 154;
    exp_47_ram[1548] = 244;
    exp_47_ram[1549] = 112;
    exp_47_ram[1550] = 207;
    exp_47_ram[1551] = 164;
    exp_47_ram[1552] = 68;
    exp_47_ram[1553] = 193;
    exp_47_ram[1554] = 4;
    exp_47_ram[1555] = 129;
    exp_47_ram[1556] = 65;
    exp_47_ram[1557] = 1;
    exp_47_ram[1558] = 193;
    exp_47_ram[1559] = 129;
    exp_47_ram[1560] = 65;
    exp_47_ram[1561] = 1;
    exp_47_ram[1562] = 193;
    exp_47_ram[1563] = 129;
    exp_47_ram[1564] = 65;
    exp_47_ram[1565] = 1;
    exp_47_ram[1566] = 0;
    exp_47_ram[1567] = 1;
    exp_47_ram[1568] = 81;
    exp_47_ram[1569] = 69;
    exp_47_ram[1570] = 144;
    exp_47_ram[1571] = 145;
    exp_47_ram[1572] = 33;
    exp_47_ram[1573] = 65;
    exp_47_ram[1574] = 240;
    exp_47_ram[1575] = 16;
    exp_47_ram[1576] = 64;
    exp_47_ram[1577] = 5;
    exp_47_ram[1578] = 129;
    exp_47_ram[1579] = 1;
    exp_47_ram[1580] = 17;
    exp_47_ram[1581] = 241;
    exp_47_ram[1582] = 129;
    exp_47_ram[1583] = 49;
    exp_47_ram[1584] = 65;
    exp_47_ram[1585] = 145;
    exp_47_ram[1586] = 81;
    exp_47_ram[1587] = 1;
    exp_47_ram[1588] = 1;
    exp_47_ram[1589] = 1;
    exp_47_ram[1590] = 15;
    exp_47_ram[1591] = 1;
    exp_47_ram[1592] = 159;
    exp_47_ram[1593] = 5;
    exp_47_ram[1594] = 5;
    exp_47_ram[1595] = 129;
    exp_47_ram[1596] = 223;
    exp_47_ram[1597] = 1;
    exp_47_ram[1598] = 65;
    exp_47_ram[1599] = 64;
    exp_47_ram[1600] = 129;
    exp_47_ram[1601] = 231;
    exp_47_ram[1602] = 1;
    exp_47_ram[1603] = 241;
    exp_47_ram[1604] = 143;
    exp_47_ram[1605] = 1;
    exp_47_ram[1606] = 31;
    exp_47_ram[1607] = 32;
    exp_47_ram[1608] = 64;
    exp_47_ram[1609] = 5;
    exp_47_ram[1610] = 5;
    exp_47_ram[1611] = 1;
    exp_47_ram[1612] = 193;
    exp_47_ram[1613] = 241;
    exp_47_ram[1614] = 65;
    exp_47_ram[1615] = 145;
    exp_47_ram[1616] = 81;
    exp_47_ram[1617] = 1;
    exp_47_ram[1618] = 1;
    exp_47_ram[1619] = 207;
    exp_47_ram[1620] = 1;
    exp_47_ram[1621] = 95;
    exp_47_ram[1622] = 5;
    exp_47_ram[1623] = 5;
    exp_47_ram[1624] = 193;
    exp_47_ram[1625] = 159;
    exp_47_ram[1626] = 65;
    exp_47_ram[1627] = 129;
    exp_47_ram[1628] = 64;
    exp_47_ram[1629] = 193;
    exp_47_ram[1630] = 231;
    exp_47_ram[1631] = 1;
    exp_47_ram[1632] = 241;
    exp_47_ram[1633] = 79;
    exp_47_ram[1634] = 1;
    exp_47_ram[1635] = 223;
    exp_47_ram[1636] = 5;
    exp_47_ram[1637] = 5;
    exp_47_ram[1638] = 64;
    exp_47_ram[1639] = 9;
    exp_47_ram[1640] = 1;
    exp_47_ram[1641] = 79;
    exp_47_ram[1642] = 1;
    exp_47_ram[1643] = 223;
    exp_47_ram[1644] = 149;
    exp_47_ram[1645] = 5;
    exp_47_ram[1646] = 5;
    exp_47_ram[1647] = 180;
    exp_47_ram[1648] = 69;
    exp_47_ram[1649] = 16;
    exp_47_ram[1650] = 135;
    exp_47_ram[1651] = 244;
    exp_47_ram[1652] = 55;
    exp_47_ram[1653] = 0;
    exp_47_ram[1654] = 193;
    exp_47_ram[1655] = 129;
    exp_47_ram[1656] = 65;
    exp_47_ram[1657] = 1;
    exp_47_ram[1658] = 193;
    exp_47_ram[1659] = 129;
    exp_47_ram[1660] = 65;
    exp_47_ram[1661] = 1;
    exp_47_ram[1662] = 0;
    exp_47_ram[1663] = 1;
    exp_47_ram[1664] = 5;
    exp_47_ram[1665] = 33;
    exp_47_ram[1666] = 64;
    exp_47_ram[1667] = 5;
    exp_47_ram[1668] = 193;
    exp_47_ram[1669] = 17;
    exp_47_ram[1670] = 129;
    exp_47_ram[1671] = 145;
    exp_47_ram[1672] = 49;
    exp_47_ram[1673] = 79;
    exp_47_ram[1674] = 64;
    exp_47_ram[1675] = 193;
    exp_47_ram[1676] = 1;
    exp_47_ram[1677] = 9;
    exp_47_ram[1678] = 15;
    exp_47_ram[1679] = 1;
    exp_47_ram[1680] = 159;
    exp_47_ram[1681] = 5;
    exp_47_ram[1682] = 5;
    exp_47_ram[1683] = 48;
    exp_47_ram[1684] = 255;
    exp_47_ram[1685] = 7;
    exp_47_ram[1686] = 245;
    exp_47_ram[1687] = 167;
    exp_47_ram[1688] = 245;
    exp_47_ram[1689] = 7;
    exp_47_ram[1690] = 135;
    exp_47_ram[1691] = 4;
    exp_47_ram[1692] = 4;
    exp_47_ram[1693] = 1;
    exp_47_ram[1694] = 95;
    exp_47_ram[1695] = 64;
    exp_47_ram[1696] = 1;
    exp_47_ram[1697] = 9;
    exp_47_ram[1698] = 15;
    exp_47_ram[1699] = 48;
    exp_47_ram[1700] = 16;
    exp_47_ram[1701] = 249;
    exp_47_ram[1702] = 193;
    exp_47_ram[1703] = 4;
    exp_47_ram[1704] = 129;
    exp_47_ram[1705] = 1;
    exp_47_ram[1706] = 193;
    exp_47_ram[1707] = 4;
    exp_47_ram[1708] = 65;
    exp_47_ram[1709] = 1;
    exp_47_ram[1710] = 0;
    exp_47_ram[1711] = 9;
    exp_47_ram[1712] = 64;
    exp_47_ram[1713] = 193;
    exp_47_ram[1714] = 1;
    exp_47_ram[1715] = 207;
    exp_47_ram[1716] = 1;
    exp_47_ram[1717] = 159;
    exp_47_ram[1718] = 0;
    exp_47_ram[1719] = 5;
    exp_47_ram[1720] = 0;
    exp_47_ram[1721] = 7;
    exp_47_ram[1722] = 244;
    exp_47_ram[1723] = 244;
    exp_47_ram[1724] = 228;
    exp_47_ram[1725] = 7;
    exp_47_ram[1726] = 95;
    exp_47_ram[1727] = 9;
    exp_47_ram[1728] = 64;
    exp_47_ram[1729] = 193;
    exp_47_ram[1730] = 1;
    exp_47_ram[1731] = 207;
    exp_47_ram[1732] = 1;
    exp_47_ram[1733] = 159;
    exp_47_ram[1734] = 169;
    exp_47_ram[1735] = 223;
    exp_47_ram[1736] = 9;
    exp_47_ram[1737] = 95;
    exp_47_ram[1738] = 1;
    exp_47_ram[1739] = 5;
    exp_47_ram[1740] = 5;
    exp_47_ram[1741] = 193;
    exp_47_ram[1742] = 17;
    exp_47_ram[1743] = 31;
    exp_47_ram[1744] = 193;
    exp_47_ram[1745] = 64;
    exp_47_ram[1746] = 1;
    exp_47_ram[1747] = 207;
    exp_47_ram[1748] = 1;
    exp_47_ram[1749] = 159;
    exp_47_ram[1750] = 193;
    exp_47_ram[1751] = 1;
    exp_47_ram[1752] = 0;
    exp_47_ram[1753] = 5;
    exp_47_ram[1754] = 69;
    exp_47_ram[1755] = 1;
    exp_47_ram[1756] = 1;
    exp_47_ram[1757] = 17;
    exp_47_ram[1758] = 129;
    exp_47_ram[1759] = 31;
    exp_47_ram[1760] = 0;
    exp_47_ram[1761] = 1;
    exp_47_ram[1762] = 68;
    exp_47_ram[1763] = 64;
    exp_47_ram[1764] = 143;
    exp_47_ram[1765] = 193;
    exp_47_ram[1766] = 68;
    exp_47_ram[1767] = 129;
    exp_47_ram[1768] = 1;
    exp_47_ram[1769] = 0;
    exp_47_ram[1770] = 1;
    exp_47_ram[1771] = 145;
    exp_47_ram[1772] = 33;
    exp_47_ram[1773] = 69;
    exp_47_ram[1774] = 5;
    exp_47_ram[1775] = 17;
    exp_47_ram[1776] = 4;
    exp_47_ram[1777] = 9;
    exp_47_ram[1778] = 129;
    exp_47_ram[1779] = 49;
    exp_47_ram[1780] = 159;
    exp_47_ram[1781] = 0;
    exp_47_ram[1782] = 5;
    exp_47_ram[1783] = 0;
    exp_47_ram[1784] = 6;
    exp_47_ram[1785] = 38;
    exp_47_ram[1786] = 197;
    exp_47_ram[1787] = 150;
    exp_47_ram[1788] = 1;
    exp_47_ram[1789] = 159;
    exp_47_ram[1790] = 0;
    exp_47_ram[1791] = 1;
    exp_47_ram[1792] = 64;
    exp_47_ram[1793] = 68;
    exp_47_ram[1794] = 15;
    exp_47_ram[1795] = 9;
    exp_47_ram[1796] = 4;
    exp_47_ram[1797] = 95;
    exp_47_ram[1798] = 68;
    exp_47_ram[1799] = 169;
    exp_47_ram[1800] = 193;
    exp_47_ram[1801] = 68;
    exp_47_ram[1802] = 129;
    exp_47_ram[1803] = 65;
    exp_47_ram[1804] = 1;
    exp_47_ram[1805] = 193;
    exp_47_ram[1806] = 1;
    exp_47_ram[1807] = 0;
    exp_47_ram[1808] = 1;
    exp_47_ram[1809] = 17;
    exp_47_ram[1810] = 31;
    exp_47_ram[1811] = 193;
    exp_47_ram[1812] = 1;
    exp_47_ram[1813] = 223;
    exp_47_ram[1814] = 1;
    exp_47_ram[1815] = 17;
    exp_47_ram[1816] = 129;
    exp_47_ram[1817] = 1;
    exp_47_ram[1818] = 0;
    exp_47_ram[1819] = 7;
    exp_47_ram[1820] = 15;
    exp_47_ram[1821] = 68;
    exp_47_ram[1822] = 0;
    exp_47_ram[1823] = 135;
    exp_47_ram[1824] = 231;
    exp_47_ram[1825] = 7;
    exp_47_ram[1826] = 68;
    exp_47_ram[1827] = 7;
    exp_47_ram[1828] = 207;
    exp_47_ram[1829] = 5;
    exp_47_ram[1830] = 7;
    exp_47_ram[1831] = 68;
    exp_47_ram[1832] = 231;
    exp_47_ram[1833] = 0;
    exp_47_ram[1834] = 199;
    exp_47_ram[1835] = 199;
    exp_47_ram[1836] = 22;
    exp_47_ram[1837] = 199;
    exp_47_ram[1838] = 38;
    exp_47_ram[1839] = 199;
    exp_47_ram[1840] = 55;
    exp_47_ram[1841] = 183;
    exp_47_ram[1842] = 199;
    exp_47_ram[1843] = 215;
    exp_47_ram[1844] = 231;
    exp_47_ram[1845] = 68;
    exp_47_ram[1846] = 0;
    exp_47_ram[1847] = 7;
    exp_47_ram[1848] = 7;
    exp_47_ram[1849] = 79;
    exp_47_ram[1850] = 5;
    exp_47_ram[1851] = 7;
    exp_47_ram[1852] = 0;
    exp_47_ram[1853] = 135;
    exp_47_ram[1854] = 159;
    exp_47_ram[1855] = 208;
    exp_47_ram[1856] = 4;
    exp_47_ram[1857] = 68;
    exp_47_ram[1858] = 7;
    exp_47_ram[1859] = 15;
    exp_47_ram[1860] = 5;
    exp_47_ram[1861] = 7;
    exp_47_ram[1862] = 68;
    exp_47_ram[1863] = 231;
    exp_47_ram[1864] = 0;
    exp_47_ram[1865] = 199;
    exp_47_ram[1866] = 199;
    exp_47_ram[1867] = 22;
    exp_47_ram[1868] = 199;
    exp_47_ram[1869] = 38;
    exp_47_ram[1870] = 199;
    exp_47_ram[1871] = 55;
    exp_47_ram[1872] = 183;
    exp_47_ram[1873] = 199;
    exp_47_ram[1874] = 215;
    exp_47_ram[1875] = 231;
    exp_47_ram[1876] = 68;
    exp_47_ram[1877] = 0;
    exp_47_ram[1878] = 199;
    exp_47_ram[1879] = 7;
    exp_47_ram[1880] = 143;
    exp_47_ram[1881] = 5;
    exp_47_ram[1882] = 7;
    exp_47_ram[1883] = 0;
    exp_47_ram[1884] = 7;
    exp_47_ram[1885] = 223;
    exp_47_ram[1886] = 16;
    exp_47_ram[1887] = 68;
    exp_47_ram[1888] = 0;
    exp_47_ram[1889] = 135;
    exp_47_ram[1890] = 231;
    exp_47_ram[1891] = 7;
    exp_47_ram[1892] = 68;
    exp_47_ram[1893] = 0;
    exp_47_ram[1894] = 135;
    exp_47_ram[1895] = 7;
    exp_47_ram[1896] = 143;
    exp_47_ram[1897] = 5;
    exp_47_ram[1898] = 7;
    exp_47_ram[1899] = 0;
    exp_47_ram[1900] = 199;
    exp_47_ram[1901] = 223;
    exp_47_ram[1902] = 16;
    exp_47_ram[1903] = 4;
    exp_47_ram[1904] = 68;
    exp_47_ram[1905] = 7;
    exp_47_ram[1906] = 7;
    exp_47_ram[1907] = 0;
    exp_47_ram[1908] = 71;
    exp_47_ram[1909] = 223;
    exp_47_ram[1910] = 16;
    exp_47_ram[1911] = 0;
    exp_47_ram[1912] = 199;
    exp_47_ram[1913] = 223;
    exp_47_ram[1914] = 0;
    exp_47_ram[1915] = 71;
    exp_47_ram[1916] = 31;
    exp_47_ram[1917] = 68;
    exp_47_ram[1918] = 0;
    exp_47_ram[1919] = 135;
    exp_47_ram[1920] = 231;
    exp_47_ram[1921] = 7;
    exp_47_ram[1922] = 68;
    exp_47_ram[1923] = 48;
    exp_47_ram[1924] = 0;
    exp_47_ram[1925] = 7;
    exp_47_ram[1926] = 7;
    exp_47_ram[1927] = 95;
    exp_47_ram[1928] = 5;
    exp_47_ram[1929] = 0;
    exp_47_ram[1930] = 7;
    exp_47_ram[1931] = 7;
    exp_47_ram[1932] = 159;
    exp_47_ram[1933] = 5;
    exp_47_ram[1934] = 7;
    exp_47_ram[1935] = 0;
    exp_47_ram[1936] = 135;
    exp_47_ram[1937] = 223;
    exp_47_ram[1938] = 16;
    exp_47_ram[1939] = 4;
    exp_47_ram[1940] = 68;
    exp_47_ram[1941] = 48;
    exp_47_ram[1942] = 0;
    exp_47_ram[1943] = 7;
    exp_47_ram[1944] = 7;
    exp_47_ram[1945] = 223;
    exp_47_ram[1946] = 5;
    exp_47_ram[1947] = 0;
    exp_47_ram[1948] = 199;
    exp_47_ram[1949] = 7;
    exp_47_ram[1950] = 31;
    exp_47_ram[1951] = 5;
    exp_47_ram[1952] = 7;
    exp_47_ram[1953] = 0;
    exp_47_ram[1954] = 7;
    exp_47_ram[1955] = 95;
    exp_47_ram[1956] = 144;
    exp_47_ram[1957] = 68;
    exp_47_ram[1958] = 0;
    exp_47_ram[1959] = 135;
    exp_47_ram[1960] = 231;
    exp_47_ram[1961] = 7;
    exp_47_ram[1962] = 68;
    exp_47_ram[1963] = 0;
    exp_47_ram[1964] = 135;
    exp_47_ram[1965] = 7;
    exp_47_ram[1966] = 31;
    exp_47_ram[1967] = 5;
    exp_47_ram[1968] = 7;
    exp_47_ram[1969] = 0;
    exp_47_ram[1970] = 199;
    exp_47_ram[1971] = 95;
    exp_47_ram[1972] = 144;
    exp_47_ram[1973] = 4;
    exp_47_ram[1974] = 68;
    exp_47_ram[1975] = 7;
    exp_47_ram[1976] = 7;
    exp_47_ram[1977] = 0;
    exp_47_ram[1978] = 71;
    exp_47_ram[1979] = 95;
    exp_47_ram[1980] = 144;
    exp_47_ram[1981] = 0;
    exp_47_ram[1982] = 199;
    exp_47_ram[1983] = 95;
    exp_47_ram[1984] = 0;
    exp_47_ram[1985] = 135;
    exp_47_ram[1986] = 159;
    exp_47_ram[1987] = 0;
    exp_47_ram[1988] = 199;
    exp_47_ram[1989] = 223;
    exp_47_ram[1990] = 0;
    exp_47_ram[1991] = 71;
    exp_47_ram[1992] = 31;
    exp_47_ram[1993] = 0;
    exp_47_ram[1994] = 199;
    exp_47_ram[1995] = 95;
    exp_47_ram[1996] = 0;
    exp_47_ram[1997] = 7;
    exp_47_ram[1998] = 159;
    exp_47_ram[1999] = 0;
    exp_47_ram[2000] = 199;
    exp_47_ram[2001] = 223;
    exp_47_ram[2002] = 0;
    exp_47_ram[2003] = 199;
    exp_47_ram[2004] = 31;
    exp_47_ram[2005] = 68;
    exp_47_ram[2006] = 51;
    exp_47_ram[2007] = 23;
    exp_47_ram[2008] = 231;
    exp_47_ram[2009] = 7;
    exp_47_ram[2010] = 68;
    exp_47_ram[2011] = 80;
    exp_47_ram[2012] = 16;
    exp_47_ram[2013] = 7;
    exp_47_ram[2014] = 31;
    exp_47_ram[2015] = 5;
    exp_47_ram[2016] = 68;
    exp_47_ram[2017] = 247;
    exp_47_ram[2018] = 0;
    exp_47_ram[2019] = 135;
    exp_47_ram[2020] = 31;
    exp_47_ram[2021] = 80;
    exp_47_ram[2022] = 68;
    exp_47_ram[2023] = 80;
    exp_47_ram[2024] = 32;
    exp_47_ram[2025] = 7;
    exp_47_ram[2026] = 31;
    exp_47_ram[2027] = 5;
    exp_47_ram[2028] = 68;
    exp_47_ram[2029] = 247;
    exp_47_ram[2030] = 16;
    exp_47_ram[2031] = 247;
    exp_47_ram[2032] = 0;
    exp_47_ram[2033] = 7;
    exp_47_ram[2034] = 159;
    exp_47_ram[2035] = 208;
    exp_47_ram[2036] = 68;
    exp_47_ram[2037] = 80;
    exp_47_ram[2038] = 48;
    exp_47_ram[2039] = 7;
    exp_47_ram[2040] = 159;
    exp_47_ram[2041] = 5;
    exp_47_ram[2042] = 68;
    exp_47_ram[2043] = 247;
    exp_47_ram[2044] = 32;
    exp_47_ram[2045] = 247;
    exp_47_ram[2046] = 0;
    exp_47_ram[2047] = 199;
    exp_47_ram[2048] = 31;
    exp_47_ram[2049] = 80;
    exp_47_ram[2050] = 68;
    exp_47_ram[2051] = 80;
    exp_47_ram[2052] = 64;
    exp_47_ram[2053] = 7;
    exp_47_ram[2054] = 31;
    exp_47_ram[2055] = 5;
    exp_47_ram[2056] = 68;
    exp_47_ram[2057] = 247;
    exp_47_ram[2058] = 48;
    exp_47_ram[2059] = 247;
    exp_47_ram[2060] = 0;
    exp_47_ram[2061] = 71;
    exp_47_ram[2062] = 159;
    exp_47_ram[2063] = 208;
    exp_47_ram[2064] = 68;
    exp_47_ram[2065] = 80;
    exp_47_ram[2066] = 80;
    exp_47_ram[2067] = 7;
    exp_47_ram[2068] = 159;
    exp_47_ram[2069] = 5;
    exp_47_ram[2070] = 7;
    exp_47_ram[2071] = 0;
    exp_47_ram[2072] = 135;
    exp_47_ram[2073] = 223;
    exp_47_ram[2074] = 16;
    exp_47_ram[2075] = 0;
    exp_47_ram[2076] = 199;
    exp_47_ram[2077] = 223;
    exp_47_ram[2078] = 0;
    exp_47_ram[2079] = 7;
    exp_47_ram[2080] = 31;
    exp_47_ram[2081] = 68;
    exp_47_ram[2082] = 51;
    exp_47_ram[2083] = 23;
    exp_47_ram[2084] = 231;
    exp_47_ram[2085] = 51;
    exp_47_ram[2086] = 23;
    exp_47_ram[2087] = 231;
    exp_47_ram[2088] = 7;
    exp_47_ram[2089] = 68;
    exp_47_ram[2090] = 16;
    exp_47_ram[2091] = 7;
    exp_47_ram[2092] = 31;
    exp_47_ram[2093] = 5;
    exp_47_ram[2094] = 68;
    exp_47_ram[2095] = 247;
    exp_47_ram[2096] = 0;
    exp_47_ram[2097] = 135;
    exp_47_ram[2098] = 159;
    exp_47_ram[2099] = 208;
    exp_47_ram[2100] = 68;
    exp_47_ram[2101] = 32;
    exp_47_ram[2102] = 7;
    exp_47_ram[2103] = 95;
    exp_47_ram[2104] = 5;
    exp_47_ram[2105] = 68;
    exp_47_ram[2106] = 247;
    exp_47_ram[2107] = 16;
    exp_47_ram[2108] = 247;
    exp_47_ram[2109] = 0;
    exp_47_ram[2110] = 7;
    exp_47_ram[2111] = 95;
    exp_47_ram[2112] = 128;
    exp_47_ram[2113] = 68;
    exp_47_ram[2114] = 48;
    exp_47_ram[2115] = 7;
    exp_47_ram[2116] = 31;
    exp_47_ram[2117] = 5;
    exp_47_ram[2118] = 68;
    exp_47_ram[2119] = 247;
    exp_47_ram[2120] = 32;
    exp_47_ram[2121] = 247;
    exp_47_ram[2122] = 0;
    exp_47_ram[2123] = 199;
    exp_47_ram[2124] = 31;
    exp_47_ram[2125] = 64;
    exp_47_ram[2126] = 68;
    exp_47_ram[2127] = 64;
    exp_47_ram[2128] = 7;
    exp_47_ram[2129] = 223;
    exp_47_ram[2130] = 5;
    exp_47_ram[2131] = 68;
    exp_47_ram[2132] = 247;
    exp_47_ram[2133] = 48;
    exp_47_ram[2134] = 247;
    exp_47_ram[2135] = 0;
    exp_47_ram[2136] = 71;
    exp_47_ram[2137] = 223;
    exp_47_ram[2138] = 0;
    exp_47_ram[2139] = 68;
    exp_47_ram[2140] = 7;
    exp_47_ram[2141] = 159;
    exp_47_ram[2142] = 5;
    exp_47_ram[2143] = 7;
    exp_47_ram[2144] = 68;
    exp_47_ram[2145] = 231;
    exp_47_ram[2146] = 68;
    exp_47_ram[2147] = 247;
    exp_47_ram[2148] = 128;
    exp_47_ram[2149] = 247;
    exp_47_ram[2150] = 0;
    exp_47_ram[2151] = 135;
    exp_47_ram[2152] = 31;
    exp_47_ram[2153] = 64;
    exp_47_ram[2154] = 68;
    exp_47_ram[2155] = 80;
    exp_47_ram[2156] = 7;
    exp_47_ram[2157] = 223;
    exp_47_ram[2158] = 5;
    exp_47_ram[2159] = 7;
    exp_47_ram[2160] = 0;
    exp_47_ram[2161] = 199;
    exp_47_ram[2162] = 159;
    exp_47_ram[2163] = 192;
    exp_47_ram[2164] = 0;
    exp_47_ram[2165] = 199;
    exp_47_ram[2166] = 159;
    exp_47_ram[2167] = 0;
    exp_47_ram[2168] = 71;
    exp_47_ram[2169] = 223;
    exp_47_ram[2170] = 68;
    exp_47_ram[2171] = 51;
    exp_47_ram[2172] = 23;
    exp_47_ram[2173] = 231;
    exp_47_ram[2174] = 7;
    exp_47_ram[2175] = 68;
    exp_47_ram[2176] = 0;
    exp_47_ram[2177] = 7;
    exp_47_ram[2178] = 7;
    exp_47_ram[2179] = 31;
    exp_47_ram[2180] = 5;
    exp_47_ram[2181] = 7;
    exp_47_ram[2182] = 0;
    exp_47_ram[2183] = 135;
    exp_47_ram[2184] = 31;
    exp_47_ram[2185] = 64;
    exp_47_ram[2186] = 68;
    exp_47_ram[2187] = 0;
    exp_47_ram[2188] = 135;
    exp_47_ram[2189] = 7;
    exp_47_ram[2190] = 95;
    exp_47_ram[2191] = 5;
    exp_47_ram[2192] = 16;
    exp_47_ram[2193] = 247;
    exp_47_ram[2194] = 0;
    exp_47_ram[2195] = 7;
    exp_47_ram[2196] = 31;
    exp_47_ram[2197] = 64;
    exp_47_ram[2198] = 68;
    exp_47_ram[2199] = 0;
    exp_47_ram[2200] = 71;
    exp_47_ram[2201] = 7;
    exp_47_ram[2202] = 95;
    exp_47_ram[2203] = 5;
    exp_47_ram[2204] = 32;
    exp_47_ram[2205] = 247;
    exp_47_ram[2206] = 0;
    exp_47_ram[2207] = 199;
    exp_47_ram[2208] = 31;
    exp_47_ram[2209] = 64;
    exp_47_ram[2210] = 68;
    exp_47_ram[2211] = 0;
    exp_47_ram[2212] = 7;
    exp_47_ram[2213] = 7;
    exp_47_ram[2214] = 95;
    exp_47_ram[2215] = 5;
    exp_47_ram[2216] = 48;
    exp_47_ram[2217] = 247;
    exp_47_ram[2218] = 0;
    exp_47_ram[2219] = 71;
    exp_47_ram[2220] = 31;
    exp_47_ram[2221] = 64;
    exp_47_ram[2222] = 68;
    exp_47_ram[2223] = 0;
    exp_47_ram[2224] = 199;
    exp_47_ram[2225] = 7;
    exp_47_ram[2226] = 95;
    exp_47_ram[2227] = 5;
    exp_47_ram[2228] = 64;
    exp_47_ram[2229] = 247;
    exp_47_ram[2230] = 0;
    exp_47_ram[2231] = 199;
    exp_47_ram[2232] = 31;
    exp_47_ram[2233] = 64;
    exp_47_ram[2234] = 0;
    exp_47_ram[2235] = 199;
    exp_47_ram[2236] = 31;
    exp_47_ram[2237] = 0;
    exp_47_ram[2238] = 135;
    exp_47_ram[2239] = 95;
    exp_47_ram[2240] = 68;
    exp_47_ram[2241] = 51;
    exp_47_ram[2242] = 23;
    exp_47_ram[2243] = 231;
    exp_47_ram[2244] = 7;
    exp_47_ram[2245] = 68;
    exp_47_ram[2246] = 0;
    exp_47_ram[2247] = 71;
    exp_47_ram[2248] = 7;
    exp_47_ram[2249] = 223;
    exp_47_ram[2250] = 5;
    exp_47_ram[2251] = 68;
    exp_47_ram[2252] = 247;
    exp_47_ram[2253] = 0;
    exp_47_ram[2254] = 135;
    exp_47_ram[2255] = 95;
    exp_47_ram[2256] = 128;
    exp_47_ram[2257] = 68;
    exp_47_ram[2258] = 0;
    exp_47_ram[2259] = 7;
    exp_47_ram[2260] = 7;
    exp_47_ram[2261] = 223;
    exp_47_ram[2262] = 5;
    exp_47_ram[2263] = 68;
    exp_47_ram[2264] = 247;
    exp_47_ram[2265] = 16;
    exp_47_ram[2266] = 247;
    exp_47_ram[2267] = 0;
    exp_47_ram[2268] = 7;
    exp_47_ram[2269] = 223;
    exp_47_ram[2270] = 0;
    exp_47_ram[2271] = 68;
    exp_47_ram[2272] = 0;
    exp_47_ram[2273] = 135;
    exp_47_ram[2274] = 7;
    exp_47_ram[2275] = 95;
    exp_47_ram[2276] = 5;
    exp_47_ram[2277] = 68;
    exp_47_ram[2278] = 247;
    exp_47_ram[2279] = 32;
    exp_47_ram[2280] = 247;
    exp_47_ram[2281] = 0;
    exp_47_ram[2282] = 199;
    exp_47_ram[2283] = 95;
    exp_47_ram[2284] = 128;
    exp_47_ram[2285] = 68;
    exp_47_ram[2286] = 0;
    exp_47_ram[2287] = 7;
    exp_47_ram[2288] = 7;
    exp_47_ram[2289] = 223;
    exp_47_ram[2290] = 5;
    exp_47_ram[2291] = 68;
    exp_47_ram[2292] = 247;
    exp_47_ram[2293] = 48;
    exp_47_ram[2294] = 247;
    exp_47_ram[2295] = 0;
    exp_47_ram[2296] = 71;
    exp_47_ram[2297] = 223;
    exp_47_ram[2298] = 0;
    exp_47_ram[2299] = 68;
    exp_47_ram[2300] = 0;
    exp_47_ram[2301] = 135;
    exp_47_ram[2302] = 7;
    exp_47_ram[2303] = 95;
    exp_47_ram[2304] = 5;
    exp_47_ram[2305] = 7;
    exp_47_ram[2306] = 0;
    exp_47_ram[2307] = 135;
    exp_47_ram[2308] = 31;
    exp_47_ram[2309] = 64;
    exp_47_ram[2310] = 0;
    exp_47_ram[2311] = 199;
    exp_47_ram[2312] = 31;
    exp_47_ram[2313] = 0;
    exp_47_ram[2314] = 71;
    exp_47_ram[2315] = 95;
    exp_47_ram[2316] = 68;
    exp_47_ram[2317] = 51;
    exp_47_ram[2318] = 23;
    exp_47_ram[2319] = 231;
    exp_47_ram[2320] = 51;
    exp_47_ram[2321] = 23;
    exp_47_ram[2322] = 231;
    exp_47_ram[2323] = 7;
    exp_47_ram[2324] = 68;
    exp_47_ram[2325] = 16;
    exp_47_ram[2326] = 7;
    exp_47_ram[2327] = 159;
    exp_47_ram[2328] = 5;
    exp_47_ram[2329] = 68;
    exp_47_ram[2330] = 247;
    exp_47_ram[2331] = 64;
    exp_47_ram[2332] = 247;
    exp_47_ram[2333] = 0;
    exp_47_ram[2334] = 135;
    exp_47_ram[2335] = 95;
    exp_47_ram[2336] = 128;
    exp_47_ram[2337] = 68;
    exp_47_ram[2338] = 32;
    exp_47_ram[2339] = 7;
    exp_47_ram[2340] = 95;
    exp_47_ram[2341] = 5;
    exp_47_ram[2342] = 68;
    exp_47_ram[2343] = 247;
    exp_47_ram[2344] = 80;
    exp_47_ram[2345] = 247;
    exp_47_ram[2346] = 0;
    exp_47_ram[2347] = 7;
    exp_47_ram[2348] = 31;
    exp_47_ram[2349] = 64;
    exp_47_ram[2350] = 68;
    exp_47_ram[2351] = 48;
    exp_47_ram[2352] = 7;
    exp_47_ram[2353] = 31;
    exp_47_ram[2354] = 5;
    exp_47_ram[2355] = 68;
    exp_47_ram[2356] = 247;
    exp_47_ram[2357] = 96;
    exp_47_ram[2358] = 247;
    exp_47_ram[2359] = 0;
    exp_47_ram[2360] = 199;
    exp_47_ram[2361] = 223;
    exp_47_ram[2362] = 0;
    exp_47_ram[2363] = 68;
    exp_47_ram[2364] = 64;
    exp_47_ram[2365] = 7;
    exp_47_ram[2366] = 223;
    exp_47_ram[2367] = 5;
    exp_47_ram[2368] = 68;
    exp_47_ram[2369] = 247;
    exp_47_ram[2370] = 112;
    exp_47_ram[2371] = 247;
    exp_47_ram[2372] = 0;
    exp_47_ram[2373] = 71;
    exp_47_ram[2374] = 143;
    exp_47_ram[2375] = 192;
    exp_47_ram[2376] = 68;
    exp_47_ram[2377] = 7;
    exp_47_ram[2378] = 95;
    exp_47_ram[2379] = 5;
    exp_47_ram[2380] = 7;
    exp_47_ram[2381] = 68;
    exp_47_ram[2382] = 231;
    exp_47_ram[2383] = 68;
    exp_47_ram[2384] = 247;
    exp_47_ram[2385] = 128;
    exp_47_ram[2386] = 247;
    exp_47_ram[2387] = 0;
    exp_47_ram[2388] = 135;
    exp_47_ram[2389] = 207;
    exp_47_ram[2390] = 0;
    exp_47_ram[2391] = 68;
    exp_47_ram[2392] = 80;
    exp_47_ram[2393] = 7;
    exp_47_ram[2394] = 223;
    exp_47_ram[2395] = 5;
    exp_47_ram[2396] = 7;
    exp_47_ram[2397] = 0;
    exp_47_ram[2398] = 199;
    exp_47_ram[2399] = 79;
    exp_47_ram[2400] = 128;
    exp_47_ram[2401] = 0;
    exp_47_ram[2402] = 199;
    exp_47_ram[2403] = 79;
    exp_47_ram[2404] = 0;
    exp_47_ram[2405] = 7;
    exp_47_ram[2406] = 143;
    exp_47_ram[2407] = 68;
    exp_47_ram[2408] = 51;
    exp_47_ram[2409] = 23;
    exp_47_ram[2410] = 231;
    exp_47_ram[2411] = 7;
    exp_47_ram[2412] = 68;
    exp_47_ram[2413] = 0;
    exp_47_ram[2414] = 199;
    exp_47_ram[2415] = 7;
    exp_47_ram[2416] = 159;
    exp_47_ram[2417] = 5;
    exp_47_ram[2418] = 16;
    exp_47_ram[2419] = 247;
    exp_47_ram[2420] = 0;
    exp_47_ram[2421] = 135;
    exp_47_ram[2422] = 143;
    exp_47_ram[2423] = 192;
    exp_47_ram[2424] = 68;
    exp_47_ram[2425] = 0;
    exp_47_ram[2426] = 71;
    exp_47_ram[2427] = 7;
    exp_47_ram[2428] = 159;
    exp_47_ram[2429] = 5;
    exp_47_ram[2430] = 32;
    exp_47_ram[2431] = 247;
    exp_47_ram[2432] = 0;
    exp_47_ram[2433] = 7;
    exp_47_ram[2434] = 143;
    exp_47_ram[2435] = 192;
    exp_47_ram[2436] = 68;
    exp_47_ram[2437] = 0;
    exp_47_ram[2438] = 7;
    exp_47_ram[2439] = 7;
    exp_47_ram[2440] = 159;
    exp_47_ram[2441] = 5;
    exp_47_ram[2442] = 48;
    exp_47_ram[2443] = 247;
    exp_47_ram[2444] = 0;
    exp_47_ram[2445] = 199;
    exp_47_ram[2446] = 143;
    exp_47_ram[2447] = 192;
    exp_47_ram[2448] = 68;
    exp_47_ram[2449] = 0;
    exp_47_ram[2450] = 7;
    exp_47_ram[2451] = 7;
    exp_47_ram[2452] = 159;
    exp_47_ram[2453] = 5;
    exp_47_ram[2454] = 7;
    exp_47_ram[2455] = 0;
    exp_47_ram[2456] = 71;
    exp_47_ram[2457] = 207;
    exp_47_ram[2458] = 0;
    exp_47_ram[2459] = 68;
    exp_47_ram[2460] = 0;
    exp_47_ram[2461] = 199;
    exp_47_ram[2462] = 7;
    exp_47_ram[2463] = 223;
    exp_47_ram[2464] = 5;
    exp_47_ram[2465] = 64;
    exp_47_ram[2466] = 247;
    exp_47_ram[2467] = 0;
    exp_47_ram[2468] = 199;
    exp_47_ram[2469] = 207;
    exp_47_ram[2470] = 0;
    exp_47_ram[2471] = 0;
    exp_47_ram[2472] = 199;
    exp_47_ram[2473] = 207;
    exp_47_ram[2474] = 0;
    exp_47_ram[2475] = 199;
    exp_47_ram[2476] = 15;
    exp_47_ram[2477] = 68;
    exp_47_ram[2478] = 51;
    exp_47_ram[2479] = 23;
    exp_47_ram[2480] = 231;
    exp_47_ram[2481] = 7;
    exp_47_ram[2482] = 68;
    exp_47_ram[2483] = 0;
    exp_47_ram[2484] = 135;
    exp_47_ram[2485] = 7;
    exp_47_ram[2486] = 95;
    exp_47_ram[2487] = 5;
    exp_47_ram[2488] = 68;
    exp_47_ram[2489] = 247;
    exp_47_ram[2490] = 0;
    exp_47_ram[2491] = 135;
    exp_47_ram[2492] = 15;
    exp_47_ram[2493] = 64;
    exp_47_ram[2494] = 68;
    exp_47_ram[2495] = 0;
    exp_47_ram[2496] = 7;
    exp_47_ram[2497] = 7;
    exp_47_ram[2498] = 95;
    exp_47_ram[2499] = 5;
    exp_47_ram[2500] = 68;
    exp_47_ram[2501] = 247;
    exp_47_ram[2502] = 16;
    exp_47_ram[2503] = 247;
    exp_47_ram[2504] = 0;
    exp_47_ram[2505] = 7;
    exp_47_ram[2506] = 143;
    exp_47_ram[2507] = 192;
    exp_47_ram[2508] = 68;
    exp_47_ram[2509] = 0;
    exp_47_ram[2510] = 71;
    exp_47_ram[2511] = 7;
    exp_47_ram[2512] = 223;
    exp_47_ram[2513] = 5;
    exp_47_ram[2514] = 68;
    exp_47_ram[2515] = 247;
    exp_47_ram[2516] = 32;
    exp_47_ram[2517] = 247;
    exp_47_ram[2518] = 0;
    exp_47_ram[2519] = 199;
    exp_47_ram[2520] = 15;
    exp_47_ram[2521] = 64;
    exp_47_ram[2522] = 68;
    exp_47_ram[2523] = 64;
    exp_47_ram[2524] = 7;
    exp_47_ram[2525] = 207;
    exp_47_ram[2526] = 5;
    exp_47_ram[2527] = 68;
    exp_47_ram[2528] = 247;
    exp_47_ram[2529] = 48;
    exp_47_ram[2530] = 247;
    exp_47_ram[2531] = 0;
    exp_47_ram[2532] = 71;
    exp_47_ram[2533] = 207;
    exp_47_ram[2534] = 0;
    exp_47_ram[2535] = 68;
    exp_47_ram[2536] = 0;
    exp_47_ram[2537] = 199;
    exp_47_ram[2538] = 7;
    exp_47_ram[2539] = 31;
    exp_47_ram[2540] = 5;
    exp_47_ram[2541] = 7;
    exp_47_ram[2542] = 0;
    exp_47_ram[2543] = 199;
    exp_47_ram[2544] = 15;
    exp_47_ram[2545] = 64;
    exp_47_ram[2546] = 0;
    exp_47_ram[2547] = 199;
    exp_47_ram[2548] = 15;
    exp_47_ram[2549] = 0;
    exp_47_ram[2550] = 135;
    exp_47_ram[2551] = 79;
    exp_47_ram[2552] = 16;
    exp_47_ram[2553] = 244;
    exp_47_ram[2554] = 68;
    exp_47_ram[2555] = 0;
    exp_47_ram[2556] = 71;
    exp_47_ram[2557] = 7;
    exp_47_ram[2558] = 15;
    exp_47_ram[2559] = 5;
    exp_47_ram[2560] = 7;
    exp_47_ram[2561] = 0;
    exp_47_ram[2562] = 135;
    exp_47_ram[2563] = 79;
    exp_47_ram[2564] = 128;
    exp_47_ram[2565] = 68;
    exp_47_ram[2566] = 32;
    exp_47_ram[2567] = 32;
    exp_47_ram[2568] = 7;
    exp_47_ram[2569] = 143;
    exp_47_ram[2570] = 5;
    exp_47_ram[2571] = 0;
    exp_47_ram[2572] = 199;
    exp_47_ram[2573] = 7;
    exp_47_ram[2574] = 15;
    exp_47_ram[2575] = 5;
    exp_47_ram[2576] = 7;
    exp_47_ram[2577] = 0;
    exp_47_ram[2578] = 7;
    exp_47_ram[2579] = 79;
    exp_47_ram[2580] = 128;
    exp_47_ram[2581] = 68;
    exp_47_ram[2582] = 48;
    exp_47_ram[2583] = 48;
    exp_47_ram[2584] = 7;
    exp_47_ram[2585] = 143;
    exp_47_ram[2586] = 5;
    exp_47_ram[2587] = 0;
    exp_47_ram[2588] = 71;
    exp_47_ram[2589] = 7;
    exp_47_ram[2590] = 15;
    exp_47_ram[2591] = 5;
    exp_47_ram[2592] = 7;
    exp_47_ram[2593] = 0;
    exp_47_ram[2594] = 199;
    exp_47_ram[2595] = 79;
    exp_47_ram[2596] = 128;
    exp_47_ram[2597] = 68;
    exp_47_ram[2598] = 64;
    exp_47_ram[2599] = 64;
    exp_47_ram[2600] = 7;
    exp_47_ram[2601] = 143;
    exp_47_ram[2602] = 5;
    exp_47_ram[2603] = 0;
    exp_47_ram[2604] = 199;
    exp_47_ram[2605] = 7;
    exp_47_ram[2606] = 15;
    exp_47_ram[2607] = 5;
    exp_47_ram[2608] = 7;
    exp_47_ram[2609] = 0;
    exp_47_ram[2610] = 71;
    exp_47_ram[2611] = 79;
    exp_47_ram[2612] = 128;
    exp_47_ram[2613] = 0;
    exp_47_ram[2614] = 199;
    exp_47_ram[2615] = 79;
    exp_47_ram[2616] = 0;
    exp_47_ram[2617] = 71;
    exp_47_ram[2618] = 143;
    exp_47_ram[2619] = 0;
    exp_47_ram[2620] = 199;
    exp_47_ram[2621] = 207;
    exp_47_ram[2622] = 193;
    exp_47_ram[2623] = 129;
    exp_47_ram[2624] = 1;
    exp_47_ram[2625] = 0;
    exp_47_ram[2626] = 1;
    exp_47_ram[2627] = 17;
    exp_47_ram[2628] = 129;
    exp_47_ram[2629] = 33;
    exp_47_ram[2630] = 49;
    exp_47_ram[2631] = 65;
    exp_47_ram[2632] = 81;
    exp_47_ram[2633] = 97;
    exp_47_ram[2634] = 113;
    exp_47_ram[2635] = 1;
    exp_47_ram[2636] = 0;
    exp_47_ram[2637] = 7;
    exp_47_ram[2638] = 143;
    exp_47_ram[2639] = 128;
    exp_47_ram[2640] = 244;
    exp_47_ram[2641] = 128;
    exp_47_ram[2642] = 244;
    exp_47_ram[2643] = 16;
    exp_47_ram[2644] = 244;
    exp_47_ram[2645] = 16;
    exp_47_ram[2646] = 244;
    exp_47_ram[2647] = 80;
    exp_47_ram[2648] = 244;
    exp_47_ram[2649] = 4;
    exp_47_ram[2650] = 240;
    exp_47_ram[2651] = 244;
    exp_47_ram[2652] = 196;
    exp_47_ram[2653] = 7;
    exp_47_ram[2654] = 79;
    exp_47_ram[2655] = 5;
    exp_47_ram[2656] = 5;
    exp_47_ram[2657] = 228;
    exp_47_ram[2658] = 244;
    exp_47_ram[2659] = 196;
    exp_47_ram[2660] = 7;
    exp_47_ram[2661] = 223;
    exp_47_ram[2662] = 5;
    exp_47_ram[2663] = 0;
    exp_47_ram[2664] = 135;
    exp_47_ram[2665] = 7;
    exp_47_ram[2666] = 15;
    exp_47_ram[2667] = 5;
    exp_47_ram[2668] = 7;
    exp_47_ram[2669] = 0;
    exp_47_ram[2670] = 135;
    exp_47_ram[2671] = 79;
    exp_47_ram[2672] = 0;
    exp_47_ram[2673] = 4;
    exp_47_ram[2674] = 7;
    exp_47_ram[2675] = 207;
    exp_47_ram[2676] = 5;
    exp_47_ram[2677] = 7;
    exp_47_ram[2678] = 159;
    exp_47_ram[2679] = 5;
    exp_47_ram[2680] = 0;
    exp_47_ram[2681] = 71;
    exp_47_ram[2682] = 7;
    exp_47_ram[2683] = 207;
    exp_47_ram[2684] = 5;
    exp_47_ram[2685] = 7;
    exp_47_ram[2686] = 0;
    exp_47_ram[2687] = 7;
    exp_47_ram[2688] = 15;
    exp_47_ram[2689] = 192;
    exp_47_ram[2690] = 4;
    exp_47_ram[2691] = 7;
    exp_47_ram[2692] = 79;
    exp_47_ram[2693] = 5;
    exp_47_ram[2694] = 7;
    exp_47_ram[2695] = 95;
    exp_47_ram[2696] = 5;
    exp_47_ram[2697] = 0;
    exp_47_ram[2698] = 135;
    exp_47_ram[2699] = 7;
    exp_47_ram[2700] = 143;
    exp_47_ram[2701] = 5;
    exp_47_ram[2702] = 7;
    exp_47_ram[2703] = 0;
    exp_47_ram[2704] = 199;
    exp_47_ram[2705] = 207;
    exp_47_ram[2706] = 128;
    exp_47_ram[2707] = 4;
    exp_47_ram[2708] = 7;
    exp_47_ram[2709] = 207;
    exp_47_ram[2710] = 5;
    exp_47_ram[2711] = 0;
    exp_47_ram[2712] = 71;
    exp_47_ram[2713] = 7;
    exp_47_ram[2714] = 15;
    exp_47_ram[2715] = 5;
    exp_47_ram[2716] = 7;
    exp_47_ram[2717] = 0;
    exp_47_ram[2718] = 71;
    exp_47_ram[2719] = 79;
    exp_47_ram[2720] = 0;
    exp_47_ram[2721] = 128;
    exp_47_ram[2722] = 244;
    exp_47_ram[2723] = 128;
    exp_47_ram[2724] = 244;
    exp_47_ram[2725] = 16;
    exp_47_ram[2726] = 244;
    exp_47_ram[2727] = 16;
    exp_47_ram[2728] = 244;
    exp_47_ram[2729] = 80;
    exp_47_ram[2730] = 244;
    exp_47_ram[2731] = 4;
    exp_47_ram[2732] = 16;
    exp_47_ram[2733] = 244;
    exp_47_ram[2734] = 196;
    exp_47_ram[2735] = 7;
    exp_47_ram[2736] = 223;
    exp_47_ram[2737] = 5;
    exp_47_ram[2738] = 5;
    exp_47_ram[2739] = 228;
    exp_47_ram[2740] = 244;
    exp_47_ram[2741] = 196;
    exp_47_ram[2742] = 7;
    exp_47_ram[2743] = 95;
    exp_47_ram[2744] = 5;
    exp_47_ram[2745] = 0;
    exp_47_ram[2746] = 135;
    exp_47_ram[2747] = 7;
    exp_47_ram[2748] = 143;
    exp_47_ram[2749] = 5;
    exp_47_ram[2750] = 7;
    exp_47_ram[2751] = 0;
    exp_47_ram[2752] = 135;
    exp_47_ram[2753] = 207;
    exp_47_ram[2754] = 128;
    exp_47_ram[2755] = 4;
    exp_47_ram[2756] = 7;
    exp_47_ram[2757] = 79;
    exp_47_ram[2758] = 5;
    exp_47_ram[2759] = 7;
    exp_47_ram[2760] = 31;
    exp_47_ram[2761] = 5;
    exp_47_ram[2762] = 0;
    exp_47_ram[2763] = 71;
    exp_47_ram[2764] = 7;
    exp_47_ram[2765] = 79;
    exp_47_ram[2766] = 5;
    exp_47_ram[2767] = 7;
    exp_47_ram[2768] = 0;
    exp_47_ram[2769] = 199;
    exp_47_ram[2770] = 143;
    exp_47_ram[2771] = 64;
    exp_47_ram[2772] = 4;
    exp_47_ram[2773] = 7;
    exp_47_ram[2774] = 207;
    exp_47_ram[2775] = 5;
    exp_47_ram[2776] = 7;
    exp_47_ram[2777] = 223;
    exp_47_ram[2778] = 5;
    exp_47_ram[2779] = 0;
    exp_47_ram[2780] = 135;
    exp_47_ram[2781] = 7;
    exp_47_ram[2782] = 15;
    exp_47_ram[2783] = 5;
    exp_47_ram[2784] = 7;
    exp_47_ram[2785] = 0;
    exp_47_ram[2786] = 7;
    exp_47_ram[2787] = 79;
    exp_47_ram[2788] = 0;
    exp_47_ram[2789] = 4;
    exp_47_ram[2790] = 7;
    exp_47_ram[2791] = 79;
    exp_47_ram[2792] = 5;
    exp_47_ram[2793] = 0;
    exp_47_ram[2794] = 71;
    exp_47_ram[2795] = 7;
    exp_47_ram[2796] = 143;
    exp_47_ram[2797] = 5;
    exp_47_ram[2798] = 7;
    exp_47_ram[2799] = 0;
    exp_47_ram[2800] = 135;
    exp_47_ram[2801] = 207;
    exp_47_ram[2802] = 128;
    exp_47_ram[2803] = 128;
    exp_47_ram[2804] = 244;
    exp_47_ram[2805] = 128;
    exp_47_ram[2806] = 244;
    exp_47_ram[2807] = 16;
    exp_47_ram[2808] = 244;
    exp_47_ram[2809] = 16;
    exp_47_ram[2810] = 244;
    exp_47_ram[2811] = 80;
    exp_47_ram[2812] = 244;
    exp_47_ram[2813] = 4;
    exp_47_ram[2814] = 4;
    exp_47_ram[2815] = 196;
    exp_47_ram[2816] = 7;
    exp_47_ram[2817] = 159;
    exp_47_ram[2818] = 5;
    exp_47_ram[2819] = 5;
    exp_47_ram[2820] = 228;
    exp_47_ram[2821] = 244;
    exp_47_ram[2822] = 196;
    exp_47_ram[2823] = 7;
    exp_47_ram[2824] = 31;
    exp_47_ram[2825] = 5;
    exp_47_ram[2826] = 0;
    exp_47_ram[2827] = 71;
    exp_47_ram[2828] = 7;
    exp_47_ram[2829] = 79;
    exp_47_ram[2830] = 5;
    exp_47_ram[2831] = 7;
    exp_47_ram[2832] = 0;
    exp_47_ram[2833] = 7;
    exp_47_ram[2834] = 143;
    exp_47_ram[2835] = 64;
    exp_47_ram[2836] = 4;
    exp_47_ram[2837] = 7;
    exp_47_ram[2838] = 31;
    exp_47_ram[2839] = 5;
    exp_47_ram[2840] = 7;
    exp_47_ram[2841] = 223;
    exp_47_ram[2842] = 5;
    exp_47_ram[2843] = 0;
    exp_47_ram[2844] = 135;
    exp_47_ram[2845] = 7;
    exp_47_ram[2846] = 15;
    exp_47_ram[2847] = 5;
    exp_47_ram[2848] = 7;
    exp_47_ram[2849] = 0;
    exp_47_ram[2850] = 71;
    exp_47_ram[2851] = 79;
    exp_47_ram[2852] = 0;
    exp_47_ram[2853] = 4;
    exp_47_ram[2854] = 7;
    exp_47_ram[2855] = 159;
    exp_47_ram[2856] = 5;
    exp_47_ram[2857] = 7;
    exp_47_ram[2858] = 159;
    exp_47_ram[2859] = 5;
    exp_47_ram[2860] = 0;
    exp_47_ram[2861] = 71;
    exp_47_ram[2862] = 7;
    exp_47_ram[2863] = 207;
    exp_47_ram[2864] = 5;
    exp_47_ram[2865] = 7;
    exp_47_ram[2866] = 0;
    exp_47_ram[2867] = 199;
    exp_47_ram[2868] = 15;
    exp_47_ram[2869] = 192;
    exp_47_ram[2870] = 4;
    exp_47_ram[2871] = 7;
    exp_47_ram[2872] = 31;
    exp_47_ram[2873] = 5;
    exp_47_ram[2874] = 0;
    exp_47_ram[2875] = 135;
    exp_47_ram[2876] = 7;
    exp_47_ram[2877] = 79;
    exp_47_ram[2878] = 5;
    exp_47_ram[2879] = 7;
    exp_47_ram[2880] = 0;
    exp_47_ram[2881] = 71;
    exp_47_ram[2882] = 159;
    exp_47_ram[2883] = 64;
    exp_47_ram[2884] = 0;
    exp_47_ram[2885] = 199;
    exp_47_ram[2886] = 159;
    exp_47_ram[2887] = 128;
    exp_47_ram[2888] = 244;
    exp_47_ram[2889] = 32;
    exp_47_ram[2890] = 244;
    exp_47_ram[2891] = 208;
    exp_47_ram[2892] = 244;
    exp_47_ram[2893] = 4;
    exp_47_ram[2894] = 176;
    exp_47_ram[2895] = 244;
    exp_47_ram[2896] = 112;
    exp_47_ram[2897] = 244;
    exp_47_ram[2898] = 240;
    exp_47_ram[2899] = 244;
    exp_47_ram[2900] = 196;
    exp_47_ram[2901] = 7;
    exp_47_ram[2902] = 95;
    exp_47_ram[2903] = 5;
    exp_47_ram[2904] = 5;
    exp_47_ram[2905] = 228;
    exp_47_ram[2906] = 244;
    exp_47_ram[2907] = 4;
    exp_47_ram[2908] = 68;
    exp_47_ram[2909] = 7;
    exp_47_ram[2910] = 7;
    exp_47_ram[2911] = 207;
    exp_47_ram[2912] = 207;
    exp_47_ram[2913] = 164;
    exp_47_ram[2914] = 180;
    exp_47_ram[2915] = 4;
    exp_47_ram[2916] = 128;
    exp_47_ram[2917] = 0;
    exp_47_ram[2918] = 79;
    exp_47_ram[2919] = 5;
    exp_47_ram[2920] = 5;
    exp_47_ram[2921] = 132;
    exp_47_ram[2922] = 196;
    exp_47_ram[2923] = 7;
    exp_47_ram[2924] = 7;
    exp_47_ram[2925] = 143;
    exp_47_ram[2926] = 5;
    exp_47_ram[2927] = 5;
    exp_47_ram[2928] = 0;
    exp_47_ram[2929] = 7;
    exp_47_ram[2930] = 7;
    exp_47_ram[2931] = 143;
    exp_47_ram[2932] = 5;
    exp_47_ram[2933] = 5;
    exp_47_ram[2934] = 7;
    exp_47_ram[2935] = 7;
    exp_47_ram[2936] = 11;
    exp_47_ram[2937] = 11;
    exp_47_ram[2938] = 143;
    exp_47_ram[2939] = 5;
    exp_47_ram[2940] = 7;
    exp_47_ram[2941] = 0;
    exp_47_ram[2942] = 7;
    exp_47_ram[2943] = 7;
    exp_47_ram[2944] = 0;
    exp_47_ram[2945] = 132;
    exp_47_ram[2946] = 196;
    exp_47_ram[2947] = 70;
    exp_47_ram[2948] = 7;
    exp_47_ram[2949] = 197;
    exp_47_ram[2950] = 86;
    exp_47_ram[2951] = 245;
    exp_47_ram[2952] = 6;
    exp_47_ram[2953] = 228;
    exp_47_ram[2954] = 244;
    exp_47_ram[2955] = 0;
    exp_47_ram[2956] = 143;
    exp_47_ram[2957] = 5;
    exp_47_ram[2958] = 5;
    exp_47_ram[2959] = 228;
    exp_47_ram[2960] = 244;
    exp_47_ram[2961] = 4;
    exp_47_ram[2962] = 7;
    exp_47_ram[2963] = 95;
    exp_47_ram[2964] = 5;
    exp_47_ram[2965] = 7;
    exp_47_ram[2966] = 159;
    exp_47_ram[2967] = 68;
    exp_47_ram[2968] = 23;
    exp_47_ram[2969] = 244;
    exp_47_ram[2970] = 68;
    exp_47_ram[2971] = 144;
    exp_47_ram[2972] = 231;
    exp_47_ram[2973] = 128;
    exp_47_ram[2974] = 244;
    exp_47_ram[2975] = 144;
    exp_47_ram[2976] = 244;
    exp_47_ram[2977] = 144;
    exp_47_ram[2978] = 244;
    exp_47_ram[2979] = 16;
    exp_47_ram[2980] = 244;
    exp_47_ram[2981] = 176;
    exp_47_ram[2982] = 244;
    exp_47_ram[2983] = 112;
    exp_47_ram[2984] = 244;
    exp_47_ram[2985] = 16;
    exp_47_ram[2986] = 244;
    exp_47_ram[2987] = 196;
    exp_47_ram[2988] = 7;
    exp_47_ram[2989] = 159;
    exp_47_ram[2990] = 5;
    exp_47_ram[2991] = 5;
    exp_47_ram[2992] = 228;
    exp_47_ram[2993] = 244;
    exp_47_ram[2994] = 196;
    exp_47_ram[2995] = 7;
    exp_47_ram[2996] = 15;
    exp_47_ram[2997] = 5;
    exp_47_ram[2998] = 7;
    exp_47_ram[2999] = 95;
    exp_47_ram[3000] = 4;
    exp_47_ram[3001] = 7;
    exp_47_ram[3002] = 159;
    exp_47_ram[3003] = 5;
    exp_47_ram[3004] = 7;
    exp_47_ram[3005] = 223;
    exp_47_ram[3006] = 4;
    exp_47_ram[3007] = 68;
    exp_47_ram[3008] = 7;
    exp_47_ram[3009] = 7;
    exp_47_ram[3010] = 15;
    exp_47_ram[3011] = 0;
    exp_47_ram[3012] = 143;
    exp_47_ram[3013] = 5;
    exp_47_ram[3014] = 5;
    exp_47_ram[3015] = 228;
    exp_47_ram[3016] = 244;
    exp_47_ram[3017] = 4;
    exp_47_ram[3018] = 7;
    exp_47_ram[3019] = 95;
    exp_47_ram[3020] = 5;
    exp_47_ram[3021] = 7;
    exp_47_ram[3022] = 159;
    exp_47_ram[3023] = 15;
    exp_47_ram[3024] = 164;
    exp_47_ram[3025] = 180;
    exp_47_ram[3026] = 4;
    exp_47_ram[3027] = 128;
    exp_47_ram[3028] = 0;
    exp_47_ram[3029] = 143;
    exp_47_ram[3030] = 5;
    exp_47_ram[3031] = 5;
    exp_47_ram[3032] = 132;
    exp_47_ram[3033] = 196;
    exp_47_ram[3034] = 7;
    exp_47_ram[3035] = 7;
    exp_47_ram[3036] = 207;
    exp_47_ram[3037] = 5;
    exp_47_ram[3038] = 5;
    exp_47_ram[3039] = 0;
    exp_47_ram[3040] = 7;
    exp_47_ram[3041] = 7;
    exp_47_ram[3042] = 207;
    exp_47_ram[3043] = 5;
    exp_47_ram[3044] = 5;
    exp_47_ram[3045] = 7;
    exp_47_ram[3046] = 7;
    exp_47_ram[3047] = 10;
    exp_47_ram[3048] = 10;
    exp_47_ram[3049] = 207;
    exp_47_ram[3050] = 5;
    exp_47_ram[3051] = 7;
    exp_47_ram[3052] = 0;
    exp_47_ram[3053] = 7;
    exp_47_ram[3054] = 7;
    exp_47_ram[3055] = 0;
    exp_47_ram[3056] = 132;
    exp_47_ram[3057] = 196;
    exp_47_ram[3058] = 38;
    exp_47_ram[3059] = 7;
    exp_47_ram[3060] = 197;
    exp_47_ram[3061] = 54;
    exp_47_ram[3062] = 245;
    exp_47_ram[3063] = 6;
    exp_47_ram[3064] = 228;
    exp_47_ram[3065] = 244;
    exp_47_ram[3066] = 0;
    exp_47_ram[3067] = 207;
    exp_47_ram[3068] = 5;
    exp_47_ram[3069] = 5;
    exp_47_ram[3070] = 228;
    exp_47_ram[3071] = 244;
    exp_47_ram[3072] = 4;
    exp_47_ram[3073] = 7;
    exp_47_ram[3074] = 159;
    exp_47_ram[3075] = 5;
    exp_47_ram[3076] = 7;
    exp_47_ram[3077] = 223;
    exp_47_ram[3078] = 4;
    exp_47_ram[3079] = 23;
    exp_47_ram[3080] = 244;
    exp_47_ram[3081] = 4;
    exp_47_ram[3082] = 144;
    exp_47_ram[3083] = 231;
    exp_47_ram[3084] = 193;
    exp_47_ram[3085] = 129;
    exp_47_ram[3086] = 65;
    exp_47_ram[3087] = 1;
    exp_47_ram[3088] = 193;
    exp_47_ram[3089] = 129;
    exp_47_ram[3090] = 65;
    exp_47_ram[3091] = 1;
    exp_47_ram[3092] = 1;
    exp_47_ram[3093] = 0;
    exp_47_ram[3094] = 1;
    exp_47_ram[3095] = 17;
    exp_47_ram[3096] = 129;
    exp_47_ram[3097] = 1;
    exp_47_ram[3098] = 31;
    exp_47_ram[3099] = 223;
    exp_47_ram[3100] = 0;
    exp_47_ram[3101] = 193;
    exp_47_ram[3102] = 129;
    exp_47_ram[3103] = 1;
    exp_47_ram[3104] = 0;
    exp_47_ram[3105] = 5;
    exp_47_ram[3106] = 5;
    exp_47_ram[3107] = 181;
    exp_47_ram[3108] = 1;
    exp_47_ram[3109] = 183;
    exp_47_ram[3110] = 7;
    exp_47_ram[3111] = 5;
    exp_47_ram[3112] = 21;
    exp_47_ram[3113] = 245;
    exp_47_ram[3114] = 1;
    exp_47_ram[3115] = 0;
    exp_47_ram[3116] = 176;
    exp_47_ram[3117] = 245;
    exp_47_ram[3118] = 245;
    exp_47_ram[3119] = 223;
    exp_47_ram[3120] = 250;
    exp_47_ram[3121] = 0;
    exp_47_ram[3122] = 110;
    exp_47_ram[3123] = 84;
    exp_47_ram[3124] = 101;
    exp_47_ram[3125] = 117;
    exp_47_ram[3126] = 83;
    exp_47_ram[3127] = 0;
    exp_47_ram[3128] = 110;
    exp_47_ram[3129] = 77;
    exp_47_ram[3130] = 112;
    exp_47_ram[3131] = 121;
    exp_47_ram[3132] = 74;
    exp_47_ram[3133] = 117;
    exp_47_ram[3134] = 112;
    exp_47_ram[3135] = 78;
    exp_47_ram[3136] = 101;
    exp_47_ram[3137] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 65;
    exp_40_ram[32] = 1;
    exp_40_ram[33] = 32;
    exp_40_ram[34] = 0;
    exp_40_ram[35] = 8;
    exp_40_ram[36] = 135;
    exp_40_ram[37] = 8;
    exp_40_ram[38] = 133;
    exp_40_ram[39] = 131;
    exp_40_ram[40] = 148;
    exp_40_ram[41] = 22;
    exp_40_ram[42] = 134;
    exp_40_ram[43] = 246;
    exp_40_ram[44] = 7;
    exp_40_ram[45] = 120;
    exp_40_ram[46] = 7;
    exp_40_ram[47] = 55;
    exp_40_ram[48] = 23;
    exp_40_ram[49] = 85;
    exp_40_ram[50] = 134;
    exp_40_ram[51] = 198;
    exp_40_ram[52] = 5;
    exp_40_ram[53] = 135;
    exp_40_ram[54] = 6;
    exp_40_ram[55] = 12;
    exp_40_ram[56] = 149;
    exp_40_ram[57] = 215;
    exp_40_ram[58] = 24;
    exp_40_ram[59] = 101;
    exp_40_ram[60] = 147;
    exp_40_ram[61] = 88;
    exp_40_ram[62] = 214;
    exp_40_ram[63] = 22;
    exp_40_ram[64] = 86;
    exp_40_ram[65] = 87;
    exp_40_ram[66] = 247;
    exp_40_ram[67] = 133;
    exp_40_ram[68] = 5;
    exp_40_ram[69] = 23;
    exp_40_ram[70] = 103;
    exp_40_ram[71] = 254;
    exp_40_ram[72] = 135;
    exp_40_ram[73] = 133;
    exp_40_ram[74] = 232;
    exp_40_ram[75] = 246;
    exp_40_ram[76] = 133;
    exp_40_ram[77] = 135;
    exp_40_ram[78] = 135;
    exp_40_ram[79] = 247;
    exp_40_ram[80] = 19;
    exp_40_ram[81] = 83;
    exp_40_ram[82] = 215;
    exp_40_ram[83] = 23;
    exp_40_ram[84] = 99;
    exp_40_ram[85] = 6;
    exp_40_ram[86] = 134;
    exp_40_ram[87] = 124;
    exp_40_ram[88] = 3;
    exp_40_ram[89] = 134;
    exp_40_ram[90] = 102;
    exp_40_ram[91] = 116;
    exp_40_ram[92] = 134;
    exp_40_ram[93] = 21;
    exp_40_ram[94] = 101;
    exp_40_ram[95] = 5;
    exp_40_ram[96] = 0;
    exp_40_ram[97] = 5;
    exp_40_ram[98] = 7;
    exp_40_ram[99] = 108;
    exp_40_ram[100] = 7;
    exp_40_ram[101] = 240;
    exp_40_ram[102] = 22;
    exp_40_ram[103] = 7;
    exp_40_ram[104] = 88;
    exp_40_ram[105] = 7;
    exp_40_ram[106] = 112;
    exp_40_ram[107] = 7;
    exp_40_ram[108] = 116;
    exp_40_ram[109] = 5;
    exp_40_ram[110] = 87;
    exp_40_ram[111] = 134;
    exp_40_ram[112] = 199;
    exp_40_ram[113] = 6;
    exp_40_ram[114] = 7;
    exp_40_ram[115] = 6;
    exp_40_ram[116] = 22;
    exp_40_ram[117] = 135;
    exp_40_ram[118] = 5;
    exp_40_ram[119] = 88;
    exp_40_ram[120] = 22;
    exp_40_ram[121] = 86;
    exp_40_ram[122] = 87;
    exp_40_ram[123] = 246;
    exp_40_ram[124] = 215;
    exp_40_ram[125] = 150;
    exp_40_ram[126] = 231;
    exp_40_ram[127] = 14;
    exp_40_ram[128] = 133;
    exp_40_ram[129] = 126;
    exp_40_ram[130] = 7;
    exp_40_ram[131] = 133;
    exp_40_ram[132] = 104;
    exp_40_ram[133] = 118;
    exp_40_ram[134] = 133;
    exp_40_ram[135] = 7;
    exp_40_ram[136] = 7;
    exp_40_ram[137] = 119;
    exp_40_ram[138] = 19;
    exp_40_ram[139] = 83;
    exp_40_ram[140] = 87;
    exp_40_ram[141] = 151;
    exp_40_ram[142] = 227;
    exp_40_ram[143] = 6;
    exp_40_ram[144] = 6;
    exp_40_ram[145] = 124;
    exp_40_ram[146] = 3;
    exp_40_ram[147] = 6;
    exp_40_ram[148] = 102;
    exp_40_ram[149] = 116;
    exp_40_ram[150] = 6;
    exp_40_ram[151] = 21;
    exp_40_ram[152] = 101;
    exp_40_ram[153] = 128;
    exp_40_ram[154] = 7;
    exp_40_ram[155] = 5;
    exp_40_ram[156] = 100;
    exp_40_ram[157] = 5;
    exp_40_ram[158] = 240;
    exp_40_ram[159] = 24;
    exp_40_ram[160] = 213;
    exp_40_ram[161] = 147;
    exp_40_ram[162] = 151;
    exp_40_ram[163] = 215;
    exp_40_ram[164] = 88;
    exp_40_ram[165] = 102;
    exp_40_ram[166] = 119;
    exp_40_ram[167] = 23;
    exp_40_ram[168] = 215;
    exp_40_ram[169] = 85;
    exp_40_ram[170] = 85;
    exp_40_ram[171] = 23;
    exp_40_ram[172] = 103;
    exp_40_ram[173] = 134;
    exp_40_ram[174] = 5;
    exp_40_ram[175] = 126;
    exp_40_ram[176] = 7;
    exp_40_ram[177] = 5;
    exp_40_ram[178] = 104;
    exp_40_ram[179] = 118;
    exp_40_ram[180] = 5;
    exp_40_ram[181] = 7;
    exp_40_ram[182] = 6;
    exp_40_ram[183] = 247;
    exp_40_ram[184] = 22;
    exp_40_ram[185] = 86;
    exp_40_ram[186] = 214;
    exp_40_ram[187] = 23;
    exp_40_ram[188] = 133;
    exp_40_ram[189] = 103;
    exp_40_ram[190] = 135;
    exp_40_ram[191] = 254;
    exp_40_ram[192] = 135;
    exp_40_ram[193] = 135;
    exp_40_ram[194] = 232;
    exp_40_ram[195] = 246;
    exp_40_ram[196] = 135;
    exp_40_ram[197] = 135;
    exp_40_ram[198] = 149;
    exp_40_ram[199] = 135;
    exp_40_ram[200] = 229;
    exp_40_ram[201] = 240;
    exp_40_ram[202] = 230;
    exp_40_ram[203] = 7;
    exp_40_ram[204] = 244;
    exp_40_ram[205] = 7;
    exp_40_ram[206] = 53;
    exp_40_ram[207] = 149;
    exp_40_ram[208] = 23;
    exp_40_ram[209] = 213;
    exp_40_ram[210] = 7;
    exp_40_ram[211] = 7;
    exp_40_ram[212] = 71;
    exp_40_ram[213] = 5;
    exp_40_ram[214] = 7;
    exp_40_ram[215] = 5;
    exp_40_ram[216] = 22;
    exp_40_ram[217] = 5;
    exp_40_ram[218] = 238;
    exp_40_ram[219] = 181;
    exp_40_ram[220] = 69;
    exp_40_ram[221] = 240;
    exp_40_ram[222] = 7;
    exp_40_ram[223] = 5;
    exp_40_ram[224] = 224;
    exp_40_ram[225] = 5;
    exp_40_ram[226] = 240;
    exp_40_ram[227] = 88;
    exp_40_ram[228] = 150;
    exp_40_ram[229] = 104;
    exp_40_ram[230] = 222;
    exp_40_ram[231] = 94;
    exp_40_ram[232] = 118;
    exp_40_ram[233] = 151;
    exp_40_ram[234] = 215;
    exp_40_ram[235] = 19;
    exp_40_ram[236] = 102;
    exp_40_ram[237] = 23;
    exp_40_ram[238] = 215;
    exp_40_ram[239] = 87;
    exp_40_ram[240] = 94;
    exp_40_ram[241] = 150;
    exp_40_ram[242] = 231;
    exp_40_ram[243] = 143;
    exp_40_ram[244] = 5;
    exp_40_ram[245] = 126;
    exp_40_ram[246] = 7;
    exp_40_ram[247] = 5;
    exp_40_ram[248] = 104;
    exp_40_ram[249] = 118;
    exp_40_ram[250] = 5;
    exp_40_ram[251] = 7;
    exp_40_ram[252] = 7;
    exp_40_ram[253] = 118;
    exp_40_ram[254] = 87;
    exp_40_ram[255] = 150;
    exp_40_ram[256] = 142;
    exp_40_ram[257] = 23;
    exp_40_ram[258] = 215;
    exp_40_ram[259] = 231;
    exp_40_ram[260] = 6;
    exp_40_ram[261] = 254;
    exp_40_ram[262] = 135;
    exp_40_ram[263] = 6;
    exp_40_ram[264] = 232;
    exp_40_ram[265] = 246;
    exp_40_ram[266] = 6;
    exp_40_ram[267] = 135;
    exp_40_ram[268] = 21;
    exp_40_ram[269] = 14;
    exp_40_ram[270] = 101;
    exp_40_ram[271] = 134;
    exp_40_ram[272] = 120;
    exp_40_ram[273] = 86;
    exp_40_ram[274] = 118;
    exp_40_ram[275] = 83;
    exp_40_ram[276] = 135;
    exp_40_ram[277] = 14;
    exp_40_ram[278] = 6;
    exp_40_ram[279] = 87;
    exp_40_ram[280] = 8;
    exp_40_ram[281] = 8;
    exp_40_ram[282] = 7;
    exp_40_ram[283] = 6;
    exp_40_ram[284] = 116;
    exp_40_ram[285] = 6;
    exp_40_ram[286] = 86;
    exp_40_ram[287] = 134;
    exp_40_ram[288] = 230;
    exp_40_ram[289] = 156;
    exp_40_ram[290] = 7;
    exp_40_ram[291] = 135;
    exp_40_ram[292] = 119;
    exp_40_ram[293] = 23;
    exp_40_ram[294] = 126;
    exp_40_ram[295] = 152;
    exp_40_ram[296] = 7;
    exp_40_ram[297] = 5;
    exp_40_ram[298] = 254;
    exp_40_ram[299] = 5;
    exp_40_ram[300] = 240;
    exp_40_ram[301] = 5;
    exp_40_ram[302] = 5;
    exp_40_ram[303] = 240;
    exp_40_ram[304] = 7;
    exp_40_ram[305] = 7;
    exp_40_ram[306] = 216;
    exp_40_ram[307] = 120;
    exp_40_ram[308] = 7;
    exp_40_ram[309] = 3;
    exp_40_ram[310] = 120;
    exp_40_ram[311] = 213;
    exp_40_ram[312] = 14;
    exp_40_ram[313] = 213;
    exp_40_ram[314] = 119;
    exp_40_ram[315] = 14;
    exp_40_ram[316] = 245;
    exp_40_ram[317] = 214;
    exp_40_ram[318] = 26;
    exp_40_ram[319] = 238;
    exp_40_ram[320] = 138;
    exp_40_ram[321] = 5;
    exp_40_ram[322] = 128;
    exp_40_ram[323] = 150;
    exp_40_ram[324] = 110;
    exp_40_ram[325] = 152;
    exp_40_ram[326] = 16;
    exp_40_ram[327] = 231;
    exp_40_ram[328] = 183;
    exp_40_ram[329] = 150;
    exp_40_ram[330] = 102;
    exp_40_ram[331] = 12;
    exp_40_ram[332] = 156;
    exp_40_ram[333] = 20;
    exp_40_ram[334] = 208;
    exp_40_ram[335] = 0;
    exp_40_ram[336] = 5;
    exp_40_ram[337] = 128;
    exp_40_ram[338] = 5;
    exp_40_ram[339] = 138;
    exp_40_ram[340] = 133;
    exp_40_ram[341] = 128;
    exp_40_ram[342] = 86;
    exp_40_ram[343] = 2;
    exp_40_ram[344] = 128;
    exp_40_ram[345] = 108;
    exp_40_ram[346] = 146;
    exp_40_ram[347] = 104;
    exp_40_ram[348] = 102;
    exp_40_ram[349] = 5;
    exp_40_ram[350] = 128;
    exp_40_ram[351] = 5;
    exp_40_ram[352] = 128;
    exp_40_ram[353] = 152;
    exp_40_ram[354] = 240;
    exp_40_ram[355] = 232;
    exp_40_ram[356] = 240;
    exp_40_ram[357] = 142;
    exp_40_ram[358] = 158;
    exp_40_ram[359] = 7;
    exp_40_ram[360] = 240;
    exp_40_ram[361] = 1;
    exp_40_ram[362] = 36;
    exp_40_ram[363] = 38;
    exp_40_ram[364] = 4;
    exp_40_ram[365] = 2;
    exp_40_ram[366] = 0;
    exp_40_ram[367] = 7;
    exp_40_ram[368] = 7;
    exp_40_ram[369] = 7;
    exp_40_ram[370] = 192;
    exp_40_ram[371] = 7;
    exp_40_ram[372] = 135;
    exp_40_ram[373] = 5;
    exp_40_ram[374] = 87;
    exp_40_ram[375] = 20;
    exp_40_ram[376] = 32;
    exp_40_ram[377] = 5;
    exp_40_ram[378] = 151;
    exp_40_ram[379] = 36;
    exp_40_ram[380] = 23;
    exp_40_ram[381] = 215;
    exp_40_ram[382] = 102;
    exp_40_ram[383] = 133;
    exp_40_ram[384] = 1;
    exp_40_ram[385] = 128;
    exp_40_ram[386] = 7;
    exp_40_ram[387] = 23;
    exp_40_ram[388] = 4;
    exp_40_ram[389] = 240;
    exp_40_ram[390] = 7;
    exp_40_ram[391] = 7;
    exp_40_ram[392] = 240;
    exp_40_ram[393] = 1;
    exp_40_ram[394] = 46;
    exp_40_ram[395] = 44;
    exp_40_ram[396] = 42;
    exp_40_ram[397] = 40;
    exp_40_ram[398] = 38;
    exp_40_ram[399] = 36;
    exp_40_ram[400] = 103;
    exp_40_ram[401] = 140;
    exp_40_ram[402] = 4;
    exp_40_ram[403] = 137;
    exp_40_ram[404] = 132;
    exp_40_ram[405] = 132;
    exp_40_ram[406] = 133;
    exp_40_ram[407] = 0;
    exp_40_ram[408] = 9;
    exp_40_ram[409] = 10;
    exp_40_ram[410] = 10;
    exp_40_ram[411] = 7;
    exp_40_ram[412] = 196;
    exp_40_ram[413] = 7;
    exp_40_ram[414] = 7;
    exp_40_ram[415] = 84;
    exp_40_ram[416] = 7;
    exp_40_ram[417] = 66;
    exp_40_ram[418] = 4;
    exp_40_ram[419] = 135;
    exp_40_ram[420] = 132;
    exp_40_ram[421] = 84;
    exp_40_ram[422] = 21;
    exp_40_ram[423] = 228;
    exp_40_ram[424] = 23;
    exp_40_ram[425] = 32;
    exp_40_ram[426] = 36;
    exp_40_ram[427] = 149;
    exp_40_ram[428] = 26;
    exp_40_ram[429] = 213;
    exp_40_ram[430] = 103;
    exp_40_ram[431] = 36;
    exp_40_ram[432] = 41;
    exp_40_ram[433] = 41;
    exp_40_ram[434] = 42;
    exp_40_ram[435] = 133;
    exp_40_ram[436] = 5;
    exp_40_ram[437] = 1;
    exp_40_ram[438] = 128;
    exp_40_ram[439] = 0;
    exp_40_ram[440] = 9;
    exp_40_ram[441] = 240;
    exp_40_ram[442] = 133;
    exp_40_ram[443] = 20;
    exp_40_ram[444] = 7;
    exp_40_ram[445] = 240;
    exp_40_ram[446] = 7;
    exp_40_ram[447] = 220;
    exp_40_ram[448] = 134;
    exp_40_ram[449] = 5;
    exp_40_ram[450] = 5;
    exp_40_ram[451] = 0;
    exp_40_ram[452] = 101;
    exp_40_ram[453] = 6;
    exp_40_ram[454] = 52;
    exp_40_ram[455] = 5;
    exp_40_ram[456] = 5;
    exp_40_ram[457] = 6;
    exp_40_ram[458] = 0;
    exp_40_ram[459] = 228;
    exp_40_ram[460] = 137;
    exp_40_ram[461] = 7;
    exp_40_ram[462] = 7;
    exp_40_ram[463] = 5;
    exp_40_ram[464] = 84;
    exp_40_ram[465] = 7;
    exp_40_ram[466] = 66;
    exp_40_ram[467] = 135;
    exp_40_ram[468] = 21;
    exp_40_ram[469] = 9;
    exp_40_ram[470] = 9;
    exp_40_ram[471] = 89;
    exp_40_ram[472] = 101;
    exp_40_ram[473] = 23;
    exp_40_ram[474] = 7;
    exp_40_ram[475] = 7;
    exp_40_ram[476] = 245;
    exp_40_ram[477] = 247;
    exp_40_ram[478] = 0;
    exp_40_ram[479] = 247;
    exp_40_ram[480] = 6;
    exp_40_ram[481] = 10;
    exp_40_ram[482] = 135;
    exp_40_ram[483] = 55;
    exp_40_ram[484] = 133;
    exp_40_ram[485] = 7;
    exp_40_ram[486] = 7;
    exp_40_ram[487] = 247;
    exp_40_ram[488] = 12;
    exp_40_ram[489] = 7;
    exp_40_ram[490] = 7;
    exp_40_ram[491] = 10;
    exp_40_ram[492] = 245;
    exp_40_ram[493] = 10;
    exp_40_ram[494] = 215;
    exp_40_ram[495] = 149;
    exp_40_ram[496] = 103;
    exp_40_ram[497] = 212;
    exp_40_ram[498] = 240;
    exp_40_ram[499] = 133;
    exp_40_ram[500] = 21;
    exp_40_ram[501] = 7;
    exp_40_ram[502] = 240;
    exp_40_ram[503] = 4;
    exp_40_ram[504] = 7;
    exp_40_ram[505] = 10;
    exp_40_ram[506] = 240;
    exp_40_ram[507] = 6;
    exp_40_ram[508] = 5;
    exp_40_ram[509] = 246;
    exp_40_ram[510] = 132;
    exp_40_ram[511] = 5;
    exp_40_ram[512] = 213;
    exp_40_ram[513] = 22;
    exp_40_ram[514] = 150;
    exp_40_ram[515] = 128;
    exp_40_ram[516] = 64;
    exp_40_ram[517] = 198;
    exp_40_ram[518] = 134;
    exp_40_ram[519] = 5;
    exp_40_ram[520] = 5;
    exp_40_ram[521] = 12;
    exp_40_ram[522] = 6;
    exp_40_ram[523] = 122;
    exp_40_ram[524] = 88;
    exp_40_ram[525] = 22;
    exp_40_ram[526] = 150;
    exp_40_ram[527] = 106;
    exp_40_ram[528] = 5;
    exp_40_ram[529] = 230;
    exp_40_ram[530] = 133;
    exp_40_ram[531] = 101;
    exp_40_ram[532] = 214;
    exp_40_ram[533] = 86;
    exp_40_ram[534] = 150;
    exp_40_ram[535] = 128;
    exp_40_ram[536] = 130;
    exp_40_ram[537] = 240;
    exp_40_ram[538] = 133;
    exp_40_ram[539] = 128;
    exp_40_ram[540] = 5;
    exp_40_ram[541] = 72;
    exp_40_ram[542] = 5;
    exp_40_ram[543] = 240;
    exp_40_ram[544] = 5;
    exp_40_ram[545] = 130;
    exp_40_ram[546] = 240;
    exp_40_ram[547] = 5;
    exp_40_ram[548] = 128;
    exp_40_ram[549] = 130;
    exp_40_ram[550] = 202;
    exp_40_ram[551] = 76;
    exp_40_ram[552] = 240;
    exp_40_ram[553] = 133;
    exp_40_ram[554] = 128;
    exp_40_ram[555] = 5;
    exp_40_ram[556] = 88;
    exp_40_ram[557] = 5;
    exp_40_ram[558] = 240;
    exp_40_ram[559] = 5;
    exp_40_ram[560] = 128;
    exp_40_ram[561] = 0;
    exp_40_ram[562] = 7;
    exp_40_ram[563] = 135;
    exp_40_ram[564] = 76;
    exp_40_ram[565] = 5;
    exp_40_ram[566] = 7;
    exp_40_ram[567] = 213;
    exp_40_ram[568] = 5;
    exp_40_ram[569] = 128;
    exp_40_ram[570] = 215;
    exp_40_ram[571] = 85;
    exp_40_ram[572] = 149;
    exp_40_ram[573] = 101;
    exp_40_ram[574] = 240;
    exp_40_ram[575] = 0;
    exp_40_ram[576] = 7;
    exp_40_ram[577] = 135;
    exp_40_ram[578] = 76;
    exp_40_ram[579] = 5;
    exp_40_ram[580] = 7;
    exp_40_ram[581] = 21;
    exp_40_ram[582] = 5;
    exp_40_ram[583] = 128;
    exp_40_ram[584] = 23;
    exp_40_ram[585] = 149;
    exp_40_ram[586] = 85;
    exp_40_ram[587] = 229;
    exp_40_ram[588] = 240;
    exp_40_ram[589] = 7;
    exp_40_ram[590] = 122;
    exp_40_ram[591] = 7;
    exp_40_ram[592] = 183;
    exp_40_ram[593] = 151;
    exp_40_ram[594] = 23;
    exp_40_ram[595] = 6;
    exp_40_ram[596] = 134;
    exp_40_ram[597] = 85;
    exp_40_ram[598] = 7;
    exp_40_ram[599] = 133;
    exp_40_ram[600] = 69;
    exp_40_ram[601] = 133;
    exp_40_ram[602] = 128;
    exp_40_ram[603] = 7;
    exp_40_ram[604] = 7;
    exp_40_ram[605] = 106;
    exp_40_ram[606] = 7;
    exp_40_ram[607] = 240;
    exp_40_ram[608] = 116;
    exp_40_ram[609] = 116;
    exp_40_ram[610] = 0;
    exp_40_ram[611] = 108;
    exp_40_ram[612] = 101;
    exp_40_ram[613] = 0;
    exp_40_ram[614] = 32;
    exp_40_ram[615] = 108;
    exp_40_ram[616] = 32;
    exp_40_ram[617] = 108;
    exp_40_ram[618] = 101;
    exp_40_ram[619] = 32;
    exp_40_ram[620] = 108;
    exp_40_ram[621] = 32;
    exp_40_ram[622] = 108;
    exp_40_ram[623] = 97;
    exp_40_ram[624] = 0;
    exp_40_ram[625] = 116;
    exp_40_ram[626] = 97;
    exp_40_ram[627] = 46;
    exp_40_ram[628] = 108;
    exp_40_ram[629] = 122;
    exp_40_ram[630] = 101;
    exp_40_ram[631] = 112;
    exp_40_ram[632] = 0;
    exp_40_ram[633] = 116;
    exp_40_ram[634] = 112;
    exp_40_ram[635] = 0;
    exp_40_ram[636] = 116;
    exp_40_ram[637] = 109;
    exp_40_ram[638] = 46;
    exp_40_ram[639] = 101;
    exp_40_ram[640] = 114;
    exp_40_ram[641] = 0;
    exp_40_ram[642] = 32;
    exp_40_ram[643] = 108;
    exp_40_ram[644] = 116;
    exp_40_ram[645] = 114;
    exp_40_ram[646] = 0;
    exp_40_ram[647] = 32;
    exp_40_ram[648] = 108;
    exp_40_ram[649] = 116;
    exp_40_ram[650] = 112;
    exp_40_ram[651] = 46;
    exp_40_ram[652] = 115;
    exp_40_ram[653] = 0;
    exp_40_ram[654] = 115;
    exp_40_ram[655] = 115;
    exp_40_ram[656] = 0;
    exp_40_ram[657] = 115;
    exp_40_ram[658] = 115;
    exp_40_ram[659] = 0;
    exp_40_ram[660] = 115;
    exp_40_ram[661] = 100;
    exp_40_ram[662] = 0;
    exp_40_ram[663] = 115;
    exp_40_ram[664] = 115;
    exp_40_ram[665] = 0;
    exp_40_ram[666] = 116;
    exp_40_ram[667] = 114;
    exp_40_ram[668] = 46;
    exp_40_ram[669] = 115;
    exp_40_ram[670] = 115;
    exp_40_ram[671] = 0;
    exp_40_ram[672] = 100;
    exp_40_ram[673] = 115;
    exp_40_ram[674] = 107;
    exp_40_ram[675] = 107;
    exp_40_ram[676] = 97;
    exp_40_ram[677] = 0;
    exp_40_ram[678] = 115;
    exp_40_ram[679] = 115;
    exp_40_ram[680] = 0;
    exp_40_ram[681] = 116;
    exp_40_ram[682] = 104;
    exp_40_ram[683] = 46;
    exp_40_ram[684] = 116;
    exp_40_ram[685] = 110;
    exp_40_ram[686] = 0;
    exp_40_ram[687] = 115;
    exp_40_ram[688] = 102;
    exp_40_ram[689] = 115;
    exp_40_ram[690] = 49;
    exp_40_ram[691] = 102;
    exp_40_ram[692] = 115;
    exp_40_ram[693] = 97;
    exp_40_ram[694] = 102;
    exp_40_ram[695] = 115;
    exp_40_ram[696] = 50;
    exp_40_ram[697] = 51;
    exp_40_ram[698] = 0;
    exp_40_ram[699] = 116;
    exp_40_ram[700] = 114;
    exp_40_ram[701] = 0;
    exp_40_ram[702] = 50;
    exp_40_ram[703] = 0;
    exp_40_ram[704] = 51;
    exp_40_ram[705] = 52;
    exp_40_ram[706] = 101;
    exp_40_ram[707] = 116;
    exp_40_ram[708] = 0;
    exp_40_ram[709] = 50;
    exp_40_ram[710] = 0;
    exp_40_ram[711] = 98;
    exp_40_ram[712] = 0;
    exp_40_ram[713] = 99;
    exp_40_ram[714] = 0;
    exp_40_ram[715] = 100;
    exp_40_ram[716] = 0;
    exp_40_ram[717] = 116;
    exp_40_ram[718] = 110;
    exp_40_ram[719] = 0;
    exp_40_ram[720] = 105;
    exp_40_ram[721] = 46;
    exp_40_ram[722] = 104;
    exp_40_ram[723] = 101;
    exp_40_ram[724] = 55;
    exp_40_ram[725] = 58;
    exp_40_ram[726] = 48;
    exp_40_ram[727] = 48;
    exp_40_ram[728] = 0;
    exp_40_ram[729] = 104;
    exp_40_ram[730] = 101;
    exp_40_ram[731] = 55;
    exp_40_ram[732] = 58;
    exp_40_ram[733] = 48;
    exp_40_ram[734] = 48;
    exp_40_ram[735] = 0;
    exp_40_ram[736] = 32;
    exp_40_ram[737] = 108;
    exp_40_ram[738] = 32;
    exp_40_ram[739] = 108;
    exp_40_ram[740] = 32;
    exp_40_ram[741] = 108;
    exp_40_ram[742] = 104;
    exp_40_ram[743] = 101;
    exp_40_ram[744] = 55;
    exp_40_ram[745] = 58;
    exp_40_ram[746] = 48;
    exp_40_ram[747] = 48;
    exp_40_ram[748] = 0;
    exp_40_ram[749] = 48;
    exp_40_ram[750] = 105;
    exp_40_ram[751] = 49;
    exp_40_ram[752] = 105;
    exp_40_ram[753] = 50;
    exp_40_ram[754] = 105;
    exp_40_ram[755] = 1;
    exp_40_ram[756] = 3;
    exp_40_ram[757] = 4;
    exp_40_ram[758] = 4;
    exp_40_ram[759] = 5;
    exp_40_ram[760] = 5;
    exp_40_ram[761] = 5;
    exp_40_ram[762] = 5;
    exp_40_ram[763] = 6;
    exp_40_ram[764] = 6;
    exp_40_ram[765] = 6;
    exp_40_ram[766] = 6;
    exp_40_ram[767] = 6;
    exp_40_ram[768] = 6;
    exp_40_ram[769] = 6;
    exp_40_ram[770] = 6;
    exp_40_ram[771] = 7;
    exp_40_ram[772] = 7;
    exp_40_ram[773] = 7;
    exp_40_ram[774] = 7;
    exp_40_ram[775] = 7;
    exp_40_ram[776] = 7;
    exp_40_ram[777] = 7;
    exp_40_ram[778] = 7;
    exp_40_ram[779] = 7;
    exp_40_ram[780] = 7;
    exp_40_ram[781] = 7;
    exp_40_ram[782] = 7;
    exp_40_ram[783] = 7;
    exp_40_ram[784] = 7;
    exp_40_ram[785] = 7;
    exp_40_ram[786] = 7;
    exp_40_ram[787] = 8;
    exp_40_ram[788] = 8;
    exp_40_ram[789] = 8;
    exp_40_ram[790] = 8;
    exp_40_ram[791] = 8;
    exp_40_ram[792] = 8;
    exp_40_ram[793] = 8;
    exp_40_ram[794] = 8;
    exp_40_ram[795] = 8;
    exp_40_ram[796] = 8;
    exp_40_ram[797] = 8;
    exp_40_ram[798] = 8;
    exp_40_ram[799] = 8;
    exp_40_ram[800] = 8;
    exp_40_ram[801] = 8;
    exp_40_ram[802] = 8;
    exp_40_ram[803] = 8;
    exp_40_ram[804] = 8;
    exp_40_ram[805] = 8;
    exp_40_ram[806] = 8;
    exp_40_ram[807] = 8;
    exp_40_ram[808] = 8;
    exp_40_ram[809] = 8;
    exp_40_ram[810] = 8;
    exp_40_ram[811] = 8;
    exp_40_ram[812] = 8;
    exp_40_ram[813] = 8;
    exp_40_ram[814] = 8;
    exp_40_ram[815] = 8;
    exp_40_ram[816] = 8;
    exp_40_ram[817] = 8;
    exp_40_ram[818] = 8;
    exp_40_ram[819] = 7;
    exp_40_ram[820] = 5;
    exp_40_ram[821] = 135;
    exp_40_ram[822] = 71;
    exp_40_ram[823] = 20;
    exp_40_ram[824] = 128;
    exp_40_ram[825] = 5;
    exp_40_ram[826] = 160;
    exp_40_ram[827] = 240;
    exp_40_ram[828] = 1;
    exp_40_ram[829] = 55;
    exp_40_ram[830] = 36;
    exp_40_ram[831] = 164;
    exp_40_ram[832] = 38;
    exp_40_ram[833] = 5;
    exp_40_ram[834] = 240;
    exp_40_ram[835] = 7;
    exp_40_ram[836] = 32;
    exp_40_ram[837] = 32;
    exp_40_ram[838] = 36;
    exp_40_ram[839] = 5;
    exp_40_ram[840] = 1;
    exp_40_ram[841] = 128;
    exp_40_ram[842] = 103;
    exp_40_ram[843] = 247;
    exp_40_ram[844] = 6;
    exp_40_ram[845] = 152;
    exp_40_ram[846] = 135;
    exp_40_ram[847] = 131;
    exp_40_ram[848] = 8;
    exp_40_ram[849] = 0;
    exp_40_ram[850] = 40;
    exp_40_ram[851] = 7;
    exp_40_ram[852] = 134;
    exp_40_ram[853] = 168;
    exp_40_ram[854] = 40;
    exp_40_ram[855] = 170;
    exp_40_ram[856] = 40;
    exp_40_ram[857] = 172;
    exp_40_ram[858] = 40;
    exp_40_ram[859] = 174;
    exp_40_ram[860] = 8;
    exp_40_ram[861] = 106;
    exp_40_ram[862] = 119;
    exp_40_ram[863] = 118;
    exp_40_ram[864] = 6;
    exp_40_ram[865] = 133;
    exp_40_ram[866] = 6;
    exp_40_ram[867] = 8;
    exp_40_ram[868] = 96;
    exp_40_ram[869] = 118;
    exp_40_ram[870] = 119;
    exp_40_ram[871] = 134;
    exp_40_ram[872] = 133;
    exp_40_ram[873] = 7;
    exp_40_ram[874] = 16;
    exp_40_ram[875] = 128;
    exp_40_ram[876] = 136;
    exp_40_ram[877] = 40;
    exp_40_ram[878] = 136;
    exp_40_ram[879] = 135;
    exp_40_ram[880] = 32;
    exp_40_ram[881] = 240;
    exp_40_ram[882] = 135;
    exp_40_ram[883] = 72;
    exp_40_ram[884] = 135;
    exp_40_ram[885] = 135;
    exp_40_ram[886] = 0;
    exp_40_ram[887] = 240;
    exp_40_ram[888] = 7;
    exp_40_ram[889] = 199;
    exp_40_ram[890] = 30;
    exp_40_ram[891] = 134;
    exp_40_ram[892] = 199;
    exp_40_ram[893] = 28;
    exp_40_ram[894] = 199;
    exp_40_ram[895] = 18;
    exp_40_ram[896] = 128;
    exp_40_ram[897] = 135;
    exp_40_ram[898] = 240;
    exp_40_ram[899] = 134;
    exp_40_ram[900] = 135;
    exp_40_ram[901] = 133;
    exp_40_ram[902] = 143;
    exp_40_ram[903] = 240;
    exp_40_ram[904] = 128;
    exp_40_ram[905] = 128;
    exp_40_ram[906] = 103;
    exp_40_ram[907] = 247;
    exp_40_ram[908] = 144;
    exp_40_ram[909] = 6;
    exp_40_ram[910] = 134;
    exp_40_ram[911] = 134;
    exp_40_ram[912] = 6;
    exp_40_ram[913] = 167;
    exp_40_ram[914] = 39;
    exp_40_ram[915] = 142;
    exp_40_ram[916] = 71;
    exp_40_ram[917] = 199;
    exp_40_ram[918] = 132;
    exp_40_ram[919] = 134;
    exp_40_ram[920] = 133;
    exp_40_ram[921] = 128;
    exp_40_ram[922] = 135;
    exp_40_ram[923] = 199;
    exp_40_ram[924] = 119;
    exp_40_ram[925] = 247;
    exp_40_ram[926] = 158;
    exp_40_ram[927] = 5;
    exp_40_ram[928] = 133;
    exp_40_ram[929] = 240;
    exp_40_ram[930] = 5;
    exp_40_ram[931] = 133;
    exp_40_ram[932] = 240;
    exp_40_ram[933] = 5;
    exp_40_ram[934] = 128;
    exp_40_ram[935] = 7;
    exp_40_ram[936] = 5;
    exp_40_ram[937] = 135;
    exp_40_ram[938] = 71;
    exp_40_ram[939] = 20;
    exp_40_ram[940] = 128;
    exp_40_ram[941] = 5;
    exp_40_ram[942] = 240;
    exp_40_ram[943] = 7;
    exp_40_ram[944] = 148;
    exp_40_ram[945] = 128;
    exp_40_ram[946] = 7;
    exp_40_ram[947] = 0;
    exp_40_ram[948] = 135;
    exp_40_ram[949] = 240;
    exp_40_ram[950] = 7;
    exp_40_ram[951] = 6;
    exp_40_ram[952] = 150;
    exp_40_ram[953] = 5;
    exp_40_ram[954] = 0;
    exp_40_ram[955] = 133;
    exp_40_ram[956] = 71;
    exp_40_ram[957] = 135;
    exp_40_ram[958] = 20;
    exp_40_ram[959] = 128;
    exp_40_ram[960] = 1;
    exp_40_ram[961] = 36;
    exp_40_ram[962] = 34;
    exp_40_ram[963] = 4;
    exp_40_ram[964] = 38;
    exp_40_ram[965] = 132;
    exp_40_ram[966] = 240;
    exp_40_ram[967] = 7;
    exp_40_ram[968] = 7;
    exp_40_ram[969] = 150;
    exp_40_ram[970] = 5;
    exp_40_ram[971] = 0;
    exp_40_ram[972] = 133;
    exp_40_ram[973] = 70;
    exp_40_ram[974] = 135;
    exp_40_ram[975] = 148;
    exp_40_ram[976] = 32;
    exp_40_ram[977] = 36;
    exp_40_ram[978] = 36;
    exp_40_ram[979] = 1;
    exp_40_ram[980] = 128;
    exp_40_ram[981] = 1;
    exp_40_ram[982] = 36;
    exp_40_ram[983] = 34;
    exp_40_ram[984] = 4;
    exp_40_ram[985] = 38;
    exp_40_ram[986] = 132;
    exp_40_ram[987] = 240;
    exp_40_ram[988] = 7;
    exp_40_ram[989] = 7;
    exp_40_ram[990] = 22;
    exp_40_ram[991] = 5;
    exp_40_ram[992] = 0;
    exp_40_ram[993] = 133;
    exp_40_ram[994] = 71;
    exp_40_ram[995] = 135;
    exp_40_ram[996] = 20;
    exp_40_ram[997] = 32;
    exp_40_ram[998] = 36;
    exp_40_ram[999] = 36;
    exp_40_ram[1000] = 1;
    exp_40_ram[1001] = 128;
    exp_40_ram[1002] = 1;
    exp_40_ram[1003] = 44;
    exp_40_ram[1004] = 42;
    exp_40_ram[1005] = 40;
    exp_40_ram[1006] = 38;
    exp_40_ram[1007] = 46;
    exp_40_ram[1008] = 9;
    exp_40_ram[1009] = 132;
    exp_40_ram[1010] = 240;
    exp_40_ram[1011] = 9;
    exp_40_ram[1012] = 4;
    exp_40_ram[1013] = 8;
    exp_40_ram[1014] = 133;
    exp_40_ram[1015] = 240;
    exp_40_ram[1016] = 7;
    exp_40_ram[1017] = 134;
    exp_40_ram[1018] = 0;
    exp_40_ram[1019] = 135;
    exp_40_ram[1020] = 198;
    exp_40_ram[1021] = 71;
    exp_40_ram[1022] = 6;
    exp_40_ram[1023] = 135;
    exp_40_ram[1024] = 22;
    exp_40_ram[1025] = 32;
    exp_40_ram[1026] = 5;
    exp_40_ram[1027] = 36;
    exp_40_ram[1028] = 36;
    exp_40_ram[1029] = 41;
    exp_40_ram[1030] = 41;
    exp_40_ram[1031] = 1;
    exp_40_ram[1032] = 128;
    exp_40_ram[1033] = 4;
    exp_40_ram[1034] = 240;
    exp_40_ram[1035] = 1;
    exp_40_ram[1036] = 44;
    exp_40_ram[1037] = 42;
    exp_40_ram[1038] = 40;
    exp_40_ram[1039] = 38;
    exp_40_ram[1040] = 46;
    exp_40_ram[1041] = 9;
    exp_40_ram[1042] = 132;
    exp_40_ram[1043] = 240;
    exp_40_ram[1044] = 9;
    exp_40_ram[1045] = 4;
    exp_40_ram[1046] = 12;
    exp_40_ram[1047] = 133;
    exp_40_ram[1048] = 240;
    exp_40_ram[1049] = 7;
    exp_40_ram[1050] = 134;
    exp_40_ram[1051] = 0;
    exp_40_ram[1052] = 135;
    exp_40_ram[1053] = 198;
    exp_40_ram[1054] = 71;
    exp_40_ram[1055] = 10;
    exp_40_ram[1056] = 135;
    exp_40_ram[1057] = 22;
    exp_40_ram[1058] = 4;
    exp_40_ram[1059] = 240;
    exp_40_ram[1060] = 32;
    exp_40_ram[1061] = 5;
    exp_40_ram[1062] = 36;
    exp_40_ram[1063] = 36;
    exp_40_ram[1064] = 41;
    exp_40_ram[1065] = 41;
    exp_40_ram[1066] = 1;
    exp_40_ram[1067] = 128;
    exp_40_ram[1068] = 1;
    exp_40_ram[1069] = 36;
    exp_40_ram[1070] = 34;
    exp_40_ram[1071] = 32;
    exp_40_ram[1072] = 4;
    exp_40_ram[1073] = 38;
    exp_40_ram[1074] = 132;
    exp_40_ram[1075] = 240;
    exp_40_ram[1076] = 9;
    exp_40_ram[1077] = 14;
    exp_40_ram[1078] = 133;
    exp_40_ram[1079] = 240;
    exp_40_ram[1080] = 7;
    exp_40_ram[1081] = 7;
    exp_40_ram[1082] = 0;
    exp_40_ram[1083] = 134;
    exp_40_ram[1084] = 70;
    exp_40_ram[1085] = 198;
    exp_40_ram[1086] = 5;
    exp_40_ram[1087] = 12;
    exp_40_ram[1088] = 135;
    exp_40_ram[1089] = 20;
    exp_40_ram[1090] = 4;
    exp_40_ram[1091] = 240;
    exp_40_ram[1092] = 5;
    exp_40_ram[1093] = 32;
    exp_40_ram[1094] = 36;
    exp_40_ram[1095] = 36;
    exp_40_ram[1096] = 41;
    exp_40_ram[1097] = 1;
    exp_40_ram[1098] = 128;
    exp_40_ram[1099] = 1;
    exp_40_ram[1100] = 44;
    exp_40_ram[1101] = 42;
    exp_40_ram[1102] = 40;
    exp_40_ram[1103] = 38;
    exp_40_ram[1104] = 46;
    exp_40_ram[1105] = 9;
    exp_40_ram[1106] = 132;
    exp_40_ram[1107] = 240;
    exp_40_ram[1108] = 9;
    exp_40_ram[1109] = 4;
    exp_40_ram[1110] = 10;
    exp_40_ram[1111] = 133;
    exp_40_ram[1112] = 240;
    exp_40_ram[1113] = 7;
    exp_40_ram[1114] = 7;
    exp_40_ram[1115] = 133;
    exp_40_ram[1116] = 0;
    exp_40_ram[1117] = 6;
    exp_40_ram[1118] = 134;
    exp_40_ram[1119] = 70;
    exp_40_ram[1120] = 198;
    exp_40_ram[1121] = 24;
    exp_40_ram[1122] = 135;
    exp_40_ram[1123] = 20;
    exp_40_ram[1124] = 32;
    exp_40_ram[1125] = 36;
    exp_40_ram[1126] = 36;
    exp_40_ram[1127] = 41;
    exp_40_ram[1128] = 41;
    exp_40_ram[1129] = 1;
    exp_40_ram[1130] = 128;
    exp_40_ram[1131] = 5;
    exp_40_ram[1132] = 240;
    exp_40_ram[1133] = 4;
    exp_40_ram[1134] = 240;
    exp_40_ram[1135] = 119;
    exp_40_ram[1136] = 148;
    exp_40_ram[1137] = 1;
    exp_40_ram[1138] = 5;
    exp_40_ram[1139] = 36;
    exp_40_ram[1140] = 38;
    exp_40_ram[1141] = 4;
    exp_40_ram[1142] = 240;
    exp_40_ram[1143] = 7;
    exp_40_ram[1144] = 26;
    exp_40_ram[1145] = 5;
    exp_40_ram[1146] = 5;
    exp_40_ram[1147] = 240;
    exp_40_ram[1148] = 55;
    exp_40_ram[1149] = 32;
    exp_40_ram[1150] = 36;
    exp_40_ram[1151] = 133;
    exp_40_ram[1152] = 1;
    exp_40_ram[1153] = 128;
    exp_40_ram[1154] = 7;
    exp_40_ram[1155] = 133;
    exp_40_ram[1156] = 128;
    exp_40_ram[1157] = 135;
    exp_40_ram[1158] = 247;
    exp_40_ram[1159] = 130;
    exp_40_ram[1160] = 247;
    exp_40_ram[1161] = 6;
    exp_40_ram[1162] = 7;
    exp_40_ram[1163] = 12;
    exp_40_ram[1164] = 7;
    exp_40_ram[1165] = 7;
    exp_40_ram[1166] = 150;
    exp_40_ram[1167] = 1;
    exp_40_ram[1168] = 38;
    exp_40_ram[1169] = 240;
    exp_40_ram[1170] = 32;
    exp_40_ram[1171] = 55;
    exp_40_ram[1172] = 135;
    exp_40_ram[1173] = 133;
    exp_40_ram[1174] = 1;
    exp_40_ram[1175] = 128;
    exp_40_ram[1176] = 7;
    exp_40_ram[1177] = 133;
    exp_40_ram[1178] = 128;
    exp_40_ram[1179] = 7;
    exp_40_ram[1180] = 166;
    exp_40_ram[1181] = 166;
    exp_40_ram[1182] = 165;
    exp_40_ram[1183] = 5;
    exp_40_ram[1184] = 167;
    exp_40_ram[1185] = 229;
    exp_40_ram[1186] = 128;
    exp_40_ram[1187] = 7;
    exp_40_ram[1188] = 5;
    exp_40_ram[1189] = 183;
    exp_40_ram[1190] = 133;
    exp_40_ram[1191] = 1;
    exp_40_ram[1192] = 133;
    exp_40_ram[1193] = 38;
    exp_40_ram[1194] = 240;
    exp_40_ram[1195] = 32;
    exp_40_ram[1196] = 1;
    exp_40_ram[1197] = 128;
    exp_40_ram[1198] = 1;
    exp_40_ram[1199] = 34;
    exp_40_ram[1200] = 42;
    exp_40_ram[1201] = 42;
    exp_40_ram[1202] = 84;
    exp_40_ram[1203] = 44;
    exp_40_ram[1204] = 40;
    exp_40_ram[1205] = 38;
    exp_40_ram[1206] = 36;
    exp_40_ram[1207] = 46;
    exp_40_ram[1208] = 32;
    exp_40_ram[1209] = 10;
    exp_40_ram[1210] = 4;
    exp_40_ram[1211] = 9;
    exp_40_ram[1212] = 9;
    exp_40_ram[1213] = 138;
    exp_40_ram[1214] = 132;
    exp_40_ram[1215] = 146;
    exp_40_ram[1216] = 43;
    exp_40_ram[1217] = 90;
    exp_40_ram[1218] = 4;
    exp_40_ram[1219] = 138;
    exp_40_ram[1220] = 0;
    exp_40_ram[1221] = 133;
    exp_40_ram[1222] = 5;
    exp_40_ram[1223] = 240;
    exp_40_ram[1224] = 133;
    exp_40_ram[1225] = 240;
    exp_40_ram[1226] = 5;
    exp_40_ram[1227] = 55;
    exp_40_ram[1228] = 137;
    exp_40_ram[1229] = 9;
    exp_40_ram[1230] = 132;
    exp_40_ram[1231] = 240;
    exp_40_ram[1232] = 5;
    exp_40_ram[1233] = 240;
    exp_40_ram[1234] = 53;
    exp_40_ram[1235] = 133;
    exp_40_ram[1236] = 5;
    exp_40_ram[1237] = 240;
    exp_40_ram[1238] = 5;
    exp_40_ram[1239] = 55;
    exp_40_ram[1240] = 137;
    exp_40_ram[1241] = 9;
    exp_40_ram[1242] = 4;
    exp_40_ram[1243] = 240;
    exp_40_ram[1244] = 39;
    exp_40_ram[1245] = 38;
    exp_40_ram[1246] = 36;
    exp_40_ram[1247] = 23;
    exp_40_ram[1248] = 135;
    exp_40_ram[1249] = 151;
    exp_40_ram[1250] = 135;
    exp_40_ram[1251] = 23;
    exp_40_ram[1252] = 7;
    exp_40_ram[1253] = 151;
    exp_40_ram[1254] = 23;
    exp_40_ram[1255] = 37;
    exp_40_ram[1256] = 86;
    exp_40_ram[1257] = 214;
    exp_40_ram[1258] = 135;
    exp_40_ram[1259] = 134;
    exp_40_ram[1260] = 55;
    exp_40_ram[1261] = 135;
    exp_40_ram[1262] = 85;
    exp_40_ram[1263] = 214;
    exp_40_ram[1264] = 4;
    exp_40_ram[1265] = 183;
    exp_40_ram[1266] = 135;
    exp_40_ram[1267] = 133;
    exp_40_ram[1268] = 5;
    exp_40_ram[1269] = 4;
    exp_40_ram[1270] = 240;
    exp_40_ram[1271] = 133;
    exp_40_ram[1272] = 87;
    exp_40_ram[1273] = 180;
    exp_40_ram[1274] = 7;
    exp_40_ram[1275] = 133;
    exp_40_ram[1276] = 132;
    exp_40_ram[1277] = 4;
    exp_40_ram[1278] = 53;
    exp_40_ram[1279] = 32;
    exp_40_ram[1280] = 133;
    exp_40_ram[1281] = 36;
    exp_40_ram[1282] = 36;
    exp_40_ram[1283] = 41;
    exp_40_ram[1284] = 41;
    exp_40_ram[1285] = 42;
    exp_40_ram[1286] = 42;
    exp_40_ram[1287] = 43;
    exp_40_ram[1288] = 1;
    exp_40_ram[1289] = 128;
    exp_40_ram[1290] = 1;
    exp_40_ram[1291] = 38;
    exp_40_ram[1292] = 36;
    exp_40_ram[1293] = 4;
    exp_40_ram[1294] = 240;
    exp_40_ram[1295] = 55;
    exp_40_ram[1296] = 166;
    exp_40_ram[1297] = 6;
    exp_40_ram[1298] = 224;
    exp_40_ram[1299] = 55;
    exp_40_ram[1300] = 167;
    exp_40_ram[1301] = 5;
    exp_40_ram[1302] = 6;
    exp_40_ram[1303] = 32;
    exp_40_ram[1304] = 34;
    exp_40_ram[1305] = 32;
    exp_40_ram[1306] = 36;
    exp_40_ram[1307] = 5;
    exp_40_ram[1308] = 1;
    exp_40_ram[1309] = 128;
    exp_40_ram[1310] = 1;
    exp_40_ram[1311] = 38;
    exp_40_ram[1312] = 36;
    exp_40_ram[1313] = 34;
    exp_40_ram[1314] = 32;
    exp_40_ram[1315] = 4;
    exp_40_ram[1316] = 132;
    exp_40_ram[1317] = 240;
    exp_40_ram[1318] = 55;
    exp_40_ram[1319] = 166;
    exp_40_ram[1320] = 6;
    exp_40_ram[1321] = 57;
    exp_40_ram[1322] = 224;
    exp_40_ram[1323] = 133;
    exp_40_ram[1324] = 180;
    exp_40_ram[1325] = 4;
    exp_40_ram[1326] = 9;
    exp_40_ram[1327] = 4;
    exp_40_ram[1328] = 34;
    exp_40_ram[1329] = 32;
    exp_40_ram[1330] = 36;
    exp_40_ram[1331] = 32;
    exp_40_ram[1332] = 36;
    exp_40_ram[1333] = 41;
    exp_40_ram[1334] = 1;
    exp_40_ram[1335] = 128;
    exp_40_ram[1336] = 1;
    exp_40_ram[1337] = 53;
    exp_40_ram[1338] = 34;
    exp_40_ram[1339] = 6;
    exp_40_ram[1340] = 4;
    exp_40_ram[1341] = 133;
    exp_40_ram[1342] = 5;
    exp_40_ram[1343] = 38;
    exp_40_ram[1344] = 36;
    exp_40_ram[1345] = 32;
    exp_40_ram[1346] = 46;
    exp_40_ram[1347] = 44;
    exp_40_ram[1348] = 240;
    exp_40_ram[1349] = 53;
    exp_40_ram[1350] = 6;
    exp_40_ram[1351] = 133;
    exp_40_ram[1352] = 5;
    exp_40_ram[1353] = 240;
    exp_40_ram[1354] = 167;
    exp_40_ram[1355] = 57;
    exp_40_ram[1356] = 132;
    exp_40_ram[1357] = 149;
    exp_40_ram[1358] = 133;
    exp_40_ram[1359] = 7;
    exp_40_ram[1360] = 9;
    exp_40_ram[1361] = 133;
    exp_40_ram[1362] = 6;
    exp_40_ram[1363] = 133;
    exp_40_ram[1364] = 240;
    exp_40_ram[1365] = 1;
    exp_40_ram[1366] = 167;
    exp_40_ram[1367] = 6;
    exp_40_ram[1368] = 5;
    exp_40_ram[1369] = 149;
    exp_40_ram[1370] = 133;
    exp_40_ram[1371] = 7;
    exp_40_ram[1372] = 133;
    exp_40_ram[1373] = 240;
    exp_40_ram[1374] = 3;
    exp_40_ram[1375] = 165;
    exp_40_ram[1376] = 5;
    exp_40_ram[1377] = 10;
    exp_40_ram[1378] = 16;
    exp_40_ram[1379] = 36;
    exp_40_ram[1380] = 39;
    exp_40_ram[1381] = 38;
    exp_40_ram[1382] = 5;
    exp_40_ram[1383] = 135;
    exp_40_ram[1384] = 4;
    exp_40_ram[1385] = 39;
    exp_40_ram[1386] = 5;
    exp_40_ram[1387] = 135;
    exp_40_ram[1388] = 4;
    exp_40_ram[1389] = 165;
    exp_40_ram[1390] = 16;
    exp_40_ram[1391] = 36;
    exp_40_ram[1392] = 39;
    exp_40_ram[1393] = 38;
    exp_40_ram[1394] = 6;
    exp_40_ram[1395] = 135;
    exp_40_ram[1396] = 5;
    exp_40_ram[1397] = 39;
    exp_40_ram[1398] = 5;
    exp_40_ram[1399] = 135;
    exp_40_ram[1400] = 6;
    exp_40_ram[1401] = 165;
    exp_40_ram[1402] = 16;
    exp_40_ram[1403] = 36;
    exp_40_ram[1404] = 39;
    exp_40_ram[1405] = 38;
    exp_40_ram[1406] = 8;
    exp_40_ram[1407] = 135;
    exp_40_ram[1408] = 7;
    exp_40_ram[1409] = 39;
    exp_40_ram[1410] = 5;
    exp_40_ram[1411] = 135;
    exp_40_ram[1412] = 7;
    exp_40_ram[1413] = 165;
    exp_40_ram[1414] = 16;
    exp_40_ram[1415] = 36;
    exp_40_ram[1416] = 39;
    exp_40_ram[1417] = 38;
    exp_40_ram[1418] = 9;
    exp_40_ram[1419] = 135;
    exp_40_ram[1420] = 8;
    exp_40_ram[1421] = 39;
    exp_40_ram[1422] = 5;
    exp_40_ram[1423] = 135;
    exp_40_ram[1424] = 9;
    exp_40_ram[1425] = 165;
    exp_40_ram[1426] = 5;
    exp_40_ram[1427] = 16;
    exp_40_ram[1428] = 36;
    exp_40_ram[1429] = 38;
    exp_40_ram[1430] = 39;
    exp_40_ram[1431] = 37;
    exp_40_ram[1432] = 5;
    exp_40_ram[1433] = 135;
    exp_40_ram[1434] = 10;
    exp_40_ram[1435] = 16;
    exp_40_ram[1436] = 36;
    exp_40_ram[1437] = 38;
    exp_40_ram[1438] = 39;
    exp_40_ram[1439] = 37;
    exp_40_ram[1440] = 5;
    exp_40_ram[1441] = 135;
    exp_40_ram[1442] = 10;
    exp_40_ram[1443] = 16;
    exp_40_ram[1444] = 36;
    exp_40_ram[1445] = 39;
    exp_40_ram[1446] = 38;
    exp_40_ram[1447] = 32;
    exp_40_ram[1448] = 135;
    exp_40_ram[1449] = 11;
    exp_40_ram[1450] = 39;
    exp_40_ram[1451] = 36;
    exp_40_ram[1452] = 41;
    exp_40_ram[1453] = 135;
    exp_40_ram[1454] = 11;
    exp_40_ram[1455] = 7;
    exp_40_ram[1456] = 28;
    exp_40_ram[1457] = 36;
    exp_40_ram[1458] = 42;
    exp_40_ram[1459] = 133;
    exp_40_ram[1460] = 41;
    exp_40_ram[1461] = 1;
    exp_40_ram[1462] = 128;
    exp_40_ram[1463] = 1;
    exp_40_ram[1464] = 32;
    exp_40_ram[1465] = 91;
    exp_40_ram[1466] = 44;
    exp_40_ram[1467] = 42;
    exp_40_ram[1468] = 40;
    exp_40_ram[1469] = 38;
    exp_40_ram[1470] = 34;
    exp_40_ram[1471] = 46;
    exp_40_ram[1472] = 36;
    exp_40_ram[1473] = 46;
    exp_40_ram[1474] = 44;
    exp_40_ram[1475] = 42;
    exp_40_ram[1476] = 4;
    exp_40_ram[1477] = 132;
    exp_40_ram[1478] = 9;
    exp_40_ram[1479] = 9;
    exp_40_ram[1480] = 10;
    exp_40_ram[1481] = 11;
    exp_40_ram[1482] = 133;
    exp_40_ram[1483] = 240;
    exp_40_ram[1484] = 58;
    exp_40_ram[1485] = 10;
    exp_40_ram[1486] = 5;
    exp_40_ram[1487] = 5;
    exp_40_ram[1488] = 240;
    exp_40_ram[1489] = 135;
    exp_40_ram[1490] = 20;
    exp_40_ram[1491] = 224;
    exp_40_ram[1492] = 133;
    exp_40_ram[1493] = 183;
    exp_40_ram[1494] = 138;
    exp_40_ram[1495] = 4;
    exp_40_ram[1496] = 9;
    exp_40_ram[1497] = 137;
    exp_40_ram[1498] = 240;
    exp_40_ram[1499] = 92;
    exp_40_ram[1500] = 12;
    exp_40_ram[1501] = 10;
    exp_40_ram[1502] = 12;
    exp_40_ram[1503] = 133;
    exp_40_ram[1504] = 133;
    exp_40_ram[1505] = 240;
    exp_40_ram[1506] = 5;
    exp_40_ram[1507] = 139;
    exp_40_ram[1508] = 11;
    exp_40_ram[1509] = 140;
    exp_40_ram[1510] = 240;
    exp_40_ram[1511] = 20;
    exp_40_ram[1512] = 224;
    exp_40_ram[1513] = 133;
    exp_40_ram[1514] = 183;
    exp_40_ram[1515] = 138;
    exp_40_ram[1516] = 10;
    exp_40_ram[1517] = 4;
    exp_40_ram[1518] = 9;
    exp_40_ram[1519] = 240;
    exp_40_ram[1520] = 85;
    exp_40_ram[1521] = 133;
    exp_40_ram[1522] = 133;
    exp_40_ram[1523] = 16;
    exp_40_ram[1524] = 38;
    exp_40_ram[1525] = 4;
    exp_40_ram[1526] = 36;
    exp_40_ram[1527] = 10;
    exp_40_ram[1528] = 37;
    exp_40_ram[1529] = 21;
    exp_40_ram[1530] = 133;
    exp_40_ram[1531] = 16;
    exp_40_ram[1532] = 38;
    exp_40_ram[1533] = 9;
    exp_40_ram[1534] = 36;
    exp_40_ram[1535] = 37;
    exp_40_ram[1536] = 5;
    exp_40_ram[1537] = 137;
    exp_40_ram[1538] = 16;
    exp_40_ram[1539] = 135;
    exp_40_ram[1540] = 36;
    exp_40_ram[1541] = 38;
    exp_40_ram[1542] = 32;
    exp_40_ram[1543] = 34;
    exp_40_ram[1544] = 36;
    exp_40_ram[1545] = 40;
    exp_40_ram[1546] = 42;
    exp_40_ram[1547] = 133;
    exp_40_ram[1548] = 38;
    exp_40_ram[1549] = 5;
    exp_40_ram[1550] = 240;
    exp_40_ram[1551] = 44;
    exp_40_ram[1552] = 46;
    exp_40_ram[1553] = 32;
    exp_40_ram[1554] = 5;
    exp_40_ram[1555] = 36;
    exp_40_ram[1556] = 36;
    exp_40_ram[1557] = 41;
    exp_40_ram[1558] = 41;
    exp_40_ram[1559] = 42;
    exp_40_ram[1560] = 42;
    exp_40_ram[1561] = 43;
    exp_40_ram[1562] = 43;
    exp_40_ram[1563] = 44;
    exp_40_ram[1564] = 44;
    exp_40_ram[1565] = 1;
    exp_40_ram[1566] = 128;
    exp_40_ram[1567] = 1;
    exp_40_ram[1568] = 34;
    exp_40_ram[1569] = 42;
    exp_40_ram[1570] = 7;
    exp_40_ram[1571] = 42;
    exp_40_ram[1572] = 40;
    exp_40_ram[1573] = 36;
    exp_40_ram[1574] = 4;
    exp_40_ram[1575] = 10;
    exp_40_ram[1576] = 6;
    exp_40_ram[1577] = 9;
    exp_40_ram[1578] = 5;
    exp_40_ram[1579] = 5;
    exp_40_ram[1580] = 46;
    exp_40_ram[1581] = 36;
    exp_40_ram[1582] = 44;
    exp_40_ram[1583] = 38;
    exp_40_ram[1584] = 32;
    exp_40_ram[1585] = 34;
    exp_40_ram[1586] = 38;
    exp_40_ram[1587] = 46;
    exp_40_ram[1588] = 44;
    exp_40_ram[1589] = 44;
    exp_40_ram[1590] = 240;
    exp_40_ram[1591] = 5;
    exp_40_ram[1592] = 240;
    exp_40_ram[1593] = 134;
    exp_40_ram[1594] = 5;
    exp_40_ram[1595] = 5;
    exp_40_ram[1596] = 240;
    exp_40_ram[1597] = 39;
    exp_40_ram[1598] = 39;
    exp_40_ram[1599] = 6;
    exp_40_ram[1600] = 5;
    exp_40_ram[1601] = 135;
    exp_40_ram[1602] = 5;
    exp_40_ram[1603] = 34;
    exp_40_ram[1604] = 240;
    exp_40_ram[1605] = 5;
    exp_40_ram[1606] = 240;
    exp_40_ram[1607] = 7;
    exp_40_ram[1608] = 6;
    exp_40_ram[1609] = 9;
    exp_40_ram[1610] = 132;
    exp_40_ram[1611] = 5;
    exp_40_ram[1612] = 5;
    exp_40_ram[1613] = 38;
    exp_40_ram[1614] = 34;
    exp_40_ram[1615] = 36;
    exp_40_ram[1616] = 40;
    exp_40_ram[1617] = 32;
    exp_40_ram[1618] = 46;
    exp_40_ram[1619] = 240;
    exp_40_ram[1620] = 5;
    exp_40_ram[1621] = 240;
    exp_40_ram[1622] = 134;
    exp_40_ram[1623] = 5;
    exp_40_ram[1624] = 5;
    exp_40_ram[1625] = 240;
    exp_40_ram[1626] = 39;
    exp_40_ram[1627] = 39;
    exp_40_ram[1628] = 6;
    exp_40_ram[1629] = 5;
    exp_40_ram[1630] = 135;
    exp_40_ram[1631] = 5;
    exp_40_ram[1632] = 36;
    exp_40_ram[1633] = 240;
    exp_40_ram[1634] = 5;
    exp_40_ram[1635] = 240;
    exp_40_ram[1636] = 132;
    exp_40_ram[1637] = 10;
    exp_40_ram[1638] = 6;
    exp_40_ram[1639] = 5;
    exp_40_ram[1640] = 5;
    exp_40_ram[1641] = 240;
    exp_40_ram[1642] = 5;
    exp_40_ram[1643] = 240;
    exp_40_ram[1644] = 226;
    exp_40_ram[1645] = 7;
    exp_40_ram[1646] = 135;
    exp_40_ram[1647] = 148;
    exp_40_ram[1648] = 106;
    exp_40_ram[1649] = 5;
    exp_40_ram[1650] = 232;
    exp_40_ram[1651] = 20;
    exp_40_ram[1652] = 100;
    exp_40_ram[1653] = 5;
    exp_40_ram[1654] = 32;
    exp_40_ram[1655] = 36;
    exp_40_ram[1656] = 36;
    exp_40_ram[1657] = 41;
    exp_40_ram[1658] = 41;
    exp_40_ram[1659] = 42;
    exp_40_ram[1660] = 42;
    exp_40_ram[1661] = 1;
    exp_40_ram[1662] = 128;
    exp_40_ram[1663] = 1;
    exp_40_ram[1664] = 5;
    exp_40_ram[1665] = 40;
    exp_40_ram[1666] = 6;
    exp_40_ram[1667] = 9;
    exp_40_ram[1668] = 5;
    exp_40_ram[1669] = 46;
    exp_40_ram[1670] = 44;
    exp_40_ram[1671] = 42;
    exp_40_ram[1672] = 38;
    exp_40_ram[1673] = 240;
    exp_40_ram[1674] = 6;
    exp_40_ram[1675] = 5;
    exp_40_ram[1676] = 5;
    exp_40_ram[1677] = 41;
    exp_40_ram[1678] = 240;
    exp_40_ram[1679] = 5;
    exp_40_ram[1680] = 240;
    exp_40_ram[1681] = 4;
    exp_40_ram[1682] = 132;
    exp_40_ram[1683] = 88;
    exp_40_ram[1684] = 247;
    exp_40_ram[1685] = 135;
    exp_40_ram[1686] = 7;
    exp_40_ram[1687] = 183;
    exp_40_ram[1688] = 132;
    exp_40_ram[1689] = 132;
    exp_40_ram[1690] = 4;
    exp_40_ram[1691] = 133;
    exp_40_ram[1692] = 6;
    exp_40_ram[1693] = 5;
    exp_40_ram[1694] = 240;
    exp_40_ram[1695] = 6;
    exp_40_ram[1696] = 5;
    exp_40_ram[1697] = 5;
    exp_40_ram[1698] = 240;
    exp_40_ram[1699] = 88;
    exp_40_ram[1700] = 7;
    exp_40_ram[1701] = 32;
    exp_40_ram[1702] = 32;
    exp_40_ram[1703] = 5;
    exp_40_ram[1704] = 36;
    exp_40_ram[1705] = 41;
    exp_40_ram[1706] = 41;
    exp_40_ram[1707] = 133;
    exp_40_ram[1708] = 36;
    exp_40_ram[1709] = 1;
    exp_40_ram[1710] = 128;
    exp_40_ram[1711] = 136;
    exp_40_ram[1712] = 6;
    exp_40_ram[1713] = 5;
    exp_40_ram[1714] = 5;
    exp_40_ram[1715] = 240;
    exp_40_ram[1716] = 5;
    exp_40_ram[1717] = 240;
    exp_40_ram[1718] = 7;
    exp_40_ram[1719] = 6;
    exp_40_ram[1720] = 23;
    exp_40_ram[1721] = 135;
    exp_40_ram[1722] = 135;
    exp_40_ram[1723] = 183;
    exp_40_ram[1724] = 4;
    exp_40_ram[1725] = 132;
    exp_40_ram[1726] = 240;
    exp_40_ram[1727] = 130;
    exp_40_ram[1728] = 6;
    exp_40_ram[1729] = 5;
    exp_40_ram[1730] = 5;
    exp_40_ram[1731] = 240;
    exp_40_ram[1732] = 5;
    exp_40_ram[1733] = 240;
    exp_40_ram[1734] = 32;
    exp_40_ram[1735] = 240;
    exp_40_ram[1736] = 32;
    exp_40_ram[1737] = 240;
    exp_40_ram[1738] = 1;
    exp_40_ram[1739] = 134;
    exp_40_ram[1740] = 5;
    exp_40_ram[1741] = 5;
    exp_40_ram[1742] = 38;
    exp_40_ram[1743] = 240;
    exp_40_ram[1744] = 5;
    exp_40_ram[1745] = 6;
    exp_40_ram[1746] = 5;
    exp_40_ram[1747] = 240;
    exp_40_ram[1748] = 5;
    exp_40_ram[1749] = 240;
    exp_40_ram[1750] = 32;
    exp_40_ram[1751] = 1;
    exp_40_ram[1752] = 128;
    exp_40_ram[1753] = 37;
    exp_40_ram[1754] = 38;
    exp_40_ram[1755] = 1;
    exp_40_ram[1756] = 5;
    exp_40_ram[1757] = 46;
    exp_40_ram[1758] = 44;
    exp_40_ram[1759] = 240;
    exp_40_ram[1760] = 52;
    exp_40_ram[1761] = 5;
    exp_40_ram[1762] = 5;
    exp_40_ram[1763] = 6;
    exp_40_ram[1764] = 240;
    exp_40_ram[1765] = 32;
    exp_40_ram[1766] = 5;
    exp_40_ram[1767] = 36;
    exp_40_ram[1768] = 1;
    exp_40_ram[1769] = 128;
    exp_40_ram[1770] = 1;
    exp_40_ram[1771] = 34;
    exp_40_ram[1772] = 32;
    exp_40_ram[1773] = 36;
    exp_40_ram[1774] = 41;
    exp_40_ram[1775] = 38;
    exp_40_ram[1776] = 133;
    exp_40_ram[1777] = 5;
    exp_40_ram[1778] = 36;
    exp_40_ram[1779] = 46;
    exp_40_ram[1780] = 240;
    exp_40_ram[1781] = 6;
    exp_40_ram[1782] = 6;
    exp_40_ram[1783] = 22;
    exp_40_ram[1784] = 6;
    exp_40_ram[1785] = 5;
    exp_40_ram[1786] = 182;
    exp_40_ram[1787] = 6;
    exp_40_ram[1788] = 5;
    exp_40_ram[1789] = 240;
    exp_40_ram[1790] = 52;
    exp_40_ram[1791] = 5;
    exp_40_ram[1792] = 6;
    exp_40_ram[1793] = 5;
    exp_40_ram[1794] = 240;
    exp_40_ram[1795] = 5;
    exp_40_ram[1796] = 133;
    exp_40_ram[1797] = 240;
    exp_40_ram[1798] = 9;
    exp_40_ram[1799] = 160;
    exp_40_ram[1800] = 32;
    exp_40_ram[1801] = 5;
    exp_40_ram[1802] = 36;
    exp_40_ram[1803] = 36;
    exp_40_ram[1804] = 41;
    exp_40_ram[1805] = 41;
    exp_40_ram[1806] = 1;
    exp_40_ram[1807] = 128;
    exp_40_ram[1808] = 1;
    exp_40_ram[1809] = 38;
    exp_40_ram[1810] = 240;
    exp_40_ram[1811] = 32;
    exp_40_ram[1812] = 1;
    exp_40_ram[1813] = 240;
    exp_40_ram[1814] = 1;
    exp_40_ram[1815] = 46;
    exp_40_ram[1816] = 44;
    exp_40_ram[1817] = 4;
    exp_40_ram[1818] = 23;
    exp_40_ram[1819] = 133;
    exp_40_ram[1820] = 240;
    exp_40_ram[1821] = 7;
    exp_40_ram[1822] = 103;
    exp_40_ram[1823] = 7;
    exp_40_ram[1824] = 144;
    exp_40_ram[1825] = 129;
    exp_40_ram[1826] = 7;
    exp_40_ram[1827] = 133;
    exp_40_ram[1828] = 240;
    exp_40_ram[1829] = 7;
    exp_40_ram[1830] = 135;
    exp_40_ram[1831] = 7;
    exp_40_ram[1832] = 135;
    exp_40_ram[1833] = 23;
    exp_40_ram[1834] = 69;
    exp_40_ram[1835] = 6;
    exp_40_ram[1836] = 198;
    exp_40_ram[1837] = 6;
    exp_40_ram[1838] = 198;
    exp_40_ram[1839] = 7;
    exp_40_ram[1840] = 71;
    exp_40_ram[1841] = 128;
    exp_40_ram[1842] = 128;
    exp_40_ram[1843] = 129;
    exp_40_ram[1844] = 129;
    exp_40_ram[1845] = 7;
    exp_40_ram[1846] = 23;
    exp_40_ram[1847] = 133;
    exp_40_ram[1848] = 5;
    exp_40_ram[1849] = 240;
    exp_40_ram[1850] = 7;
    exp_40_ram[1851] = 138;
    exp_40_ram[1852] = 23;
    exp_40_ram[1853] = 133;
    exp_40_ram[1854] = 224;
    exp_40_ram[1855] = 0;
    exp_40_ram[1856] = 2;
    exp_40_ram[1857] = 7;
    exp_40_ram[1858] = 133;
    exp_40_ram[1859] = 240;
    exp_40_ram[1860] = 7;
    exp_40_ram[1861] = 135;
    exp_40_ram[1862] = 7;
    exp_40_ram[1863] = 135;
    exp_40_ram[1864] = 23;
    exp_40_ram[1865] = 69;
    exp_40_ram[1866] = 6;
    exp_40_ram[1867] = 198;
    exp_40_ram[1868] = 6;
    exp_40_ram[1869] = 198;
    exp_40_ram[1870] = 7;
    exp_40_ram[1871] = 71;
    exp_40_ram[1872] = 128;
    exp_40_ram[1873] = 128;
    exp_40_ram[1874] = 129;
    exp_40_ram[1875] = 129;
    exp_40_ram[1876] = 7;
    exp_40_ram[1877] = 23;
    exp_40_ram[1878] = 133;
    exp_40_ram[1879] = 5;
    exp_40_ram[1880] = 240;
    exp_40_ram[1881] = 7;
    exp_40_ram[1882] = 138;
    exp_40_ram[1883] = 23;
    exp_40_ram[1884] = 133;
    exp_40_ram[1885] = 224;
    exp_40_ram[1886] = 0;
    exp_40_ram[1887] = 7;
    exp_40_ram[1888] = 103;
    exp_40_ram[1889] = 7;
    exp_40_ram[1890] = 144;
    exp_40_ram[1891] = 129;
    exp_40_ram[1892] = 7;
    exp_40_ram[1893] = 23;
    exp_40_ram[1894] = 133;
    exp_40_ram[1895] = 5;
    exp_40_ram[1896] = 240;
    exp_40_ram[1897] = 7;
    exp_40_ram[1898] = 138;
    exp_40_ram[1899] = 23;
    exp_40_ram[1900] = 133;
    exp_40_ram[1901] = 224;
    exp_40_ram[1902] = 0;
    exp_40_ram[1903] = 2;
    exp_40_ram[1904] = 7;
    exp_40_ram[1905] = 199;
    exp_40_ram[1906] = 138;
    exp_40_ram[1907] = 23;
    exp_40_ram[1908] = 133;
    exp_40_ram[1909] = 224;
    exp_40_ram[1910] = 0;
    exp_40_ram[1911] = 23;
    exp_40_ram[1912] = 133;
    exp_40_ram[1913] = 224;
    exp_40_ram[1914] = 23;
    exp_40_ram[1915] = 133;
    exp_40_ram[1916] = 224;
    exp_40_ram[1917] = 7;
    exp_40_ram[1918] = 103;
    exp_40_ram[1919] = 7;
    exp_40_ram[1920] = 144;
    exp_40_ram[1921] = 129;
    exp_40_ram[1922] = 7;
    exp_40_ram[1923] = 6;
    exp_40_ram[1924] = 23;
    exp_40_ram[1925] = 133;
    exp_40_ram[1926] = 5;
    exp_40_ram[1927] = 224;
    exp_40_ram[1928] = 7;
    exp_40_ram[1929] = 23;
    exp_40_ram[1930] = 133;
    exp_40_ram[1931] = 5;
    exp_40_ram[1932] = 224;
    exp_40_ram[1933] = 7;
    exp_40_ram[1934] = 138;
    exp_40_ram[1935] = 23;
    exp_40_ram[1936] = 133;
    exp_40_ram[1937] = 224;
    exp_40_ram[1938] = 0;
    exp_40_ram[1939] = 2;
    exp_40_ram[1940] = 7;
    exp_40_ram[1941] = 6;
    exp_40_ram[1942] = 23;
    exp_40_ram[1943] = 133;
    exp_40_ram[1944] = 5;
    exp_40_ram[1945] = 224;
    exp_40_ram[1946] = 7;
    exp_40_ram[1947] = 23;
    exp_40_ram[1948] = 133;
    exp_40_ram[1949] = 5;
    exp_40_ram[1950] = 224;
    exp_40_ram[1951] = 7;
    exp_40_ram[1952] = 138;
    exp_40_ram[1953] = 23;
    exp_40_ram[1954] = 133;
    exp_40_ram[1955] = 224;
    exp_40_ram[1956] = 0;
    exp_40_ram[1957] = 7;
    exp_40_ram[1958] = 103;
    exp_40_ram[1959] = 7;
    exp_40_ram[1960] = 144;
    exp_40_ram[1961] = 129;
    exp_40_ram[1962] = 7;
    exp_40_ram[1963] = 23;
    exp_40_ram[1964] = 133;
    exp_40_ram[1965] = 5;
    exp_40_ram[1966] = 224;
    exp_40_ram[1967] = 7;
    exp_40_ram[1968] = 138;
    exp_40_ram[1969] = 23;
    exp_40_ram[1970] = 133;
    exp_40_ram[1971] = 224;
    exp_40_ram[1972] = 0;
    exp_40_ram[1973] = 2;
    exp_40_ram[1974] = 7;
    exp_40_ram[1975] = 199;
    exp_40_ram[1976] = 138;
    exp_40_ram[1977] = 23;
    exp_40_ram[1978] = 133;
    exp_40_ram[1979] = 224;
    exp_40_ram[1980] = 0;
    exp_40_ram[1981] = 23;
    exp_40_ram[1982] = 133;
    exp_40_ram[1983] = 224;
    exp_40_ram[1984] = 23;
    exp_40_ram[1985] = 133;
    exp_40_ram[1986] = 224;
    exp_40_ram[1987] = 23;
    exp_40_ram[1988] = 133;
    exp_40_ram[1989] = 224;
    exp_40_ram[1990] = 23;
    exp_40_ram[1991] = 133;
    exp_40_ram[1992] = 224;
    exp_40_ram[1993] = 23;
    exp_40_ram[1994] = 133;
    exp_40_ram[1995] = 224;
    exp_40_ram[1996] = 23;
    exp_40_ram[1997] = 133;
    exp_40_ram[1998] = 224;
    exp_40_ram[1999] = 23;
    exp_40_ram[2000] = 133;
    exp_40_ram[2001] = 224;
    exp_40_ram[2002] = 23;
    exp_40_ram[2003] = 133;
    exp_40_ram[2004] = 224;
    exp_40_ram[2005] = 7;
    exp_40_ram[2006] = 55;
    exp_40_ram[2007] = 7;
    exp_40_ram[2008] = 160;
    exp_40_ram[2009] = 130;
    exp_40_ram[2010] = 7;
    exp_40_ram[2011] = 6;
    exp_40_ram[2012] = 5;
    exp_40_ram[2013] = 133;
    exp_40_ram[2014] = 224;
    exp_40_ram[2015] = 7;
    exp_40_ram[2016] = 7;
    exp_40_ram[2017] = 10;
    exp_40_ram[2018] = 23;
    exp_40_ram[2019] = 133;
    exp_40_ram[2020] = 224;
    exp_40_ram[2021] = 0;
    exp_40_ram[2022] = 7;
    exp_40_ram[2023] = 6;
    exp_40_ram[2024] = 5;
    exp_40_ram[2025] = 133;
    exp_40_ram[2026] = 224;
    exp_40_ram[2027] = 7;
    exp_40_ram[2028] = 7;
    exp_40_ram[2029] = 7;
    exp_40_ram[2030] = 7;
    exp_40_ram[2031] = 10;
    exp_40_ram[2032] = 23;
    exp_40_ram[2033] = 133;
    exp_40_ram[2034] = 224;
    exp_40_ram[2035] = 0;
    exp_40_ram[2036] = 7;
    exp_40_ram[2037] = 6;
    exp_40_ram[2038] = 5;
    exp_40_ram[2039] = 133;
    exp_40_ram[2040] = 224;
    exp_40_ram[2041] = 7;
    exp_40_ram[2042] = 7;
    exp_40_ram[2043] = 7;
    exp_40_ram[2044] = 7;
    exp_40_ram[2045] = 10;
    exp_40_ram[2046] = 23;
    exp_40_ram[2047] = 133;
    exp_40_ram[2048] = 224;
    exp_40_ram[2049] = 0;
    exp_40_ram[2050] = 7;
    exp_40_ram[2051] = 6;
    exp_40_ram[2052] = 5;
    exp_40_ram[2053] = 133;
    exp_40_ram[2054] = 224;
    exp_40_ram[2055] = 7;
    exp_40_ram[2056] = 7;
    exp_40_ram[2057] = 7;
    exp_40_ram[2058] = 7;
    exp_40_ram[2059] = 10;
    exp_40_ram[2060] = 23;
    exp_40_ram[2061] = 133;
    exp_40_ram[2062] = 224;
    exp_40_ram[2063] = 0;
    exp_40_ram[2064] = 7;
    exp_40_ram[2065] = 6;
    exp_40_ram[2066] = 5;
    exp_40_ram[2067] = 133;
    exp_40_ram[2068] = 224;
    exp_40_ram[2069] = 7;
    exp_40_ram[2070] = 138;
    exp_40_ram[2071] = 23;
    exp_40_ram[2072] = 133;
    exp_40_ram[2073] = 224;
    exp_40_ram[2074] = 0;
    exp_40_ram[2075] = 23;
    exp_40_ram[2076] = 133;
    exp_40_ram[2077] = 224;
    exp_40_ram[2078] = 23;
    exp_40_ram[2079] = 133;
    exp_40_ram[2080] = 224;
    exp_40_ram[2081] = 7;
    exp_40_ram[2082] = 55;
    exp_40_ram[2083] = 7;
    exp_40_ram[2084] = 160;
    exp_40_ram[2085] = 55;
    exp_40_ram[2086] = 7;
    exp_40_ram[2087] = 162;
    exp_40_ram[2088] = 132;
    exp_40_ram[2089] = 7;
    exp_40_ram[2090] = 5;
    exp_40_ram[2091] = 133;
    exp_40_ram[2092] = 224;
    exp_40_ram[2093] = 7;
    exp_40_ram[2094] = 7;
    exp_40_ram[2095] = 10;
    exp_40_ram[2096] = 23;
    exp_40_ram[2097] = 133;
    exp_40_ram[2098] = 224;
    exp_40_ram[2099] = 0;
    exp_40_ram[2100] = 7;
    exp_40_ram[2101] = 5;
    exp_40_ram[2102] = 133;
    exp_40_ram[2103] = 224;
    exp_40_ram[2104] = 7;
    exp_40_ram[2105] = 7;
    exp_40_ram[2106] = 7;
    exp_40_ram[2107] = 7;
    exp_40_ram[2108] = 10;
    exp_40_ram[2109] = 23;
    exp_40_ram[2110] = 133;
    exp_40_ram[2111] = 224;
    exp_40_ram[2112] = 0;
    exp_40_ram[2113] = 7;
    exp_40_ram[2114] = 5;
    exp_40_ram[2115] = 133;
    exp_40_ram[2116] = 224;
    exp_40_ram[2117] = 7;
    exp_40_ram[2118] = 7;
    exp_40_ram[2119] = 7;
    exp_40_ram[2120] = 7;
    exp_40_ram[2121] = 10;
    exp_40_ram[2122] = 23;
    exp_40_ram[2123] = 133;
    exp_40_ram[2124] = 224;
    exp_40_ram[2125] = 0;
    exp_40_ram[2126] = 7;
    exp_40_ram[2127] = 5;
    exp_40_ram[2128] = 133;
    exp_40_ram[2129] = 224;
    exp_40_ram[2130] = 7;
    exp_40_ram[2131] = 7;
    exp_40_ram[2132] = 7;
    exp_40_ram[2133] = 7;
    exp_40_ram[2134] = 10;
    exp_40_ram[2135] = 23;
    exp_40_ram[2136] = 133;
    exp_40_ram[2137] = 224;
    exp_40_ram[2138] = 0;
    exp_40_ram[2139] = 7;
    exp_40_ram[2140] = 133;
    exp_40_ram[2141] = 224;
    exp_40_ram[2142] = 7;
    exp_40_ram[2143] = 135;
    exp_40_ram[2144] = 7;
    exp_40_ram[2145] = 135;
    exp_40_ram[2146] = 7;
    exp_40_ram[2147] = 7;
    exp_40_ram[2148] = 7;
    exp_40_ram[2149] = 10;
    exp_40_ram[2150] = 23;
    exp_40_ram[2151] = 133;
    exp_40_ram[2152] = 224;
    exp_40_ram[2153] = 0;
    exp_40_ram[2154] = 7;
    exp_40_ram[2155] = 5;
    exp_40_ram[2156] = 133;
    exp_40_ram[2157] = 224;
    exp_40_ram[2158] = 7;
    exp_40_ram[2159] = 138;
    exp_40_ram[2160] = 23;
    exp_40_ram[2161] = 133;
    exp_40_ram[2162] = 224;
    exp_40_ram[2163] = 0;
    exp_40_ram[2164] = 23;
    exp_40_ram[2165] = 133;
    exp_40_ram[2166] = 224;
    exp_40_ram[2167] = 23;
    exp_40_ram[2168] = 133;
    exp_40_ram[2169] = 224;
    exp_40_ram[2170] = 7;
    exp_40_ram[2171] = 55;
    exp_40_ram[2172] = 7;
    exp_40_ram[2173] = 160;
    exp_40_ram[2174] = 130;
    exp_40_ram[2175] = 7;
    exp_40_ram[2176] = 23;
    exp_40_ram[2177] = 133;
    exp_40_ram[2178] = 5;
    exp_40_ram[2179] = 224;
    exp_40_ram[2180] = 7;
    exp_40_ram[2181] = 138;
    exp_40_ram[2182] = 23;
    exp_40_ram[2183] = 133;
    exp_40_ram[2184] = 224;
    exp_40_ram[2185] = 0;
    exp_40_ram[2186] = 7;
    exp_40_ram[2187] = 23;
    exp_40_ram[2188] = 133;
    exp_40_ram[2189] = 5;
    exp_40_ram[2190] = 224;
    exp_40_ram[2191] = 7;
    exp_40_ram[2192] = 7;
    exp_40_ram[2193] = 10;
    exp_40_ram[2194] = 23;
    exp_40_ram[2195] = 133;
    exp_40_ram[2196] = 224;
    exp_40_ram[2197] = 0;
    exp_40_ram[2198] = 7;
    exp_40_ram[2199] = 23;
    exp_40_ram[2200] = 133;
    exp_40_ram[2201] = 5;
    exp_40_ram[2202] = 224;
    exp_40_ram[2203] = 7;
    exp_40_ram[2204] = 7;
    exp_40_ram[2205] = 10;
    exp_40_ram[2206] = 23;
    exp_40_ram[2207] = 133;
    exp_40_ram[2208] = 224;
    exp_40_ram[2209] = 0;
    exp_40_ram[2210] = 7;
    exp_40_ram[2211] = 23;
    exp_40_ram[2212] = 133;
    exp_40_ram[2213] = 5;
    exp_40_ram[2214] = 224;
    exp_40_ram[2215] = 7;
    exp_40_ram[2216] = 7;
    exp_40_ram[2217] = 10;
    exp_40_ram[2218] = 23;
    exp_40_ram[2219] = 133;
    exp_40_ram[2220] = 224;
    exp_40_ram[2221] = 0;
    exp_40_ram[2222] = 7;
    exp_40_ram[2223] = 23;
    exp_40_ram[2224] = 133;
    exp_40_ram[2225] = 5;
    exp_40_ram[2226] = 224;
    exp_40_ram[2227] = 7;
    exp_40_ram[2228] = 7;
    exp_40_ram[2229] = 10;
    exp_40_ram[2230] = 23;
    exp_40_ram[2231] = 133;
    exp_40_ram[2232] = 224;
    exp_40_ram[2233] = 0;
    exp_40_ram[2234] = 23;
    exp_40_ram[2235] = 133;
    exp_40_ram[2236] = 224;
    exp_40_ram[2237] = 23;
    exp_40_ram[2238] = 133;
    exp_40_ram[2239] = 224;
    exp_40_ram[2240] = 7;
    exp_40_ram[2241] = 55;
    exp_40_ram[2242] = 7;
    exp_40_ram[2243] = 160;
    exp_40_ram[2244] = 130;
    exp_40_ram[2245] = 7;
    exp_40_ram[2246] = 23;
    exp_40_ram[2247] = 133;
    exp_40_ram[2248] = 5;
    exp_40_ram[2249] = 224;
    exp_40_ram[2250] = 7;
    exp_40_ram[2251] = 7;
    exp_40_ram[2252] = 10;
    exp_40_ram[2253] = 23;
    exp_40_ram[2254] = 133;
    exp_40_ram[2255] = 224;
    exp_40_ram[2256] = 0;
    exp_40_ram[2257] = 7;
    exp_40_ram[2258] = 23;
    exp_40_ram[2259] = 133;
    exp_40_ram[2260] = 5;
    exp_40_ram[2261] = 224;
    exp_40_ram[2262] = 7;
    exp_40_ram[2263] = 7;
    exp_40_ram[2264] = 7;
    exp_40_ram[2265] = 7;
    exp_40_ram[2266] = 10;
    exp_40_ram[2267] = 23;
    exp_40_ram[2268] = 133;
    exp_40_ram[2269] = 224;
    exp_40_ram[2270] = 0;
    exp_40_ram[2271] = 7;
    exp_40_ram[2272] = 23;
    exp_40_ram[2273] = 133;
    exp_40_ram[2274] = 5;
    exp_40_ram[2275] = 224;
    exp_40_ram[2276] = 7;
    exp_40_ram[2277] = 7;
    exp_40_ram[2278] = 7;
    exp_40_ram[2279] = 7;
    exp_40_ram[2280] = 10;
    exp_40_ram[2281] = 23;
    exp_40_ram[2282] = 133;
    exp_40_ram[2283] = 224;
    exp_40_ram[2284] = 0;
    exp_40_ram[2285] = 7;
    exp_40_ram[2286] = 23;
    exp_40_ram[2287] = 133;
    exp_40_ram[2288] = 5;
    exp_40_ram[2289] = 224;
    exp_40_ram[2290] = 7;
    exp_40_ram[2291] = 7;
    exp_40_ram[2292] = 7;
    exp_40_ram[2293] = 7;
    exp_40_ram[2294] = 10;
    exp_40_ram[2295] = 23;
    exp_40_ram[2296] = 133;
    exp_40_ram[2297] = 224;
    exp_40_ram[2298] = 0;
    exp_40_ram[2299] = 7;
    exp_40_ram[2300] = 23;
    exp_40_ram[2301] = 133;
    exp_40_ram[2302] = 5;
    exp_40_ram[2303] = 224;
    exp_40_ram[2304] = 7;
    exp_40_ram[2305] = 138;
    exp_40_ram[2306] = 23;
    exp_40_ram[2307] = 133;
    exp_40_ram[2308] = 224;
    exp_40_ram[2309] = 0;
    exp_40_ram[2310] = 23;
    exp_40_ram[2311] = 133;
    exp_40_ram[2312] = 224;
    exp_40_ram[2313] = 23;
    exp_40_ram[2314] = 133;
    exp_40_ram[2315] = 224;
    exp_40_ram[2316] = 7;
    exp_40_ram[2317] = 55;
    exp_40_ram[2318] = 7;
    exp_40_ram[2319] = 160;
    exp_40_ram[2320] = 55;
    exp_40_ram[2321] = 7;
    exp_40_ram[2322] = 162;
    exp_40_ram[2323] = 132;
    exp_40_ram[2324] = 7;
    exp_40_ram[2325] = 5;
    exp_40_ram[2326] = 133;
    exp_40_ram[2327] = 224;
    exp_40_ram[2328] = 7;
    exp_40_ram[2329] = 7;
    exp_40_ram[2330] = 7;
    exp_40_ram[2331] = 7;
    exp_40_ram[2332] = 10;
    exp_40_ram[2333] = 23;
    exp_40_ram[2334] = 133;
    exp_40_ram[2335] = 224;
    exp_40_ram[2336] = 0;
    exp_40_ram[2337] = 7;
    exp_40_ram[2338] = 5;
    exp_40_ram[2339] = 133;
    exp_40_ram[2340] = 224;
    exp_40_ram[2341] = 7;
    exp_40_ram[2342] = 7;
    exp_40_ram[2343] = 7;
    exp_40_ram[2344] = 7;
    exp_40_ram[2345] = 10;
    exp_40_ram[2346] = 23;
    exp_40_ram[2347] = 133;
    exp_40_ram[2348] = 224;
    exp_40_ram[2349] = 0;
    exp_40_ram[2350] = 7;
    exp_40_ram[2351] = 5;
    exp_40_ram[2352] = 133;
    exp_40_ram[2353] = 224;
    exp_40_ram[2354] = 7;
    exp_40_ram[2355] = 7;
    exp_40_ram[2356] = 7;
    exp_40_ram[2357] = 7;
    exp_40_ram[2358] = 10;
    exp_40_ram[2359] = 23;
    exp_40_ram[2360] = 133;
    exp_40_ram[2361] = 224;
    exp_40_ram[2362] = 0;
    exp_40_ram[2363] = 7;
    exp_40_ram[2364] = 5;
    exp_40_ram[2365] = 133;
    exp_40_ram[2366] = 224;
    exp_40_ram[2367] = 7;
    exp_40_ram[2368] = 7;
    exp_40_ram[2369] = 7;
    exp_40_ram[2370] = 7;
    exp_40_ram[2371] = 10;
    exp_40_ram[2372] = 23;
    exp_40_ram[2373] = 133;
    exp_40_ram[2374] = 224;
    exp_40_ram[2375] = 0;
    exp_40_ram[2376] = 7;
    exp_40_ram[2377] = 133;
    exp_40_ram[2378] = 224;
    exp_40_ram[2379] = 7;
    exp_40_ram[2380] = 135;
    exp_40_ram[2381] = 7;
    exp_40_ram[2382] = 135;
    exp_40_ram[2383] = 7;
    exp_40_ram[2384] = 7;
    exp_40_ram[2385] = 7;
    exp_40_ram[2386] = 10;
    exp_40_ram[2387] = 23;
    exp_40_ram[2388] = 133;
    exp_40_ram[2389] = 224;
    exp_40_ram[2390] = 0;
    exp_40_ram[2391] = 7;
    exp_40_ram[2392] = 5;
    exp_40_ram[2393] = 133;
    exp_40_ram[2394] = 224;
    exp_40_ram[2395] = 7;
    exp_40_ram[2396] = 138;
    exp_40_ram[2397] = 23;
    exp_40_ram[2398] = 133;
    exp_40_ram[2399] = 224;
    exp_40_ram[2400] = 0;
    exp_40_ram[2401] = 23;
    exp_40_ram[2402] = 133;
    exp_40_ram[2403] = 224;
    exp_40_ram[2404] = 23;
    exp_40_ram[2405] = 133;
    exp_40_ram[2406] = 224;
    exp_40_ram[2407] = 7;
    exp_40_ram[2408] = 55;
    exp_40_ram[2409] = 7;
    exp_40_ram[2410] = 160;
    exp_40_ram[2411] = 130;
    exp_40_ram[2412] = 7;
    exp_40_ram[2413] = 23;
    exp_40_ram[2414] = 133;
    exp_40_ram[2415] = 5;
    exp_40_ram[2416] = 224;
    exp_40_ram[2417] = 7;
    exp_40_ram[2418] = 7;
    exp_40_ram[2419] = 10;
    exp_40_ram[2420] = 23;
    exp_40_ram[2421] = 133;
    exp_40_ram[2422] = 224;
    exp_40_ram[2423] = 0;
    exp_40_ram[2424] = 7;
    exp_40_ram[2425] = 23;
    exp_40_ram[2426] = 133;
    exp_40_ram[2427] = 5;
    exp_40_ram[2428] = 224;
    exp_40_ram[2429] = 7;
    exp_40_ram[2430] = 7;
    exp_40_ram[2431] = 10;
    exp_40_ram[2432] = 23;
    exp_40_ram[2433] = 133;
    exp_40_ram[2434] = 224;
    exp_40_ram[2435] = 0;
    exp_40_ram[2436] = 7;
    exp_40_ram[2437] = 23;
    exp_40_ram[2438] = 133;
    exp_40_ram[2439] = 5;
    exp_40_ram[2440] = 224;
    exp_40_ram[2441] = 7;
    exp_40_ram[2442] = 7;
    exp_40_ram[2443] = 10;
    exp_40_ram[2444] = 23;
    exp_40_ram[2445] = 133;
    exp_40_ram[2446] = 224;
    exp_40_ram[2447] = 0;
    exp_40_ram[2448] = 7;
    exp_40_ram[2449] = 23;
    exp_40_ram[2450] = 133;
    exp_40_ram[2451] = 5;
    exp_40_ram[2452] = 224;
    exp_40_ram[2453] = 7;
    exp_40_ram[2454] = 138;
    exp_40_ram[2455] = 23;
    exp_40_ram[2456] = 133;
    exp_40_ram[2457] = 224;
    exp_40_ram[2458] = 0;
    exp_40_ram[2459] = 7;
    exp_40_ram[2460] = 23;
    exp_40_ram[2461] = 133;
    exp_40_ram[2462] = 5;
    exp_40_ram[2463] = 224;
    exp_40_ram[2464] = 7;
    exp_40_ram[2465] = 7;
    exp_40_ram[2466] = 10;
    exp_40_ram[2467] = 23;
    exp_40_ram[2468] = 133;
    exp_40_ram[2469] = 224;
    exp_40_ram[2470] = 0;
    exp_40_ram[2471] = 23;
    exp_40_ram[2472] = 133;
    exp_40_ram[2473] = 224;
    exp_40_ram[2474] = 23;
    exp_40_ram[2475] = 133;
    exp_40_ram[2476] = 224;
    exp_40_ram[2477] = 7;
    exp_40_ram[2478] = 55;
    exp_40_ram[2479] = 7;
    exp_40_ram[2480] = 160;
    exp_40_ram[2481] = 130;
    exp_40_ram[2482] = 7;
    exp_40_ram[2483] = 23;
    exp_40_ram[2484] = 133;
    exp_40_ram[2485] = 5;
    exp_40_ram[2486] = 224;
    exp_40_ram[2487] = 7;
    exp_40_ram[2488] = 7;
    exp_40_ram[2489] = 10;
    exp_40_ram[2490] = 23;
    exp_40_ram[2491] = 133;
    exp_40_ram[2492] = 224;
    exp_40_ram[2493] = 0;
    exp_40_ram[2494] = 7;
    exp_40_ram[2495] = 23;
    exp_40_ram[2496] = 133;
    exp_40_ram[2497] = 5;
    exp_40_ram[2498] = 224;
    exp_40_ram[2499] = 7;
    exp_40_ram[2500] = 7;
    exp_40_ram[2501] = 7;
    exp_40_ram[2502] = 7;
    exp_40_ram[2503] = 10;
    exp_40_ram[2504] = 23;
    exp_40_ram[2505] = 133;
    exp_40_ram[2506] = 224;
    exp_40_ram[2507] = 0;
    exp_40_ram[2508] = 7;
    exp_40_ram[2509] = 23;
    exp_40_ram[2510] = 133;
    exp_40_ram[2511] = 5;
    exp_40_ram[2512] = 224;
    exp_40_ram[2513] = 7;
    exp_40_ram[2514] = 7;
    exp_40_ram[2515] = 7;
    exp_40_ram[2516] = 7;
    exp_40_ram[2517] = 10;
    exp_40_ram[2518] = 23;
    exp_40_ram[2519] = 133;
    exp_40_ram[2520] = 224;
    exp_40_ram[2521] = 0;
    exp_40_ram[2522] = 7;
    exp_40_ram[2523] = 5;
    exp_40_ram[2524] = 133;
    exp_40_ram[2525] = 224;
    exp_40_ram[2526] = 7;
    exp_40_ram[2527] = 7;
    exp_40_ram[2528] = 7;
    exp_40_ram[2529] = 7;
    exp_40_ram[2530] = 10;
    exp_40_ram[2531] = 23;
    exp_40_ram[2532] = 133;
    exp_40_ram[2533] = 224;
    exp_40_ram[2534] = 0;
    exp_40_ram[2535] = 7;
    exp_40_ram[2536] = 23;
    exp_40_ram[2537] = 133;
    exp_40_ram[2538] = 5;
    exp_40_ram[2539] = 224;
    exp_40_ram[2540] = 7;
    exp_40_ram[2541] = 138;
    exp_40_ram[2542] = 23;
    exp_40_ram[2543] = 133;
    exp_40_ram[2544] = 224;
    exp_40_ram[2545] = 0;
    exp_40_ram[2546] = 23;
    exp_40_ram[2547] = 133;
    exp_40_ram[2548] = 224;
    exp_40_ram[2549] = 23;
    exp_40_ram[2550] = 133;
    exp_40_ram[2551] = 224;
    exp_40_ram[2552] = 7;
    exp_40_ram[2553] = 2;
    exp_40_ram[2554] = 7;
    exp_40_ram[2555] = 23;
    exp_40_ram[2556] = 133;
    exp_40_ram[2557] = 5;
    exp_40_ram[2558] = 224;
    exp_40_ram[2559] = 7;
    exp_40_ram[2560] = 138;
    exp_40_ram[2561] = 23;
    exp_40_ram[2562] = 133;
    exp_40_ram[2563] = 224;
    exp_40_ram[2564] = 0;
    exp_40_ram[2565] = 7;
    exp_40_ram[2566] = 6;
    exp_40_ram[2567] = 5;
    exp_40_ram[2568] = 133;
    exp_40_ram[2569] = 224;
    exp_40_ram[2570] = 7;
    exp_40_ram[2571] = 23;
    exp_40_ram[2572] = 133;
    exp_40_ram[2573] = 5;
    exp_40_ram[2574] = 224;
    exp_40_ram[2575] = 7;
    exp_40_ram[2576] = 138;
    exp_40_ram[2577] = 23;
    exp_40_ram[2578] = 133;
    exp_40_ram[2579] = 224;
    exp_40_ram[2580] = 0;
    exp_40_ram[2581] = 7;
    exp_40_ram[2582] = 6;
    exp_40_ram[2583] = 5;
    exp_40_ram[2584] = 133;
    exp_40_ram[2585] = 224;
    exp_40_ram[2586] = 7;
    exp_40_ram[2587] = 23;
    exp_40_ram[2588] = 133;
    exp_40_ram[2589] = 5;
    exp_40_ram[2590] = 224;
    exp_40_ram[2591] = 7;
    exp_40_ram[2592] = 138;
    exp_40_ram[2593] = 23;
    exp_40_ram[2594] = 133;
    exp_40_ram[2595] = 224;
    exp_40_ram[2596] = 0;
    exp_40_ram[2597] = 7;
    exp_40_ram[2598] = 6;
    exp_40_ram[2599] = 5;
    exp_40_ram[2600] = 133;
    exp_40_ram[2601] = 224;
    exp_40_ram[2602] = 7;
    exp_40_ram[2603] = 23;
    exp_40_ram[2604] = 133;
    exp_40_ram[2605] = 5;
    exp_40_ram[2606] = 224;
    exp_40_ram[2607] = 7;
    exp_40_ram[2608] = 138;
    exp_40_ram[2609] = 23;
    exp_40_ram[2610] = 133;
    exp_40_ram[2611] = 224;
    exp_40_ram[2612] = 0;
    exp_40_ram[2613] = 23;
    exp_40_ram[2614] = 133;
    exp_40_ram[2615] = 224;
    exp_40_ram[2616] = 23;
    exp_40_ram[2617] = 133;
    exp_40_ram[2618] = 224;
    exp_40_ram[2619] = 23;
    exp_40_ram[2620] = 133;
    exp_40_ram[2621] = 224;
    exp_40_ram[2622] = 32;
    exp_40_ram[2623] = 36;
    exp_40_ram[2624] = 1;
    exp_40_ram[2625] = 128;
    exp_40_ram[2626] = 1;
    exp_40_ram[2627] = 46;
    exp_40_ram[2628] = 44;
    exp_40_ram[2629] = 42;
    exp_40_ram[2630] = 40;
    exp_40_ram[2631] = 38;
    exp_40_ram[2632] = 36;
    exp_40_ram[2633] = 34;
    exp_40_ram[2634] = 32;
    exp_40_ram[2635] = 4;
    exp_40_ram[2636] = 23;
    exp_40_ram[2637] = 133;
    exp_40_ram[2638] = 224;
    exp_40_ram[2639] = 7;
    exp_40_ram[2640] = 32;
    exp_40_ram[2641] = 7;
    exp_40_ram[2642] = 46;
    exp_40_ram[2643] = 7;
    exp_40_ram[2644] = 44;
    exp_40_ram[2645] = 7;
    exp_40_ram[2646] = 42;
    exp_40_ram[2647] = 7;
    exp_40_ram[2648] = 40;
    exp_40_ram[2649] = 38;
    exp_40_ram[2650] = 7;
    exp_40_ram[2651] = 38;
    exp_40_ram[2652] = 7;
    exp_40_ram[2653] = 133;
    exp_40_ram[2654] = 240;
    exp_40_ram[2655] = 7;
    exp_40_ram[2656] = 135;
    exp_40_ram[2657] = 32;
    exp_40_ram[2658] = 34;
    exp_40_ram[2659] = 7;
    exp_40_ram[2660] = 133;
    exp_40_ram[2661] = 224;
    exp_40_ram[2662] = 7;
    exp_40_ram[2663] = 23;
    exp_40_ram[2664] = 133;
    exp_40_ram[2665] = 5;
    exp_40_ram[2666] = 224;
    exp_40_ram[2667] = 7;
    exp_40_ram[2668] = 138;
    exp_40_ram[2669] = 23;
    exp_40_ram[2670] = 133;
    exp_40_ram[2671] = 224;
    exp_40_ram[2672] = 0;
    exp_40_ram[2673] = 7;
    exp_40_ram[2674] = 133;
    exp_40_ram[2675] = 240;
    exp_40_ram[2676] = 7;
    exp_40_ram[2677] = 133;
    exp_40_ram[2678] = 224;
    exp_40_ram[2679] = 7;
    exp_40_ram[2680] = 23;
    exp_40_ram[2681] = 133;
    exp_40_ram[2682] = 5;
    exp_40_ram[2683] = 224;
    exp_40_ram[2684] = 7;
    exp_40_ram[2685] = 138;
    exp_40_ram[2686] = 23;
    exp_40_ram[2687] = 133;
    exp_40_ram[2688] = 224;
    exp_40_ram[2689] = 0;
    exp_40_ram[2690] = 7;
    exp_40_ram[2691] = 133;
    exp_40_ram[2692] = 240;
    exp_40_ram[2693] = 7;
    exp_40_ram[2694] = 133;
    exp_40_ram[2695] = 224;
    exp_40_ram[2696] = 7;
    exp_40_ram[2697] = 23;
    exp_40_ram[2698] = 133;
    exp_40_ram[2699] = 5;
    exp_40_ram[2700] = 224;
    exp_40_ram[2701] = 7;
    exp_40_ram[2702] = 138;
    exp_40_ram[2703] = 23;
    exp_40_ram[2704] = 133;
    exp_40_ram[2705] = 224;
    exp_40_ram[2706] = 0;
    exp_40_ram[2707] = 7;
    exp_40_ram[2708] = 133;
    exp_40_ram[2709] = 240;
    exp_40_ram[2710] = 7;
    exp_40_ram[2711] = 23;
    exp_40_ram[2712] = 133;
    exp_40_ram[2713] = 5;
    exp_40_ram[2714] = 224;
    exp_40_ram[2715] = 7;
    exp_40_ram[2716] = 138;
    exp_40_ram[2717] = 23;
    exp_40_ram[2718] = 133;
    exp_40_ram[2719] = 224;
    exp_40_ram[2720] = 0;
    exp_40_ram[2721] = 7;
    exp_40_ram[2722] = 32;
    exp_40_ram[2723] = 7;
    exp_40_ram[2724] = 46;
    exp_40_ram[2725] = 7;
    exp_40_ram[2726] = 44;
    exp_40_ram[2727] = 7;
    exp_40_ram[2728] = 42;
    exp_40_ram[2729] = 7;
    exp_40_ram[2730] = 40;
    exp_40_ram[2731] = 38;
    exp_40_ram[2732] = 7;
    exp_40_ram[2733] = 38;
    exp_40_ram[2734] = 7;
    exp_40_ram[2735] = 133;
    exp_40_ram[2736] = 224;
    exp_40_ram[2737] = 7;
    exp_40_ram[2738] = 135;
    exp_40_ram[2739] = 32;
    exp_40_ram[2740] = 34;
    exp_40_ram[2741] = 7;
    exp_40_ram[2742] = 133;
    exp_40_ram[2743] = 224;
    exp_40_ram[2744] = 7;
    exp_40_ram[2745] = 23;
    exp_40_ram[2746] = 133;
    exp_40_ram[2747] = 5;
    exp_40_ram[2748] = 224;
    exp_40_ram[2749] = 7;
    exp_40_ram[2750] = 138;
    exp_40_ram[2751] = 23;
    exp_40_ram[2752] = 133;
    exp_40_ram[2753] = 224;
    exp_40_ram[2754] = 0;
    exp_40_ram[2755] = 7;
    exp_40_ram[2756] = 133;
    exp_40_ram[2757] = 240;
    exp_40_ram[2758] = 7;
    exp_40_ram[2759] = 133;
    exp_40_ram[2760] = 224;
    exp_40_ram[2761] = 7;
    exp_40_ram[2762] = 23;
    exp_40_ram[2763] = 133;
    exp_40_ram[2764] = 5;
    exp_40_ram[2765] = 224;
    exp_40_ram[2766] = 7;
    exp_40_ram[2767] = 138;
    exp_40_ram[2768] = 23;
    exp_40_ram[2769] = 133;
    exp_40_ram[2770] = 224;
    exp_40_ram[2771] = 0;
    exp_40_ram[2772] = 7;
    exp_40_ram[2773] = 133;
    exp_40_ram[2774] = 240;
    exp_40_ram[2775] = 7;
    exp_40_ram[2776] = 133;
    exp_40_ram[2777] = 224;
    exp_40_ram[2778] = 7;
    exp_40_ram[2779] = 23;
    exp_40_ram[2780] = 133;
    exp_40_ram[2781] = 5;
    exp_40_ram[2782] = 224;
    exp_40_ram[2783] = 7;
    exp_40_ram[2784] = 138;
    exp_40_ram[2785] = 23;
    exp_40_ram[2786] = 133;
    exp_40_ram[2787] = 224;
    exp_40_ram[2788] = 0;
    exp_40_ram[2789] = 7;
    exp_40_ram[2790] = 133;
    exp_40_ram[2791] = 240;
    exp_40_ram[2792] = 7;
    exp_40_ram[2793] = 23;
    exp_40_ram[2794] = 133;
    exp_40_ram[2795] = 5;
    exp_40_ram[2796] = 224;
    exp_40_ram[2797] = 7;
    exp_40_ram[2798] = 138;
    exp_40_ram[2799] = 23;
    exp_40_ram[2800] = 133;
    exp_40_ram[2801] = 224;
    exp_40_ram[2802] = 0;
    exp_40_ram[2803] = 7;
    exp_40_ram[2804] = 32;
    exp_40_ram[2805] = 7;
    exp_40_ram[2806] = 46;
    exp_40_ram[2807] = 7;
    exp_40_ram[2808] = 44;
    exp_40_ram[2809] = 7;
    exp_40_ram[2810] = 42;
    exp_40_ram[2811] = 7;
    exp_40_ram[2812] = 40;
    exp_40_ram[2813] = 38;
    exp_40_ram[2814] = 38;
    exp_40_ram[2815] = 7;
    exp_40_ram[2816] = 133;
    exp_40_ram[2817] = 224;
    exp_40_ram[2818] = 7;
    exp_40_ram[2819] = 135;
    exp_40_ram[2820] = 32;
    exp_40_ram[2821] = 34;
    exp_40_ram[2822] = 7;
    exp_40_ram[2823] = 133;
    exp_40_ram[2824] = 224;
    exp_40_ram[2825] = 7;
    exp_40_ram[2826] = 23;
    exp_40_ram[2827] = 133;
    exp_40_ram[2828] = 5;
    exp_40_ram[2829] = 224;
    exp_40_ram[2830] = 7;
    exp_40_ram[2831] = 138;
    exp_40_ram[2832] = 23;
    exp_40_ram[2833] = 133;
    exp_40_ram[2834] = 224;
    exp_40_ram[2835] = 0;
    exp_40_ram[2836] = 7;
    exp_40_ram[2837] = 133;
    exp_40_ram[2838] = 224;
    exp_40_ram[2839] = 7;
    exp_40_ram[2840] = 133;
    exp_40_ram[2841] = 224;
    exp_40_ram[2842] = 7;
    exp_40_ram[2843] = 23;
    exp_40_ram[2844] = 133;
    exp_40_ram[2845] = 5;
    exp_40_ram[2846] = 224;
    exp_40_ram[2847] = 7;
    exp_40_ram[2848] = 138;
    exp_40_ram[2849] = 23;
    exp_40_ram[2850] = 133;
    exp_40_ram[2851] = 224;
    exp_40_ram[2852] = 0;
    exp_40_ram[2853] = 7;
    exp_40_ram[2854] = 133;
    exp_40_ram[2855] = 224;
    exp_40_ram[2856] = 7;
    exp_40_ram[2857] = 133;
    exp_40_ram[2858] = 224;
    exp_40_ram[2859] = 7;
    exp_40_ram[2860] = 23;
    exp_40_ram[2861] = 133;
    exp_40_ram[2862] = 5;
    exp_40_ram[2863] = 224;
    exp_40_ram[2864] = 7;
    exp_40_ram[2865] = 138;
    exp_40_ram[2866] = 23;
    exp_40_ram[2867] = 133;
    exp_40_ram[2868] = 224;
    exp_40_ram[2869] = 0;
    exp_40_ram[2870] = 7;
    exp_40_ram[2871] = 133;
    exp_40_ram[2872] = 224;
    exp_40_ram[2873] = 7;
    exp_40_ram[2874] = 23;
    exp_40_ram[2875] = 133;
    exp_40_ram[2876] = 5;
    exp_40_ram[2877] = 224;
    exp_40_ram[2878] = 7;
    exp_40_ram[2879] = 138;
    exp_40_ram[2880] = 23;
    exp_40_ram[2881] = 133;
    exp_40_ram[2882] = 208;
    exp_40_ram[2883] = 0;
    exp_40_ram[2884] = 23;
    exp_40_ram[2885] = 133;
    exp_40_ram[2886] = 208;
    exp_40_ram[2887] = 7;
    exp_40_ram[2888] = 32;
    exp_40_ram[2889] = 7;
    exp_40_ram[2890] = 46;
    exp_40_ram[2891] = 7;
    exp_40_ram[2892] = 44;
    exp_40_ram[2893] = 42;
    exp_40_ram[2894] = 7;
    exp_40_ram[2895] = 40;
    exp_40_ram[2896] = 7;
    exp_40_ram[2897] = 38;
    exp_40_ram[2898] = 7;
    exp_40_ram[2899] = 38;
    exp_40_ram[2900] = 7;
    exp_40_ram[2901] = 133;
    exp_40_ram[2902] = 224;
    exp_40_ram[2903] = 7;
    exp_40_ram[2904] = 135;
    exp_40_ram[2905] = 32;
    exp_40_ram[2906] = 34;
    exp_40_ram[2907] = 39;
    exp_40_ram[2908] = 39;
    exp_40_ram[2909] = 5;
    exp_40_ram[2910] = 133;
    exp_40_ram[2911] = 224;
    exp_40_ram[2912] = 224;
    exp_40_ram[2913] = 44;
    exp_40_ram[2914] = 46;
    exp_40_ram[2915] = 42;
    exp_40_ram[2916] = 0;
    exp_40_ram[2917] = 0;
    exp_40_ram[2918] = 224;
    exp_40_ram[2919] = 7;
    exp_40_ram[2920] = 135;
    exp_40_ram[2921] = 38;
    exp_40_ram[2922] = 38;
    exp_40_ram[2923] = 5;
    exp_40_ram[2924] = 133;
    exp_40_ram[2925] = 224;
    exp_40_ram[2926] = 11;
    exp_40_ram[2927] = 139;
    exp_40_ram[2928] = 55;
    exp_40_ram[2929] = 167;
    exp_40_ram[2930] = 133;
    exp_40_ram[2931] = 208;
    exp_40_ram[2932] = 7;
    exp_40_ram[2933] = 135;
    exp_40_ram[2934] = 6;
    exp_40_ram[2935] = 134;
    exp_40_ram[2936] = 5;
    exp_40_ram[2937] = 133;
    exp_40_ram[2938] = 208;
    exp_40_ram[2939] = 7;
    exp_40_ram[2940] = 196;
    exp_40_ram[2941] = 55;
    exp_40_ram[2942] = 167;
    exp_40_ram[2943] = 138;
    exp_40_ram[2944] = 10;
    exp_40_ram[2945] = 38;
    exp_40_ram[2946] = 38;
    exp_40_ram[2947] = 7;
    exp_40_ram[2948] = 5;
    exp_40_ram[2949] = 181;
    exp_40_ram[2950] = 135;
    exp_40_ram[2951] = 134;
    exp_40_ram[2952] = 135;
    exp_40_ram[2953] = 44;
    exp_40_ram[2954] = 46;
    exp_40_ram[2955] = 5;
    exp_40_ram[2956] = 224;
    exp_40_ram[2957] = 7;
    exp_40_ram[2958] = 135;
    exp_40_ram[2959] = 32;
    exp_40_ram[2960] = 34;
    exp_40_ram[2961] = 7;
    exp_40_ram[2962] = 133;
    exp_40_ram[2963] = 224;
    exp_40_ram[2964] = 7;
    exp_40_ram[2965] = 133;
    exp_40_ram[2966] = 208;
    exp_40_ram[2967] = 39;
    exp_40_ram[2968] = 135;
    exp_40_ram[2969] = 42;
    exp_40_ram[2970] = 39;
    exp_40_ram[2971] = 7;
    exp_40_ram[2972] = 210;
    exp_40_ram[2973] = 7;
    exp_40_ram[2974] = 32;
    exp_40_ram[2975] = 7;
    exp_40_ram[2976] = 46;
    exp_40_ram[2977] = 7;
    exp_40_ram[2978] = 44;
    exp_40_ram[2979] = 7;
    exp_40_ram[2980] = 42;
    exp_40_ram[2981] = 7;
    exp_40_ram[2982] = 40;
    exp_40_ram[2983] = 7;
    exp_40_ram[2984] = 38;
    exp_40_ram[2985] = 7;
    exp_40_ram[2986] = 38;
    exp_40_ram[2987] = 7;
    exp_40_ram[2988] = 133;
    exp_40_ram[2989] = 224;
    exp_40_ram[2990] = 7;
    exp_40_ram[2991] = 135;
    exp_40_ram[2992] = 32;
    exp_40_ram[2993] = 34;
    exp_40_ram[2994] = 7;
    exp_40_ram[2995] = 133;
    exp_40_ram[2996] = 224;
    exp_40_ram[2997] = 7;
    exp_40_ram[2998] = 133;
    exp_40_ram[2999] = 208;
    exp_40_ram[3000] = 7;
    exp_40_ram[3001] = 133;
    exp_40_ram[3002] = 224;
    exp_40_ram[3003] = 7;
    exp_40_ram[3004] = 133;
    exp_40_ram[3005] = 208;
    exp_40_ram[3006] = 39;
    exp_40_ram[3007] = 39;
    exp_40_ram[3008] = 5;
    exp_40_ram[3009] = 133;
    exp_40_ram[3010] = 224;
    exp_40_ram[3011] = 5;
    exp_40_ram[3012] = 224;
    exp_40_ram[3013] = 7;
    exp_40_ram[3014] = 135;
    exp_40_ram[3015] = 32;
    exp_40_ram[3016] = 34;
    exp_40_ram[3017] = 7;
    exp_40_ram[3018] = 133;
    exp_40_ram[3019] = 224;
    exp_40_ram[3020] = 7;
    exp_40_ram[3021] = 133;
    exp_40_ram[3022] = 208;
    exp_40_ram[3023] = 224;
    exp_40_ram[3024] = 44;
    exp_40_ram[3025] = 46;
    exp_40_ram[3026] = 40;
    exp_40_ram[3027] = 0;
    exp_40_ram[3028] = 0;
    exp_40_ram[3029] = 224;
    exp_40_ram[3030] = 7;
    exp_40_ram[3031] = 135;
    exp_40_ram[3032] = 38;
    exp_40_ram[3033] = 38;
    exp_40_ram[3034] = 5;
    exp_40_ram[3035] = 133;
    exp_40_ram[3036] = 224;
    exp_40_ram[3037] = 10;
    exp_40_ram[3038] = 138;
    exp_40_ram[3039] = 55;
    exp_40_ram[3040] = 167;
    exp_40_ram[3041] = 133;
    exp_40_ram[3042] = 208;
    exp_40_ram[3043] = 7;
    exp_40_ram[3044] = 135;
    exp_40_ram[3045] = 6;
    exp_40_ram[3046] = 134;
    exp_40_ram[3047] = 5;
    exp_40_ram[3048] = 133;
    exp_40_ram[3049] = 208;
    exp_40_ram[3050] = 7;
    exp_40_ram[3051] = 196;
    exp_40_ram[3052] = 55;
    exp_40_ram[3053] = 167;
    exp_40_ram[3054] = 137;
    exp_40_ram[3055] = 9;
    exp_40_ram[3056] = 38;
    exp_40_ram[3057] = 38;
    exp_40_ram[3058] = 7;
    exp_40_ram[3059] = 5;
    exp_40_ram[3060] = 181;
    exp_40_ram[3061] = 135;
    exp_40_ram[3062] = 134;
    exp_40_ram[3063] = 135;
    exp_40_ram[3064] = 44;
    exp_40_ram[3065] = 46;
    exp_40_ram[3066] = 5;
    exp_40_ram[3067] = 224;
    exp_40_ram[3068] = 7;
    exp_40_ram[3069] = 135;
    exp_40_ram[3070] = 32;
    exp_40_ram[3071] = 34;
    exp_40_ram[3072] = 7;
    exp_40_ram[3073] = 133;
    exp_40_ram[3074] = 224;
    exp_40_ram[3075] = 7;
    exp_40_ram[3076] = 133;
    exp_40_ram[3077] = 208;
    exp_40_ram[3078] = 39;
    exp_40_ram[3079] = 135;
    exp_40_ram[3080] = 40;
    exp_40_ram[3081] = 39;
    exp_40_ram[3082] = 7;
    exp_40_ram[3083] = 210;
    exp_40_ram[3084] = 32;
    exp_40_ram[3085] = 36;
    exp_40_ram[3086] = 41;
    exp_40_ram[3087] = 41;
    exp_40_ram[3088] = 42;
    exp_40_ram[3089] = 42;
    exp_40_ram[3090] = 43;
    exp_40_ram[3091] = 43;
    exp_40_ram[3092] = 1;
    exp_40_ram[3093] = 128;
    exp_40_ram[3094] = 1;
    exp_40_ram[3095] = 38;
    exp_40_ram[3096] = 36;
    exp_40_ram[3097] = 4;
    exp_40_ram[3098] = 224;
    exp_40_ram[3099] = 240;
    exp_40_ram[3100] = 0;
    exp_40_ram[3101] = 32;
    exp_40_ram[3102] = 36;
    exp_40_ram[3103] = 1;
    exp_40_ram[3104] = 128;
    exp_40_ram[3105] = 7;
    exp_40_ram[3106] = 135;
    exp_40_ram[3107] = 69;
    exp_40_ram[3108] = 1;
    exp_40_ram[3109] = 101;
    exp_40_ram[3110] = 76;
    exp_40_ram[3111] = 214;
    exp_40_ram[3112] = 5;
    exp_40_ram[3113] = 133;
    exp_40_ram[3114] = 1;
    exp_40_ram[3115] = 128;
    exp_40_ram[3116] = 92;
    exp_40_ram[3117] = 5;
    exp_40_ram[3118] = 133;
    exp_40_ram[3119] = 240;
    exp_40_ram[3120] = 240;
    exp_40_ram[3121] = 0;
    exp_40_ram[3122] = 117;
    exp_40_ram[3123] = 110;
    exp_40_ram[3124] = 87;
    exp_40_ram[3125] = 104;
    exp_40_ram[3126] = 105;
    exp_40_ram[3127] = 0;
    exp_40_ram[3128] = 97;
    exp_40_ram[3129] = 98;
    exp_40_ram[3130] = 65;
    exp_40_ram[3131] = 97;
    exp_40_ram[3132] = 110;
    exp_40_ram[3133] = 65;
    exp_40_ram[3134] = 101;
    exp_40_ram[3135] = 116;
    exp_40_ram[3136] = 68;
    exp_40_ram[3137] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 55;
    exp_33_ram[32] = 19;
    exp_33_ram[33] = 239;
    exp_33_ram[34] = 111;
    exp_33_ram[35] = 147;
    exp_33_ram[36] = 147;
    exp_33_ram[37] = 19;
    exp_33_ram[38] = 19;
    exp_33_ram[39] = 19;
    exp_33_ram[40] = 99;
    exp_33_ram[41] = 183;
    exp_33_ram[42] = 147;
    exp_33_ram[43] = 99;
    exp_33_ram[44] = 55;
    exp_33_ram[45] = 99;
    exp_33_ram[46] = 19;
    exp_33_ram[47] = 51;
    exp_33_ram[48] = 19;
    exp_33_ram[49] = 51;
    exp_33_ram[50] = 179;
    exp_33_ram[51] = 131;
    exp_33_ram[52] = 19;
    exp_33_ram[53] = 51;
    exp_33_ram[54] = 179;
    exp_33_ram[55] = 99;
    exp_33_ram[56] = 179;
    exp_33_ram[57] = 51;
    exp_33_ram[58] = 51;
    exp_33_ram[59] = 179;
    exp_33_ram[60] = 51;
    exp_33_ram[61] = 147;
    exp_33_ram[62] = 179;
    exp_33_ram[63] = 19;
    exp_33_ram[64] = 19;
    exp_33_ram[65] = 147;
    exp_33_ram[66] = 51;
    exp_33_ram[67] = 19;
    exp_33_ram[68] = 179;
    exp_33_ram[69] = 19;
    exp_33_ram[70] = 179;
    exp_33_ram[71] = 99;
    exp_33_ram[72] = 179;
    exp_33_ram[73] = 19;
    exp_33_ram[74] = 99;
    exp_33_ram[75] = 99;
    exp_33_ram[76] = 19;
    exp_33_ram[77] = 179;
    exp_33_ram[78] = 179;
    exp_33_ram[79] = 51;
    exp_33_ram[80] = 19;
    exp_33_ram[81] = 19;
    exp_33_ram[82] = 179;
    exp_33_ram[83] = 19;
    exp_33_ram[84] = 51;
    exp_33_ram[85] = 179;
    exp_33_ram[86] = 19;
    exp_33_ram[87] = 99;
    exp_33_ram[88] = 51;
    exp_33_ram[89] = 19;
    exp_33_ram[90] = 99;
    exp_33_ram[91] = 99;
    exp_33_ram[92] = 19;
    exp_33_ram[93] = 19;
    exp_33_ram[94] = 51;
    exp_33_ram[95] = 147;
    exp_33_ram[96] = 111;
    exp_33_ram[97] = 55;
    exp_33_ram[98] = 19;
    exp_33_ram[99] = 227;
    exp_33_ram[100] = 19;
    exp_33_ram[101] = 111;
    exp_33_ram[102] = 99;
    exp_33_ram[103] = 19;
    exp_33_ram[104] = 51;
    exp_33_ram[105] = 55;
    exp_33_ram[106] = 99;
    exp_33_ram[107] = 19;
    exp_33_ram[108] = 99;
    exp_33_ram[109] = 19;
    exp_33_ram[110] = 51;
    exp_33_ram[111] = 179;
    exp_33_ram[112] = 3;
    exp_33_ram[113] = 19;
    exp_33_ram[114] = 51;
    exp_33_ram[115] = 179;
    exp_33_ram[116] = 99;
    exp_33_ram[117] = 179;
    exp_33_ram[118] = 147;
    exp_33_ram[119] = 147;
    exp_33_ram[120] = 19;
    exp_33_ram[121] = 19;
    exp_33_ram[122] = 19;
    exp_33_ram[123] = 179;
    exp_33_ram[124] = 179;
    exp_33_ram[125] = 147;
    exp_33_ram[126] = 51;
    exp_33_ram[127] = 51;
    exp_33_ram[128] = 19;
    exp_33_ram[129] = 99;
    exp_33_ram[130] = 51;
    exp_33_ram[131] = 19;
    exp_33_ram[132] = 99;
    exp_33_ram[133] = 99;
    exp_33_ram[134] = 19;
    exp_33_ram[135] = 51;
    exp_33_ram[136] = 51;
    exp_33_ram[137] = 179;
    exp_33_ram[138] = 19;
    exp_33_ram[139] = 19;
    exp_33_ram[140] = 51;
    exp_33_ram[141] = 147;
    exp_33_ram[142] = 51;
    exp_33_ram[143] = 179;
    exp_33_ram[144] = 19;
    exp_33_ram[145] = 99;
    exp_33_ram[146] = 51;
    exp_33_ram[147] = 19;
    exp_33_ram[148] = 99;
    exp_33_ram[149] = 99;
    exp_33_ram[150] = 19;
    exp_33_ram[151] = 19;
    exp_33_ram[152] = 51;
    exp_33_ram[153] = 103;
    exp_33_ram[154] = 55;
    exp_33_ram[155] = 19;
    exp_33_ram[156] = 227;
    exp_33_ram[157] = 19;
    exp_33_ram[158] = 111;
    exp_33_ram[159] = 51;
    exp_33_ram[160] = 51;
    exp_33_ram[161] = 51;
    exp_33_ram[162] = 179;
    exp_33_ram[163] = 51;
    exp_33_ram[164] = 147;
    exp_33_ram[165] = 51;
    exp_33_ram[166] = 51;
    exp_33_ram[167] = 147;
    exp_33_ram[168] = 147;
    exp_33_ram[169] = 147;
    exp_33_ram[170] = 51;
    exp_33_ram[171] = 19;
    exp_33_ram[172] = 51;
    exp_33_ram[173] = 179;
    exp_33_ram[174] = 147;
    exp_33_ram[175] = 99;
    exp_33_ram[176] = 51;
    exp_33_ram[177] = 147;
    exp_33_ram[178] = 99;
    exp_33_ram[179] = 99;
    exp_33_ram[180] = 147;
    exp_33_ram[181] = 51;
    exp_33_ram[182] = 179;
    exp_33_ram[183] = 51;
    exp_33_ram[184] = 19;
    exp_33_ram[185] = 19;
    exp_33_ram[186] = 179;
    exp_33_ram[187] = 19;
    exp_33_ram[188] = 51;
    exp_33_ram[189] = 179;
    exp_33_ram[190] = 19;
    exp_33_ram[191] = 99;
    exp_33_ram[192] = 179;
    exp_33_ram[193] = 19;
    exp_33_ram[194] = 99;
    exp_33_ram[195] = 99;
    exp_33_ram[196] = 19;
    exp_33_ram[197] = 179;
    exp_33_ram[198] = 147;
    exp_33_ram[199] = 179;
    exp_33_ram[200] = 179;
    exp_33_ram[201] = 111;
    exp_33_ram[202] = 99;
    exp_33_ram[203] = 55;
    exp_33_ram[204] = 99;
    exp_33_ram[205] = 19;
    exp_33_ram[206] = 179;
    exp_33_ram[207] = 147;
    exp_33_ram[208] = 55;
    exp_33_ram[209] = 51;
    exp_33_ram[210] = 19;
    exp_33_ram[211] = 51;
    exp_33_ram[212] = 3;
    exp_33_ram[213] = 19;
    exp_33_ram[214] = 51;
    exp_33_ram[215] = 179;
    exp_33_ram[216] = 99;
    exp_33_ram[217] = 19;
    exp_33_ram[218] = 227;
    exp_33_ram[219] = 51;
    exp_33_ram[220] = 19;
    exp_33_ram[221] = 111;
    exp_33_ram[222] = 55;
    exp_33_ram[223] = 147;
    exp_33_ram[224] = 227;
    exp_33_ram[225] = 147;
    exp_33_ram[226] = 111;
    exp_33_ram[227] = 51;
    exp_33_ram[228] = 179;
    exp_33_ram[229] = 51;
    exp_33_ram[230] = 51;
    exp_33_ram[231] = 147;
    exp_33_ram[232] = 179;
    exp_33_ram[233] = 179;
    exp_33_ram[234] = 51;
    exp_33_ram[235] = 51;
    exp_33_ram[236] = 51;
    exp_33_ram[237] = 147;
    exp_33_ram[238] = 147;
    exp_33_ram[239] = 19;
    exp_33_ram[240] = 51;
    exp_33_ram[241] = 147;
    exp_33_ram[242] = 51;
    exp_33_ram[243] = 51;
    exp_33_ram[244] = 19;
    exp_33_ram[245] = 99;
    exp_33_ram[246] = 51;
    exp_33_ram[247] = 19;
    exp_33_ram[248] = 99;
    exp_33_ram[249] = 99;
    exp_33_ram[250] = 19;
    exp_33_ram[251] = 51;
    exp_33_ram[252] = 51;
    exp_33_ram[253] = 179;
    exp_33_ram[254] = 51;
    exp_33_ram[255] = 147;
    exp_33_ram[256] = 51;
    exp_33_ram[257] = 147;
    exp_33_ram[258] = 147;
    exp_33_ram[259] = 179;
    exp_33_ram[260] = 19;
    exp_33_ram[261] = 99;
    exp_33_ram[262] = 179;
    exp_33_ram[263] = 19;
    exp_33_ram[264] = 99;
    exp_33_ram[265] = 99;
    exp_33_ram[266] = 19;
    exp_33_ram[267] = 179;
    exp_33_ram[268] = 19;
    exp_33_ram[269] = 183;
    exp_33_ram[270] = 51;
    exp_33_ram[271] = 147;
    exp_33_ram[272] = 51;
    exp_33_ram[273] = 19;
    exp_33_ram[274] = 179;
    exp_33_ram[275] = 19;
    exp_33_ram[276] = 179;
    exp_33_ram[277] = 51;
    exp_33_ram[278] = 179;
    exp_33_ram[279] = 19;
    exp_33_ram[280] = 51;
    exp_33_ram[281] = 51;
    exp_33_ram[282] = 51;
    exp_33_ram[283] = 51;
    exp_33_ram[284] = 99;
    exp_33_ram[285] = 51;
    exp_33_ram[286] = 147;
    exp_33_ram[287] = 51;
    exp_33_ram[288] = 99;
    exp_33_ram[289] = 227;
    exp_33_ram[290] = 183;
    exp_33_ram[291] = 147;
    exp_33_ram[292] = 51;
    exp_33_ram[293] = 19;
    exp_33_ram[294] = 51;
    exp_33_ram[295] = 179;
    exp_33_ram[296] = 51;
    exp_33_ram[297] = 147;
    exp_33_ram[298] = 227;
    exp_33_ram[299] = 19;
    exp_33_ram[300] = 111;
    exp_33_ram[301] = 147;
    exp_33_ram[302] = 19;
    exp_33_ram[303] = 111;
    exp_33_ram[304] = 55;
    exp_33_ram[305] = 19;
    exp_33_ram[306] = 19;
    exp_33_ram[307] = 179;
    exp_33_ram[308] = 147;
    exp_33_ram[309] = 19;
    exp_33_ram[310] = 19;
    exp_33_ram[311] = 19;
    exp_33_ram[312] = 147;
    exp_33_ram[313] = 147;
    exp_33_ram[314] = 51;
    exp_33_ram[315] = 19;
    exp_33_ram[316] = 147;
    exp_33_ram[317] = 147;
    exp_33_ram[318] = 99;
    exp_33_ram[319] = 179;
    exp_33_ram[320] = 99;
    exp_33_ram[321] = 19;
    exp_33_ram[322] = 103;
    exp_33_ram[323] = 99;
    exp_33_ram[324] = 179;
    exp_33_ram[325] = 227;
    exp_33_ram[326] = 99;
    exp_33_ram[327] = 179;
    exp_33_ram[328] = 147;
    exp_33_ram[329] = 99;
    exp_33_ram[330] = 51;
    exp_33_ram[331] = 99;
    exp_33_ram[332] = 99;
    exp_33_ram[333] = 99;
    exp_33_ram[334] = 99;
    exp_33_ram[335] = 99;
    exp_33_ram[336] = 19;
    exp_33_ram[337] = 103;
    exp_33_ram[338] = 19;
    exp_33_ram[339] = 99;
    exp_33_ram[340] = 19;
    exp_33_ram[341] = 103;
    exp_33_ram[342] = 99;
    exp_33_ram[343] = 227;
    exp_33_ram[344] = 103;
    exp_33_ram[345] = 227;
    exp_33_ram[346] = 99;
    exp_33_ram[347] = 227;
    exp_33_ram[348] = 227;
    exp_33_ram[349] = 19;
    exp_33_ram[350] = 103;
    exp_33_ram[351] = 19;
    exp_33_ram[352] = 103;
    exp_33_ram[353] = 227;
    exp_33_ram[354] = 111;
    exp_33_ram[355] = 227;
    exp_33_ram[356] = 111;
    exp_33_ram[357] = 227;
    exp_33_ram[358] = 227;
    exp_33_ram[359] = 147;
    exp_33_ram[360] = 111;
    exp_33_ram[361] = 19;
    exp_33_ram[362] = 35;
    exp_33_ram[363] = 35;
    exp_33_ram[364] = 19;
    exp_33_ram[365] = 99;
    exp_33_ram[366] = 239;
    exp_33_ram[367] = 19;
    exp_33_ram[368] = 147;
    exp_33_ram[369] = 51;
    exp_33_ram[370] = 99;
    exp_33_ram[371] = 147;
    exp_33_ram[372] = 179;
    exp_33_ram[373] = 19;
    exp_33_ram[374] = 179;
    exp_33_ram[375] = 51;
    exp_33_ram[376] = 131;
    exp_33_ram[377] = 19;
    exp_33_ram[378] = 147;
    exp_33_ram[379] = 3;
    exp_33_ram[380] = 19;
    exp_33_ram[381] = 147;
    exp_33_ram[382] = 179;
    exp_33_ram[383] = 147;
    exp_33_ram[384] = 19;
    exp_33_ram[385] = 103;
    exp_33_ram[386] = 147;
    exp_33_ram[387] = 179;
    exp_33_ram[388] = 19;
    exp_33_ram[389] = 111;
    exp_33_ram[390] = 147;
    exp_33_ram[391] = 19;
    exp_33_ram[392] = 111;
    exp_33_ram[393] = 19;
    exp_33_ram[394] = 35;
    exp_33_ram[395] = 35;
    exp_33_ram[396] = 35;
    exp_33_ram[397] = 35;
    exp_33_ram[398] = 35;
    exp_33_ram[399] = 35;
    exp_33_ram[400] = 179;
    exp_33_ram[401] = 99;
    exp_33_ram[402] = 19;
    exp_33_ram[403] = 19;
    exp_33_ram[404] = 147;
    exp_33_ram[405] = 99;
    exp_33_ram[406] = 19;
    exp_33_ram[407] = 239;
    exp_33_ram[408] = 147;
    exp_33_ram[409] = 19;
    exp_33_ram[410] = 51;
    exp_33_ram[411] = 147;
    exp_33_ram[412] = 99;
    exp_33_ram[413] = 19;
    exp_33_ram[414] = 147;
    exp_33_ram[415] = 99;
    exp_33_ram[416] = 19;
    exp_33_ram[417] = 99;
    exp_33_ram[418] = 147;
    exp_33_ram[419] = 19;
    exp_33_ram[420] = 179;
    exp_33_ram[421] = 179;
    exp_33_ram[422] = 179;
    exp_33_ram[423] = 179;
    exp_33_ram[424] = 179;
    exp_33_ram[425] = 131;
    exp_33_ram[426] = 3;
    exp_33_ram[427] = 147;
    exp_33_ram[428] = 19;
    exp_33_ram[429] = 147;
    exp_33_ram[430] = 51;
    exp_33_ram[431] = 131;
    exp_33_ram[432] = 3;
    exp_33_ram[433] = 131;
    exp_33_ram[434] = 3;
    exp_33_ram[435] = 19;
    exp_33_ram[436] = 147;
    exp_33_ram[437] = 19;
    exp_33_ram[438] = 103;
    exp_33_ram[439] = 239;
    exp_33_ram[440] = 147;
    exp_33_ram[441] = 111;
    exp_33_ram[442] = 147;
    exp_33_ram[443] = 179;
    exp_33_ram[444] = 147;
    exp_33_ram[445] = 111;
    exp_33_ram[446] = 147;
    exp_33_ram[447] = 99;
    exp_33_ram[448] = 19;
    exp_33_ram[449] = 19;
    exp_33_ram[450] = 147;
    exp_33_ram[451] = 239;
    exp_33_ram[452] = 51;
    exp_33_ram[453] = 19;
    exp_33_ram[454] = 179;
    exp_33_ram[455] = 147;
    exp_33_ram[456] = 19;
    exp_33_ram[457] = 51;
    exp_33_ram[458] = 239;
    exp_33_ram[459] = 51;
    exp_33_ram[460] = 19;
    exp_33_ram[461] = 19;
    exp_33_ram[462] = 147;
    exp_33_ram[463] = 147;
    exp_33_ram[464] = 99;
    exp_33_ram[465] = 19;
    exp_33_ram[466] = 99;
    exp_33_ram[467] = 19;
    exp_33_ram[468] = 179;
    exp_33_ram[469] = 19;
    exp_33_ram[470] = 51;
    exp_33_ram[471] = 51;
    exp_33_ram[472] = 179;
    exp_33_ram[473] = 179;
    exp_33_ram[474] = 55;
    exp_33_ram[475] = 19;
    exp_33_ram[476] = 179;
    exp_33_ram[477] = 19;
    exp_33_ram[478] = 99;
    exp_33_ram[479] = 19;
    exp_33_ram[480] = 147;
    exp_33_ram[481] = 99;
    exp_33_ram[482] = 19;
    exp_33_ram[483] = 179;
    exp_33_ram[484] = 179;
    exp_33_ram[485] = 147;
    exp_33_ram[486] = 55;
    exp_33_ram[487] = 51;
    exp_33_ram[488] = 99;
    exp_33_ram[489] = 55;
    exp_33_ram[490] = 19;
    exp_33_ram[491] = 19;
    exp_33_ram[492] = 179;
    exp_33_ram[493] = 51;
    exp_33_ram[494] = 147;
    exp_33_ram[495] = 19;
    exp_33_ram[496] = 179;
    exp_33_ram[497] = 147;
    exp_33_ram[498] = 111;
    exp_33_ram[499] = 147;
    exp_33_ram[500] = 179;
    exp_33_ram[501] = 147;
    exp_33_ram[502] = 111;
    exp_33_ram[503] = 147;
    exp_33_ram[504] = 147;
    exp_33_ram[505] = 19;
    exp_33_ram[506] = 111;
    exp_33_ram[507] = 19;
    exp_33_ram[508] = 19;
    exp_33_ram[509] = 147;
    exp_33_ram[510] = 99;
    exp_33_ram[511] = 51;
    exp_33_ram[512] = 147;
    exp_33_ram[513] = 19;
    exp_33_ram[514] = 227;
    exp_33_ram[515] = 103;
    exp_33_ram[516] = 99;
    exp_33_ram[517] = 99;
    exp_33_ram[518] = 19;
    exp_33_ram[519] = 147;
    exp_33_ram[520] = 19;
    exp_33_ram[521] = 99;
    exp_33_ram[522] = 147;
    exp_33_ram[523] = 99;
    exp_33_ram[524] = 99;
    exp_33_ram[525] = 19;
    exp_33_ram[526] = 147;
    exp_33_ram[527] = 227;
    exp_33_ram[528] = 19;
    exp_33_ram[529] = 99;
    exp_33_ram[530] = 179;
    exp_33_ram[531] = 51;
    exp_33_ram[532] = 147;
    exp_33_ram[533] = 19;
    exp_33_ram[534] = 227;
    exp_33_ram[535] = 103;
    exp_33_ram[536] = 147;
    exp_33_ram[537] = 239;
    exp_33_ram[538] = 19;
    exp_33_ram[539] = 103;
    exp_33_ram[540] = 51;
    exp_33_ram[541] = 99;
    exp_33_ram[542] = 179;
    exp_33_ram[543] = 111;
    exp_33_ram[544] = 179;
    exp_33_ram[545] = 147;
    exp_33_ram[546] = 239;
    exp_33_ram[547] = 51;
    exp_33_ram[548] = 103;
    exp_33_ram[549] = 147;
    exp_33_ram[550] = 99;
    exp_33_ram[551] = 99;
    exp_33_ram[552] = 239;
    exp_33_ram[553] = 19;
    exp_33_ram[554] = 103;
    exp_33_ram[555] = 179;
    exp_33_ram[556] = 227;
    exp_33_ram[557] = 51;
    exp_33_ram[558] = 239;
    exp_33_ram[559] = 51;
    exp_33_ram[560] = 103;
    exp_33_ram[561] = 99;
    exp_33_ram[562] = 147;
    exp_33_ram[563] = 179;
    exp_33_ram[564] = 99;
    exp_33_ram[565] = 19;
    exp_33_ram[566] = 19;
    exp_33_ram[567] = 51;
    exp_33_ram[568] = 147;
    exp_33_ram[569] = 103;
    exp_33_ram[570] = 51;
    exp_33_ram[571] = 51;
    exp_33_ram[572] = 179;
    exp_33_ram[573] = 51;
    exp_33_ram[574] = 111;
    exp_33_ram[575] = 99;
    exp_33_ram[576] = 147;
    exp_33_ram[577] = 179;
    exp_33_ram[578] = 99;
    exp_33_ram[579] = 147;
    exp_33_ram[580] = 19;
    exp_33_ram[581] = 179;
    exp_33_ram[582] = 19;
    exp_33_ram[583] = 103;
    exp_33_ram[584] = 51;
    exp_33_ram[585] = 179;
    exp_33_ram[586] = 51;
    exp_33_ram[587] = 179;
    exp_33_ram[588] = 111;
    exp_33_ram[589] = 183;
    exp_33_ram[590] = 99;
    exp_33_ram[591] = 147;
    exp_33_ram[592] = 179;
    exp_33_ram[593] = 147;
    exp_33_ram[594] = 55;
    exp_33_ram[595] = 147;
    exp_33_ram[596] = 179;
    exp_33_ram[597] = 51;
    exp_33_ram[598] = 147;
    exp_33_ram[599] = 51;
    exp_33_ram[600] = 3;
    exp_33_ram[601] = 51;
    exp_33_ram[602] = 103;
    exp_33_ram[603] = 55;
    exp_33_ram[604] = 147;
    exp_33_ram[605] = 227;
    exp_33_ram[606] = 147;
    exp_33_ram[607] = 111;
    exp_33_ram[608] = 115;
    exp_33_ram[609] = 97;
    exp_33_ram[610] = 46;
    exp_33_ram[611] = 108;
    exp_33_ram[612] = 72;
    exp_33_ram[613] = 111;
    exp_33_ram[614] = 49;
    exp_33_ram[615] = 105;
    exp_33_ram[616] = 50;
    exp_33_ram[617] = 105;
    exp_33_ram[618] = 72;
    exp_33_ram[619] = 51;
    exp_33_ram[620] = 105;
    exp_33_ram[621] = 52;
    exp_33_ram[622] = 105;
    exp_33_ram[623] = 112;
    exp_33_ram[624] = 0;
    exp_33_ram[625] = 115;
    exp_33_ram[626] = 99;
    exp_33_ram[627] = 46;
    exp_33_ram[628] = 108;
    exp_33_ram[629] = 121;
    exp_33_ram[630] = 109;
    exp_33_ram[631] = 109;
    exp_33_ram[632] = 46;
    exp_33_ram[633] = 115;
    exp_33_ram[634] = 109;
    exp_33_ram[635] = 46;
    exp_33_ram[636] = 115;
    exp_33_ram[637] = 99;
    exp_33_ram[638] = 46;
    exp_33_ram[639] = 109;
    exp_33_ram[640] = 104;
    exp_33_ram[641] = 46;
    exp_33_ram[642] = 53;
    exp_33_ram[643] = 105;
    exp_33_ram[644] = 115;
    exp_33_ram[645] = 104;
    exp_33_ram[646] = 46;
    exp_33_ram[647] = 54;
    exp_33_ram[648] = 105;
    exp_33_ram[649] = 115;
    exp_33_ram[650] = 115;
    exp_33_ram[651] = 46;
    exp_33_ram[652] = 97;
    exp_33_ram[653] = 49;
    exp_33_ram[654] = 97;
    exp_33_ram[655] = 97;
    exp_33_ram[656] = 50;
    exp_33_ram[657] = 97;
    exp_33_ram[658] = 97;
    exp_33_ram[659] = 51;
    exp_33_ram[660] = 97;
    exp_33_ram[661] = 115;
    exp_33_ram[662] = 0;
    exp_33_ram[663] = 97;
    exp_33_ram[664] = 97;
    exp_33_ram[665] = 0;
    exp_33_ram[666] = 115;
    exp_33_ram[667] = 98;
    exp_33_ram[668] = 46;
    exp_33_ram[669] = 97;
    exp_33_ram[670] = 97;
    exp_33_ram[671] = 0;
    exp_33_ram[672] = 97;
    exp_33_ram[673] = 97;
    exp_33_ram[674] = 108;
    exp_33_ram[675] = 108;
    exp_33_ram[676] = 52;
    exp_33_ram[677] = 102;
    exp_33_ram[678] = 97;
    exp_33_ram[679] = 97;
    exp_33_ram[680] = 0;
    exp_33_ram[681] = 115;
    exp_33_ram[682] = 99;
    exp_33_ram[683] = 46;
    exp_33_ram[684] = 115;
    exp_33_ram[685] = 112;
    exp_33_ram[686] = 46;
    exp_33_ram[687] = 97;
    exp_33_ram[688] = 52;
    exp_33_ram[689] = 97;
    exp_33_ram[690] = 102;
    exp_33_ram[691] = 100;
    exp_33_ram[692] = 97;
    exp_33_ram[693] = 49;
    exp_33_ram[694] = 100;
    exp_33_ram[695] = 97;
    exp_33_ram[696] = 102;
    exp_33_ram[697] = 115;
    exp_33_ram[698] = 0;
    exp_33_ram[699] = 115;
    exp_33_ram[700] = 116;
    exp_33_ram[701] = 46;
    exp_33_ram[702] = 49;
    exp_33_ram[703] = 0;
    exp_33_ram[704] = 50;
    exp_33_ram[705] = 51;
    exp_33_ram[706] = 109;
    exp_33_ram[707] = 101;
    exp_33_ram[708] = 46;
    exp_33_ram[709] = 97;
    exp_33_ram[710] = 0;
    exp_33_ram[711] = 98;
    exp_33_ram[712] = 0;
    exp_33_ram[713] = 99;
    exp_33_ram[714] = 0;
    exp_33_ram[715] = 100;
    exp_33_ram[716] = 0;
    exp_33_ram[717] = 115;
    exp_33_ram[718] = 101;
    exp_33_ram[719] = 46;
    exp_33_ram[720] = 116;
    exp_33_ram[721] = 46;
    exp_33_ram[722] = 84;
    exp_33_ram[723] = 83;
    exp_33_ram[724] = 49;
    exp_33_ram[725] = 48;
    exp_33_ram[726] = 58;
    exp_33_ram[727] = 50;
    exp_33_ram[728] = 10;
    exp_33_ram[729] = 84;
    exp_33_ram[730] = 83;
    exp_33_ram[731] = 49;
    exp_33_ram[732] = 49;
    exp_33_ram[733] = 58;
    exp_33_ram[734] = 50;
    exp_33_ram[735] = 10;
    exp_33_ram[736] = 55;
    exp_33_ram[737] = 105;
    exp_33_ram[738] = 56;
    exp_33_ram[739] = 105;
    exp_33_ram[740] = 57;
    exp_33_ram[741] = 105;
    exp_33_ram[742] = 84;
    exp_33_ram[743] = 83;
    exp_33_ram[744] = 49;
    exp_33_ram[745] = 50;
    exp_33_ram[746] = 58;
    exp_33_ram[747] = 50;
    exp_33_ram[748] = 10;
    exp_33_ram[749] = 49;
    exp_33_ram[750] = 97;
    exp_33_ram[751] = 49;
    exp_33_ram[752] = 97;
    exp_33_ram[753] = 49;
    exp_33_ram[754] = 97;
    exp_33_ram[755] = 0;
    exp_33_ram[756] = 3;
    exp_33_ram[757] = 4;
    exp_33_ram[758] = 4;
    exp_33_ram[759] = 5;
    exp_33_ram[760] = 5;
    exp_33_ram[761] = 5;
    exp_33_ram[762] = 5;
    exp_33_ram[763] = 6;
    exp_33_ram[764] = 6;
    exp_33_ram[765] = 6;
    exp_33_ram[766] = 6;
    exp_33_ram[767] = 6;
    exp_33_ram[768] = 6;
    exp_33_ram[769] = 6;
    exp_33_ram[770] = 6;
    exp_33_ram[771] = 7;
    exp_33_ram[772] = 7;
    exp_33_ram[773] = 7;
    exp_33_ram[774] = 7;
    exp_33_ram[775] = 7;
    exp_33_ram[776] = 7;
    exp_33_ram[777] = 7;
    exp_33_ram[778] = 7;
    exp_33_ram[779] = 7;
    exp_33_ram[780] = 7;
    exp_33_ram[781] = 7;
    exp_33_ram[782] = 7;
    exp_33_ram[783] = 7;
    exp_33_ram[784] = 7;
    exp_33_ram[785] = 7;
    exp_33_ram[786] = 7;
    exp_33_ram[787] = 8;
    exp_33_ram[788] = 8;
    exp_33_ram[789] = 8;
    exp_33_ram[790] = 8;
    exp_33_ram[791] = 8;
    exp_33_ram[792] = 8;
    exp_33_ram[793] = 8;
    exp_33_ram[794] = 8;
    exp_33_ram[795] = 8;
    exp_33_ram[796] = 8;
    exp_33_ram[797] = 8;
    exp_33_ram[798] = 8;
    exp_33_ram[799] = 8;
    exp_33_ram[800] = 8;
    exp_33_ram[801] = 8;
    exp_33_ram[802] = 8;
    exp_33_ram[803] = 8;
    exp_33_ram[804] = 8;
    exp_33_ram[805] = 8;
    exp_33_ram[806] = 8;
    exp_33_ram[807] = 8;
    exp_33_ram[808] = 8;
    exp_33_ram[809] = 8;
    exp_33_ram[810] = 8;
    exp_33_ram[811] = 8;
    exp_33_ram[812] = 8;
    exp_33_ram[813] = 8;
    exp_33_ram[814] = 8;
    exp_33_ram[815] = 8;
    exp_33_ram[816] = 8;
    exp_33_ram[817] = 8;
    exp_33_ram[818] = 8;
    exp_33_ram[819] = 147;
    exp_33_ram[820] = 19;
    exp_33_ram[821] = 51;
    exp_33_ram[822] = 3;
    exp_33_ram[823] = 99;
    exp_33_ram[824] = 103;
    exp_33_ram[825] = 19;
    exp_33_ram[826] = 35;
    exp_33_ram[827] = 111;
    exp_33_ram[828] = 19;
    exp_33_ram[829] = 183;
    exp_33_ram[830] = 35;
    exp_33_ram[831] = 3;
    exp_33_ram[832] = 35;
    exp_33_ram[833] = 147;
    exp_33_ram[834] = 239;
    exp_33_ram[835] = 147;
    exp_33_ram[836] = 131;
    exp_33_ram[837] = 35;
    exp_33_ram[838] = 3;
    exp_33_ram[839] = 19;
    exp_33_ram[840] = 19;
    exp_33_ram[841] = 103;
    exp_33_ram[842] = 179;
    exp_33_ram[843] = 147;
    exp_33_ram[844] = 147;
    exp_33_ram[845] = 99;
    exp_33_ram[846] = 19;
    exp_33_ram[847] = 51;
    exp_33_ram[848] = 19;
    exp_33_ram[849] = 111;
    exp_33_ram[850] = 131;
    exp_33_ram[851] = 19;
    exp_33_ram[852] = 147;
    exp_33_ram[853] = 35;
    exp_33_ram[854] = 131;
    exp_33_ram[855] = 35;
    exp_33_ram[856] = 131;
    exp_33_ram[857] = 35;
    exp_33_ram[858] = 131;
    exp_33_ram[859] = 35;
    exp_33_ram[860] = 179;
    exp_33_ram[861] = 227;
    exp_33_ram[862] = 19;
    exp_33_ram[863] = 19;
    exp_33_ram[864] = 179;
    exp_33_ram[865] = 179;
    exp_33_ram[866] = 19;
    exp_33_ram[867] = 51;
    exp_33_ram[868] = 99;
    exp_33_ram[869] = 19;
    exp_33_ram[870] = 19;
    exp_33_ram[871] = 179;
    exp_33_ram[872] = 179;
    exp_33_ram[873] = 147;
    exp_33_ram[874] = 99;
    exp_33_ram[875] = 103;
    exp_33_ram[876] = 51;
    exp_33_ram[877] = 131;
    exp_33_ram[878] = 51;
    exp_33_ram[879] = 147;
    exp_33_ram[880] = 35;
    exp_33_ram[881] = 111;
    exp_33_ram[882] = 51;
    exp_33_ram[883] = 3;
    exp_33_ram[884] = 51;
    exp_33_ram[885] = 147;
    exp_33_ram[886] = 35;
    exp_33_ram[887] = 111;
    exp_33_ram[888] = 147;
    exp_33_ram[889] = 3;
    exp_33_ram[890] = 99;
    exp_33_ram[891] = 51;
    exp_33_ram[892] = 3;
    exp_33_ram[893] = 99;
    exp_33_ram[894] = 3;
    exp_33_ram[895] = 99;
    exp_33_ram[896] = 103;
    exp_33_ram[897] = 147;
    exp_33_ram[898] = 111;
    exp_33_ram[899] = 227;
    exp_33_ram[900] = 147;
    exp_33_ram[901] = 147;
    exp_33_ram[902] = 163;
    exp_33_ram[903] = 111;
    exp_33_ram[904] = 35;
    exp_33_ram[905] = 103;
    exp_33_ram[906] = 179;
    exp_33_ram[907] = 147;
    exp_33_ram[908] = 99;
    exp_33_ram[909] = 183;
    exp_33_ram[910] = 55;
    exp_33_ram[911] = 147;
    exp_33_ram[912] = 19;
    exp_33_ram[913] = 3;
    exp_33_ram[914] = 131;
    exp_33_ram[915] = 99;
    exp_33_ram[916] = 131;
    exp_33_ram[917] = 3;
    exp_33_ram[918] = 99;
    exp_33_ram[919] = 99;
    exp_33_ram[920] = 51;
    exp_33_ram[921] = 103;
    exp_33_ram[922] = 51;
    exp_33_ram[923] = 147;
    exp_33_ram[924] = 179;
    exp_33_ram[925] = 179;
    exp_33_ram[926] = 99;
    exp_33_ram[927] = 19;
    exp_33_ram[928] = 147;
    exp_33_ram[929] = 111;
    exp_33_ram[930] = 19;
    exp_33_ram[931] = 147;
    exp_33_ram[932] = 111;
    exp_33_ram[933] = 19;
    exp_33_ram[934] = 103;
    exp_33_ram[935] = 147;
    exp_33_ram[936] = 19;
    exp_33_ram[937] = 51;
    exp_33_ram[938] = 3;
    exp_33_ram[939] = 99;
    exp_33_ram[940] = 103;
    exp_33_ram[941] = 19;
    exp_33_ram[942] = 111;
    exp_33_ram[943] = 147;
    exp_33_ram[944] = 99;
    exp_33_ram[945] = 103;
    exp_33_ram[946] = 51;
    exp_33_ram[947] = 35;
    exp_33_ram[948] = 147;
    exp_33_ram[949] = 111;
    exp_33_ram[950] = 147;
    exp_33_ram[951] = 51;
    exp_33_ram[952] = 99;
    exp_33_ram[953] = 19;
    exp_33_ram[954] = 111;
    exp_33_ram[955] = 19;
    exp_33_ram[956] = 3;
    exp_33_ram[957] = 147;
    exp_33_ram[958] = 227;
    exp_33_ram[959] = 103;
    exp_33_ram[960] = 19;
    exp_33_ram[961] = 35;
    exp_33_ram[962] = 35;
    exp_33_ram[963] = 19;
    exp_33_ram[964] = 35;
    exp_33_ram[965] = 147;
    exp_33_ram[966] = 239;
    exp_33_ram[967] = 147;
    exp_33_ram[968] = 51;
    exp_33_ram[969] = 99;
    exp_33_ram[970] = 19;
    exp_33_ram[971] = 111;
    exp_33_ram[972] = 19;
    exp_33_ram[973] = 131;
    exp_33_ram[974] = 147;
    exp_33_ram[975] = 227;
    exp_33_ram[976] = 131;
    exp_33_ram[977] = 3;
    exp_33_ram[978] = 131;
    exp_33_ram[979] = 19;
    exp_33_ram[980] = 103;
    exp_33_ram[981] = 19;
    exp_33_ram[982] = 35;
    exp_33_ram[983] = 35;
    exp_33_ram[984] = 19;
    exp_33_ram[985] = 35;
    exp_33_ram[986] = 147;
    exp_33_ram[987] = 239;
    exp_33_ram[988] = 147;
    exp_33_ram[989] = 179;
    exp_33_ram[990] = 99;
    exp_33_ram[991] = 19;
    exp_33_ram[992] = 111;
    exp_33_ram[993] = 19;
    exp_33_ram[994] = 3;
    exp_33_ram[995] = 147;
    exp_33_ram[996] = 227;
    exp_33_ram[997] = 131;
    exp_33_ram[998] = 3;
    exp_33_ram[999] = 131;
    exp_33_ram[1000] = 19;
    exp_33_ram[1001] = 103;
    exp_33_ram[1002] = 19;
    exp_33_ram[1003] = 35;
    exp_33_ram[1004] = 35;
    exp_33_ram[1005] = 35;
    exp_33_ram[1006] = 35;
    exp_33_ram[1007] = 35;
    exp_33_ram[1008] = 147;
    exp_33_ram[1009] = 147;
    exp_33_ram[1010] = 239;
    exp_33_ram[1011] = 19;
    exp_33_ram[1012] = 19;
    exp_33_ram[1013] = 99;
    exp_33_ram[1014] = 19;
    exp_33_ram[1015] = 239;
    exp_33_ram[1016] = 147;
    exp_33_ram[1017] = 179;
    exp_33_ram[1018] = 111;
    exp_33_ram[1019] = 51;
    exp_33_ram[1020] = 3;
    exp_33_ram[1021] = 3;
    exp_33_ram[1022] = 99;
    exp_33_ram[1023] = 147;
    exp_33_ram[1024] = 227;
    exp_33_ram[1025] = 131;
    exp_33_ram[1026] = 19;
    exp_33_ram[1027] = 3;
    exp_33_ram[1028] = 131;
    exp_33_ram[1029] = 3;
    exp_33_ram[1030] = 131;
    exp_33_ram[1031] = 19;
    exp_33_ram[1032] = 103;
    exp_33_ram[1033] = 19;
    exp_33_ram[1034] = 111;
    exp_33_ram[1035] = 19;
    exp_33_ram[1036] = 35;
    exp_33_ram[1037] = 35;
    exp_33_ram[1038] = 35;
    exp_33_ram[1039] = 35;
    exp_33_ram[1040] = 35;
    exp_33_ram[1041] = 147;
    exp_33_ram[1042] = 147;
    exp_33_ram[1043] = 239;
    exp_33_ram[1044] = 19;
    exp_33_ram[1045] = 19;
    exp_33_ram[1046] = 99;
    exp_33_ram[1047] = 19;
    exp_33_ram[1048] = 239;
    exp_33_ram[1049] = 147;
    exp_33_ram[1050] = 179;
    exp_33_ram[1051] = 111;
    exp_33_ram[1052] = 51;
    exp_33_ram[1053] = 3;
    exp_33_ram[1054] = 3;
    exp_33_ram[1055] = 99;
    exp_33_ram[1056] = 147;
    exp_33_ram[1057] = 227;
    exp_33_ram[1058] = 19;
    exp_33_ram[1059] = 111;
    exp_33_ram[1060] = 131;
    exp_33_ram[1061] = 19;
    exp_33_ram[1062] = 3;
    exp_33_ram[1063] = 131;
    exp_33_ram[1064] = 3;
    exp_33_ram[1065] = 131;
    exp_33_ram[1066] = 19;
    exp_33_ram[1067] = 103;
    exp_33_ram[1068] = 19;
    exp_33_ram[1069] = 35;
    exp_33_ram[1070] = 35;
    exp_33_ram[1071] = 35;
    exp_33_ram[1072] = 19;
    exp_33_ram[1073] = 35;
    exp_33_ram[1074] = 147;
    exp_33_ram[1075] = 239;
    exp_33_ram[1076] = 51;
    exp_33_ram[1077] = 99;
    exp_33_ram[1078] = 19;
    exp_33_ram[1079] = 239;
    exp_33_ram[1080] = 19;
    exp_33_ram[1081] = 147;
    exp_33_ram[1082] = 111;
    exp_33_ram[1083] = 179;
    exp_33_ram[1084] = 3;
    exp_33_ram[1085] = 131;
    exp_33_ram[1086] = 19;
    exp_33_ram[1087] = 99;
    exp_33_ram[1088] = 147;
    exp_33_ram[1089] = 227;
    exp_33_ram[1090] = 19;
    exp_33_ram[1091] = 111;
    exp_33_ram[1092] = 19;
    exp_33_ram[1093] = 131;
    exp_33_ram[1094] = 3;
    exp_33_ram[1095] = 131;
    exp_33_ram[1096] = 3;
    exp_33_ram[1097] = 19;
    exp_33_ram[1098] = 103;
    exp_33_ram[1099] = 19;
    exp_33_ram[1100] = 35;
    exp_33_ram[1101] = 35;
    exp_33_ram[1102] = 35;
    exp_33_ram[1103] = 35;
    exp_33_ram[1104] = 35;
    exp_33_ram[1105] = 147;
    exp_33_ram[1106] = 147;
    exp_33_ram[1107] = 239;
    exp_33_ram[1108] = 19;
    exp_33_ram[1109] = 19;
    exp_33_ram[1110] = 99;
    exp_33_ram[1111] = 19;
    exp_33_ram[1112] = 239;
    exp_33_ram[1113] = 19;
    exp_33_ram[1114] = 147;
    exp_33_ram[1115] = 51;
    exp_33_ram[1116] = 111;
    exp_33_ram[1117] = 51;
    exp_33_ram[1118] = 179;
    exp_33_ram[1119] = 3;
    exp_33_ram[1120] = 131;
    exp_33_ram[1121] = 99;
    exp_33_ram[1122] = 147;
    exp_33_ram[1123] = 227;
    exp_33_ram[1124] = 131;
    exp_33_ram[1125] = 3;
    exp_33_ram[1126] = 131;
    exp_33_ram[1127] = 3;
    exp_33_ram[1128] = 131;
    exp_33_ram[1129] = 19;
    exp_33_ram[1130] = 103;
    exp_33_ram[1131] = 19;
    exp_33_ram[1132] = 111;
    exp_33_ram[1133] = 19;
    exp_33_ram[1134] = 111;
    exp_33_ram[1135] = 147;
    exp_33_ram[1136] = 99;
    exp_33_ram[1137] = 19;
    exp_33_ram[1138] = 147;
    exp_33_ram[1139] = 35;
    exp_33_ram[1140] = 35;
    exp_33_ram[1141] = 19;
    exp_33_ram[1142] = 239;
    exp_33_ram[1143] = 147;
    exp_33_ram[1144] = 99;
    exp_33_ram[1145] = 147;
    exp_33_ram[1146] = 19;
    exp_33_ram[1147] = 239;
    exp_33_ram[1148] = 147;
    exp_33_ram[1149] = 131;
    exp_33_ram[1150] = 3;
    exp_33_ram[1151] = 19;
    exp_33_ram[1152] = 19;
    exp_33_ram[1153] = 103;
    exp_33_ram[1154] = 147;
    exp_33_ram[1155] = 19;
    exp_33_ram[1156] = 103;
    exp_33_ram[1157] = 147;
    exp_33_ram[1158] = 147;
    exp_33_ram[1159] = 99;
    exp_33_ram[1160] = 19;
    exp_33_ram[1161] = 147;
    exp_33_ram[1162] = 147;
    exp_33_ram[1163] = 99;
    exp_33_ram[1164] = 19;
    exp_33_ram[1165] = 147;
    exp_33_ram[1166] = 99;
    exp_33_ram[1167] = 19;
    exp_33_ram[1168] = 35;
    exp_33_ram[1169] = 239;
    exp_33_ram[1170] = 131;
    exp_33_ram[1171] = 179;
    exp_33_ram[1172] = 147;
    exp_33_ram[1173] = 19;
    exp_33_ram[1174] = 19;
    exp_33_ram[1175] = 103;
    exp_33_ram[1176] = 147;
    exp_33_ram[1177] = 19;
    exp_33_ram[1178] = 103;
    exp_33_ram[1179] = 183;
    exp_33_ram[1180] = 3;
    exp_33_ram[1181] = 131;
    exp_33_ram[1182] = 131;
    exp_33_ram[1183] = 19;
    exp_33_ram[1184] = 131;
    exp_33_ram[1185] = 179;
    exp_33_ram[1186] = 103;
    exp_33_ram[1187] = 147;
    exp_33_ram[1188] = 51;
    exp_33_ram[1189] = 179;
    exp_33_ram[1190] = 179;
    exp_33_ram[1191] = 19;
    exp_33_ram[1192] = 179;
    exp_33_ram[1193] = 35;
    exp_33_ram[1194] = 239;
    exp_33_ram[1195] = 131;
    exp_33_ram[1196] = 19;
    exp_33_ram[1197] = 103;
    exp_33_ram[1198] = 19;
    exp_33_ram[1199] = 35;
    exp_33_ram[1200] = 131;
    exp_33_ram[1201] = 35;
    exp_33_ram[1202] = 183;
    exp_33_ram[1203] = 35;
    exp_33_ram[1204] = 35;
    exp_33_ram[1205] = 35;
    exp_33_ram[1206] = 35;
    exp_33_ram[1207] = 35;
    exp_33_ram[1208] = 35;
    exp_33_ram[1209] = 19;
    exp_33_ram[1210] = 19;
    exp_33_ram[1211] = 19;
    exp_33_ram[1212] = 147;
    exp_33_ram[1213] = 147;
    exp_33_ram[1214] = 147;
    exp_33_ram[1215] = 99;
    exp_33_ram[1216] = 3;
    exp_33_ram[1217] = 183;
    exp_33_ram[1218] = 147;
    exp_33_ram[1219] = 147;
    exp_33_ram[1220] = 99;
    exp_33_ram[1221] = 147;
    exp_33_ram[1222] = 19;
    exp_33_ram[1223] = 239;
    exp_33_ram[1224] = 147;
    exp_33_ram[1225] = 239;
    exp_33_ram[1226] = 51;
    exp_33_ram[1227] = 179;
    exp_33_ram[1228] = 179;
    exp_33_ram[1229] = 19;
    exp_33_ram[1230] = 147;
    exp_33_ram[1231] = 111;
    exp_33_ram[1232] = 19;
    exp_33_ram[1233] = 239;
    exp_33_ram[1234] = 51;
    exp_33_ram[1235] = 147;
    exp_33_ram[1236] = 19;
    exp_33_ram[1237] = 239;
    exp_33_ram[1238] = 51;
    exp_33_ram[1239] = 179;
    exp_33_ram[1240] = 179;
    exp_33_ram[1241] = 19;
    exp_33_ram[1242] = 19;
    exp_33_ram[1243] = 111;
    exp_33_ram[1244] = 3;
    exp_33_ram[1245] = 3;
    exp_33_ram[1246] = 131;
    exp_33_ram[1247] = 147;
    exp_33_ram[1248] = 179;
    exp_33_ram[1249] = 147;
    exp_33_ram[1250] = 179;
    exp_33_ram[1251] = 19;
    exp_33_ram[1252] = 51;
    exp_33_ram[1253] = 147;
    exp_33_ram[1254] = 19;
    exp_33_ram[1255] = 3;
    exp_33_ram[1256] = 19;
    exp_33_ram[1257] = 147;
    exp_33_ram[1258] = 51;
    exp_33_ram[1259] = 179;
    exp_33_ram[1260] = 179;
    exp_33_ram[1261] = 179;
    exp_33_ram[1262] = 183;
    exp_33_ram[1263] = 147;
    exp_33_ram[1264] = 179;
    exp_33_ram[1265] = 51;
    exp_33_ram[1266] = 179;
    exp_33_ram[1267] = 147;
    exp_33_ram[1268] = 19;
    exp_33_ram[1269] = 51;
    exp_33_ram[1270] = 239;
    exp_33_ram[1271] = 179;
    exp_33_ram[1272] = 147;
    exp_33_ram[1273] = 179;
    exp_33_ram[1274] = 179;
    exp_33_ram[1275] = 51;
    exp_33_ram[1276] = 51;
    exp_33_ram[1277] = 51;
    exp_33_ram[1278] = 179;
    exp_33_ram[1279] = 131;
    exp_33_ram[1280] = 179;
    exp_33_ram[1281] = 3;
    exp_33_ram[1282] = 131;
    exp_33_ram[1283] = 3;
    exp_33_ram[1284] = 131;
    exp_33_ram[1285] = 3;
    exp_33_ram[1286] = 131;
    exp_33_ram[1287] = 3;
    exp_33_ram[1288] = 19;
    exp_33_ram[1289] = 103;
    exp_33_ram[1290] = 19;
    exp_33_ram[1291] = 35;
    exp_33_ram[1292] = 35;
    exp_33_ram[1293] = 19;
    exp_33_ram[1294] = 239;
    exp_33_ram[1295] = 183;
    exp_33_ram[1296] = 3;
    exp_33_ram[1297] = 147;
    exp_33_ram[1298] = 239;
    exp_33_ram[1299] = 183;
    exp_33_ram[1300] = 131;
    exp_33_ram[1301] = 51;
    exp_33_ram[1302] = 99;
    exp_33_ram[1303] = 35;
    exp_33_ram[1304] = 35;
    exp_33_ram[1305] = 131;
    exp_33_ram[1306] = 3;
    exp_33_ram[1307] = 147;
    exp_33_ram[1308] = 19;
    exp_33_ram[1309] = 103;
    exp_33_ram[1310] = 19;
    exp_33_ram[1311] = 35;
    exp_33_ram[1312] = 35;
    exp_33_ram[1313] = 35;
    exp_33_ram[1314] = 35;
    exp_33_ram[1315] = 147;
    exp_33_ram[1316] = 19;
    exp_33_ram[1317] = 239;
    exp_33_ram[1318] = 183;
    exp_33_ram[1319] = 3;
    exp_33_ram[1320] = 147;
    exp_33_ram[1321] = 55;
    exp_33_ram[1322] = 239;
    exp_33_ram[1323] = 51;
    exp_33_ram[1324] = 179;
    exp_33_ram[1325] = 51;
    exp_33_ram[1326] = 19;
    exp_33_ram[1327] = 51;
    exp_33_ram[1328] = 35;
    exp_33_ram[1329] = 131;
    exp_33_ram[1330] = 3;
    exp_33_ram[1331] = 35;
    exp_33_ram[1332] = 131;
    exp_33_ram[1333] = 3;
    exp_33_ram[1334] = 19;
    exp_33_ram[1335] = 103;
    exp_33_ram[1336] = 19;
    exp_33_ram[1337] = 183;
    exp_33_ram[1338] = 35;
    exp_33_ram[1339] = 19;
    exp_33_ram[1340] = 147;
    exp_33_ram[1341] = 147;
    exp_33_ram[1342] = 19;
    exp_33_ram[1343] = 35;
    exp_33_ram[1344] = 35;
    exp_33_ram[1345] = 35;
    exp_33_ram[1346] = 35;
    exp_33_ram[1347] = 35;
    exp_33_ram[1348] = 239;
    exp_33_ram[1349] = 183;
    exp_33_ram[1350] = 19;
    exp_33_ram[1351] = 147;
    exp_33_ram[1352] = 19;
    exp_33_ram[1353] = 239;
    exp_33_ram[1354] = 131;
    exp_33_ram[1355] = 183;
    exp_33_ram[1356] = 19;
    exp_33_ram[1357] = 147;
    exp_33_ram[1358] = 179;
    exp_33_ram[1359] = 147;
    exp_33_ram[1360] = 19;
    exp_33_ram[1361] = 179;
    exp_33_ram[1362] = 19;
    exp_33_ram[1363] = 19;
    exp_33_ram[1364] = 239;
    exp_33_ram[1365] = 163;
    exp_33_ram[1366] = 131;
    exp_33_ram[1367] = 19;
    exp_33_ram[1368] = 19;
    exp_33_ram[1369] = 147;
    exp_33_ram[1370] = 179;
    exp_33_ram[1371] = 147;
    exp_33_ram[1372] = 179;
    exp_33_ram[1373] = 239;
    exp_33_ram[1374] = 163;
    exp_33_ram[1375] = 3;
    exp_33_ram[1376] = 147;
    exp_33_ram[1377] = 19;
    exp_33_ram[1378] = 239;
    exp_33_ram[1379] = 35;
    exp_33_ram[1380] = 131;
    exp_33_ram[1381] = 35;
    exp_33_ram[1382] = 35;
    exp_33_ram[1383] = 147;
    exp_33_ram[1384] = 35;
    exp_33_ram[1385] = 131;
    exp_33_ram[1386] = 147;
    exp_33_ram[1387] = 147;
    exp_33_ram[1388] = 163;
    exp_33_ram[1389] = 3;
    exp_33_ram[1390] = 239;
    exp_33_ram[1391] = 35;
    exp_33_ram[1392] = 131;
    exp_33_ram[1393] = 35;
    exp_33_ram[1394] = 163;
    exp_33_ram[1395] = 147;
    exp_33_ram[1396] = 163;
    exp_33_ram[1397] = 131;
    exp_33_ram[1398] = 147;
    exp_33_ram[1399] = 147;
    exp_33_ram[1400] = 35;
    exp_33_ram[1401] = 3;
    exp_33_ram[1402] = 239;
    exp_33_ram[1403] = 35;
    exp_33_ram[1404] = 131;
    exp_33_ram[1405] = 35;
    exp_33_ram[1406] = 35;
    exp_33_ram[1407] = 147;
    exp_33_ram[1408] = 35;
    exp_33_ram[1409] = 131;
    exp_33_ram[1410] = 147;
    exp_33_ram[1411] = 147;
    exp_33_ram[1412] = 163;
    exp_33_ram[1413] = 3;
    exp_33_ram[1414] = 239;
    exp_33_ram[1415] = 35;
    exp_33_ram[1416] = 131;
    exp_33_ram[1417] = 35;
    exp_33_ram[1418] = 163;
    exp_33_ram[1419] = 147;
    exp_33_ram[1420] = 163;
    exp_33_ram[1421] = 131;
    exp_33_ram[1422] = 147;
    exp_33_ram[1423] = 147;
    exp_33_ram[1424] = 35;
    exp_33_ram[1425] = 3;
    exp_33_ram[1426] = 19;
    exp_33_ram[1427] = 239;
    exp_33_ram[1428] = 35;
    exp_33_ram[1429] = 35;
    exp_33_ram[1430] = 131;
    exp_33_ram[1431] = 3;
    exp_33_ram[1432] = 147;
    exp_33_ram[1433] = 147;
    exp_33_ram[1434] = 35;
    exp_33_ram[1435] = 239;
    exp_33_ram[1436] = 35;
    exp_33_ram[1437] = 35;
    exp_33_ram[1438] = 131;
    exp_33_ram[1439] = 3;
    exp_33_ram[1440] = 147;
    exp_33_ram[1441] = 147;
    exp_33_ram[1442] = 163;
    exp_33_ram[1443] = 239;
    exp_33_ram[1444] = 35;
    exp_33_ram[1445] = 131;
    exp_33_ram[1446] = 35;
    exp_33_ram[1447] = 131;
    exp_33_ram[1448] = 147;
    exp_33_ram[1449] = 35;
    exp_33_ram[1450] = 131;
    exp_33_ram[1451] = 131;
    exp_33_ram[1452] = 3;
    exp_33_ram[1453] = 147;
    exp_33_ram[1454] = 163;
    exp_33_ram[1455] = 147;
    exp_33_ram[1456] = 35;
    exp_33_ram[1457] = 3;
    exp_33_ram[1458] = 3;
    exp_33_ram[1459] = 19;
    exp_33_ram[1460] = 131;
    exp_33_ram[1461] = 19;
    exp_33_ram[1462] = 103;
    exp_33_ram[1463] = 19;
    exp_33_ram[1464] = 35;
    exp_33_ram[1465] = 55;
    exp_33_ram[1466] = 35;
    exp_33_ram[1467] = 35;
    exp_33_ram[1468] = 35;
    exp_33_ram[1469] = 35;
    exp_33_ram[1470] = 35;
    exp_33_ram[1471] = 35;
    exp_33_ram[1472] = 35;
    exp_33_ram[1473] = 35;
    exp_33_ram[1474] = 35;
    exp_33_ram[1475] = 35;
    exp_33_ram[1476] = 19;
    exp_33_ram[1477] = 147;
    exp_33_ram[1478] = 19;
    exp_33_ram[1479] = 147;
    exp_33_ram[1480] = 147;
    exp_33_ram[1481] = 19;
    exp_33_ram[1482] = 19;
    exp_33_ram[1483] = 239;
    exp_33_ram[1484] = 51;
    exp_33_ram[1485] = 19;
    exp_33_ram[1486] = 147;
    exp_33_ram[1487] = 19;
    exp_33_ram[1488] = 239;
    exp_33_ram[1489] = 147;
    exp_33_ram[1490] = 99;
    exp_33_ram[1491] = 99;
    exp_33_ram[1492] = 51;
    exp_33_ram[1493] = 51;
    exp_33_ram[1494] = 179;
    exp_33_ram[1495] = 147;
    exp_33_ram[1496] = 51;
    exp_33_ram[1497] = 147;
    exp_33_ram[1498] = 111;
    exp_33_ram[1499] = 55;
    exp_33_ram[1500] = 147;
    exp_33_ram[1501] = 19;
    exp_33_ram[1502] = 19;
    exp_33_ram[1503] = 147;
    exp_33_ram[1504] = 19;
    exp_33_ram[1505] = 239;
    exp_33_ram[1506] = 147;
    exp_33_ram[1507] = 19;
    exp_33_ram[1508] = 147;
    exp_33_ram[1509] = 147;
    exp_33_ram[1510] = 239;
    exp_33_ram[1511] = 99;
    exp_33_ram[1512] = 99;
    exp_33_ram[1513] = 51;
    exp_33_ram[1514] = 179;
    exp_33_ram[1515] = 179;
    exp_33_ram[1516] = 51;
    exp_33_ram[1517] = 147;
    exp_33_ram[1518] = 51;
    exp_33_ram[1519] = 111;
    exp_33_ram[1520] = 183;
    exp_33_ram[1521] = 19;
    exp_33_ram[1522] = 147;
    exp_33_ram[1523] = 239;
    exp_33_ram[1524] = 35;
    exp_33_ram[1525] = 147;
    exp_33_ram[1526] = 35;
    exp_33_ram[1527] = 51;
    exp_33_ram[1528] = 3;
    exp_33_ram[1529] = 183;
    exp_33_ram[1530] = 147;
    exp_33_ram[1531] = 239;
    exp_33_ram[1532] = 35;
    exp_33_ram[1533] = 19;
    exp_33_ram[1534] = 35;
    exp_33_ram[1535] = 3;
    exp_33_ram[1536] = 147;
    exp_33_ram[1537] = 147;
    exp_33_ram[1538] = 239;
    exp_33_ram[1539] = 147;
    exp_33_ram[1540] = 35;
    exp_33_ram[1541] = 35;
    exp_33_ram[1542] = 35;
    exp_33_ram[1543] = 35;
    exp_33_ram[1544] = 35;
    exp_33_ram[1545] = 35;
    exp_33_ram[1546] = 35;
    exp_33_ram[1547] = 51;
    exp_33_ram[1548] = 35;
    exp_33_ram[1549] = 147;
    exp_33_ram[1550] = 239;
    exp_33_ram[1551] = 35;
    exp_33_ram[1552] = 35;
    exp_33_ram[1553] = 131;
    exp_33_ram[1554] = 19;
    exp_33_ram[1555] = 3;
    exp_33_ram[1556] = 131;
    exp_33_ram[1557] = 3;
    exp_33_ram[1558] = 131;
    exp_33_ram[1559] = 3;
    exp_33_ram[1560] = 131;
    exp_33_ram[1561] = 3;
    exp_33_ram[1562] = 131;
    exp_33_ram[1563] = 3;
    exp_33_ram[1564] = 131;
    exp_33_ram[1565] = 19;
    exp_33_ram[1566] = 103;
    exp_33_ram[1567] = 19;
    exp_33_ram[1568] = 35;
    exp_33_ram[1569] = 131;
    exp_33_ram[1570] = 147;
    exp_33_ram[1571] = 35;
    exp_33_ram[1572] = 35;
    exp_33_ram[1573] = 35;
    exp_33_ram[1574] = 147;
    exp_33_ram[1575] = 19;
    exp_33_ram[1576] = 19;
    exp_33_ram[1577] = 19;
    exp_33_ram[1578] = 147;
    exp_33_ram[1579] = 19;
    exp_33_ram[1580] = 35;
    exp_33_ram[1581] = 35;
    exp_33_ram[1582] = 35;
    exp_33_ram[1583] = 35;
    exp_33_ram[1584] = 35;
    exp_33_ram[1585] = 35;
    exp_33_ram[1586] = 35;
    exp_33_ram[1587] = 35;
    exp_33_ram[1588] = 35;
    exp_33_ram[1589] = 35;
    exp_33_ram[1590] = 239;
    exp_33_ram[1591] = 19;
    exp_33_ram[1592] = 239;
    exp_33_ram[1593] = 19;
    exp_33_ram[1594] = 147;
    exp_33_ram[1595] = 19;
    exp_33_ram[1596] = 239;
    exp_33_ram[1597] = 3;
    exp_33_ram[1598] = 131;
    exp_33_ram[1599] = 19;
    exp_33_ram[1600] = 147;
    exp_33_ram[1601] = 179;
    exp_33_ram[1602] = 19;
    exp_33_ram[1603] = 35;
    exp_33_ram[1604] = 239;
    exp_33_ram[1605] = 19;
    exp_33_ram[1606] = 239;
    exp_33_ram[1607] = 147;
    exp_33_ram[1608] = 19;
    exp_33_ram[1609] = 147;
    exp_33_ram[1610] = 19;
    exp_33_ram[1611] = 19;
    exp_33_ram[1612] = 147;
    exp_33_ram[1613] = 35;
    exp_33_ram[1614] = 35;
    exp_33_ram[1615] = 35;
    exp_33_ram[1616] = 35;
    exp_33_ram[1617] = 35;
    exp_33_ram[1618] = 35;
    exp_33_ram[1619] = 239;
    exp_33_ram[1620] = 19;
    exp_33_ram[1621] = 239;
    exp_33_ram[1622] = 19;
    exp_33_ram[1623] = 147;
    exp_33_ram[1624] = 19;
    exp_33_ram[1625] = 239;
    exp_33_ram[1626] = 3;
    exp_33_ram[1627] = 131;
    exp_33_ram[1628] = 19;
    exp_33_ram[1629] = 147;
    exp_33_ram[1630] = 179;
    exp_33_ram[1631] = 19;
    exp_33_ram[1632] = 35;
    exp_33_ram[1633] = 239;
    exp_33_ram[1634] = 19;
    exp_33_ram[1635] = 239;
    exp_33_ram[1636] = 147;
    exp_33_ram[1637] = 19;
    exp_33_ram[1638] = 19;
    exp_33_ram[1639] = 147;
    exp_33_ram[1640] = 19;
    exp_33_ram[1641] = 239;
    exp_33_ram[1642] = 19;
    exp_33_ram[1643] = 239;
    exp_33_ram[1644] = 99;
    exp_33_ram[1645] = 19;
    exp_33_ram[1646] = 147;
    exp_33_ram[1647] = 99;
    exp_33_ram[1648] = 99;
    exp_33_ram[1649] = 19;
    exp_33_ram[1650] = 99;
    exp_33_ram[1651] = 99;
    exp_33_ram[1652] = 99;
    exp_33_ram[1653] = 19;
    exp_33_ram[1654] = 131;
    exp_33_ram[1655] = 3;
    exp_33_ram[1656] = 131;
    exp_33_ram[1657] = 3;
    exp_33_ram[1658] = 131;
    exp_33_ram[1659] = 3;
    exp_33_ram[1660] = 131;
    exp_33_ram[1661] = 19;
    exp_33_ram[1662] = 103;
    exp_33_ram[1663] = 19;
    exp_33_ram[1664] = 147;
    exp_33_ram[1665] = 35;
    exp_33_ram[1666] = 19;
    exp_33_ram[1667] = 19;
    exp_33_ram[1668] = 19;
    exp_33_ram[1669] = 35;
    exp_33_ram[1670] = 35;
    exp_33_ram[1671] = 35;
    exp_33_ram[1672] = 35;
    exp_33_ram[1673] = 239;
    exp_33_ram[1674] = 19;
    exp_33_ram[1675] = 147;
    exp_33_ram[1676] = 19;
    exp_33_ram[1677] = 131;
    exp_33_ram[1678] = 239;
    exp_33_ram[1679] = 19;
    exp_33_ram[1680] = 239;
    exp_33_ram[1681] = 147;
    exp_33_ram[1682] = 19;
    exp_33_ram[1683] = 99;
    exp_33_ram[1684] = 183;
    exp_33_ram[1685] = 147;
    exp_33_ram[1686] = 179;
    exp_33_ram[1687] = 51;
    exp_33_ram[1688] = 19;
    exp_33_ram[1689] = 147;
    exp_33_ram[1690] = 51;
    exp_33_ram[1691] = 147;
    exp_33_ram[1692] = 19;
    exp_33_ram[1693] = 19;
    exp_33_ram[1694] = 239;
    exp_33_ram[1695] = 19;
    exp_33_ram[1696] = 147;
    exp_33_ram[1697] = 19;
    exp_33_ram[1698] = 239;
    exp_33_ram[1699] = 99;
    exp_33_ram[1700] = 147;
    exp_33_ram[1701] = 35;
    exp_33_ram[1702] = 131;
    exp_33_ram[1703] = 147;
    exp_33_ram[1704] = 3;
    exp_33_ram[1705] = 3;
    exp_33_ram[1706] = 131;
    exp_33_ram[1707] = 19;
    exp_33_ram[1708] = 131;
    exp_33_ram[1709] = 19;
    exp_33_ram[1710] = 103;
    exp_33_ram[1711] = 227;
    exp_33_ram[1712] = 19;
    exp_33_ram[1713] = 147;
    exp_33_ram[1714] = 19;
    exp_33_ram[1715] = 239;
    exp_33_ram[1716] = 19;
    exp_33_ram[1717] = 239;
    exp_33_ram[1718] = 147;
    exp_33_ram[1719] = 99;
    exp_33_ram[1720] = 183;
    exp_33_ram[1721] = 147;
    exp_33_ram[1722] = 179;
    exp_33_ram[1723] = 51;
    exp_33_ram[1724] = 51;
    exp_33_ram[1725] = 147;
    exp_33_ram[1726] = 111;
    exp_33_ram[1727] = 99;
    exp_33_ram[1728] = 19;
    exp_33_ram[1729] = 147;
    exp_33_ram[1730] = 19;
    exp_33_ram[1731] = 239;
    exp_33_ram[1732] = 19;
    exp_33_ram[1733] = 239;
    exp_33_ram[1734] = 35;
    exp_33_ram[1735] = 111;
    exp_33_ram[1736] = 35;
    exp_33_ram[1737] = 111;
    exp_33_ram[1738] = 19;
    exp_33_ram[1739] = 19;
    exp_33_ram[1740] = 147;
    exp_33_ram[1741] = 19;
    exp_33_ram[1742] = 35;
    exp_33_ram[1743] = 239;
    exp_33_ram[1744] = 147;
    exp_33_ram[1745] = 19;
    exp_33_ram[1746] = 19;
    exp_33_ram[1747] = 239;
    exp_33_ram[1748] = 19;
    exp_33_ram[1749] = 239;
    exp_33_ram[1750] = 131;
    exp_33_ram[1751] = 19;
    exp_33_ram[1752] = 103;
    exp_33_ram[1753] = 131;
    exp_33_ram[1754] = 3;
    exp_33_ram[1755] = 19;
    exp_33_ram[1756] = 19;
    exp_33_ram[1757] = 35;
    exp_33_ram[1758] = 35;
    exp_33_ram[1759] = 239;
    exp_33_ram[1760] = 55;
    exp_33_ram[1761] = 147;
    exp_33_ram[1762] = 19;
    exp_33_ram[1763] = 19;
    exp_33_ram[1764] = 239;
    exp_33_ram[1765] = 131;
    exp_33_ram[1766] = 19;
    exp_33_ram[1767] = 3;
    exp_33_ram[1768] = 19;
    exp_33_ram[1769] = 103;
    exp_33_ram[1770] = 19;
    exp_33_ram[1771] = 35;
    exp_33_ram[1772] = 35;
    exp_33_ram[1773] = 131;
    exp_33_ram[1774] = 3;
    exp_33_ram[1775] = 35;
    exp_33_ram[1776] = 147;
    exp_33_ram[1777] = 19;
    exp_33_ram[1778] = 35;
    exp_33_ram[1779] = 35;
    exp_33_ram[1780] = 239;
    exp_33_ram[1781] = 19;
    exp_33_ram[1782] = 99;
    exp_33_ram[1783] = 55;
    exp_33_ram[1784] = 19;
    exp_33_ram[1785] = 179;
    exp_33_ram[1786] = 51;
    exp_33_ram[1787] = 51;
    exp_33_ram[1788] = 19;
    exp_33_ram[1789] = 239;
    exp_33_ram[1790] = 55;
    exp_33_ram[1791] = 147;
    exp_33_ram[1792] = 19;
    exp_33_ram[1793] = 19;
    exp_33_ram[1794] = 239;
    exp_33_ram[1795] = 19;
    exp_33_ram[1796] = 147;
    exp_33_ram[1797] = 239;
    exp_33_ram[1798] = 147;
    exp_33_ram[1799] = 35;
    exp_33_ram[1800] = 131;
    exp_33_ram[1801] = 19;
    exp_33_ram[1802] = 3;
    exp_33_ram[1803] = 131;
    exp_33_ram[1804] = 3;
    exp_33_ram[1805] = 131;
    exp_33_ram[1806] = 19;
    exp_33_ram[1807] = 103;
    exp_33_ram[1808] = 19;
    exp_33_ram[1809] = 35;
    exp_33_ram[1810] = 239;
    exp_33_ram[1811] = 131;
    exp_33_ram[1812] = 19;
    exp_33_ram[1813] = 111;
    exp_33_ram[1814] = 19;
    exp_33_ram[1815] = 35;
    exp_33_ram[1816] = 35;
    exp_33_ram[1817] = 19;
    exp_33_ram[1818] = 183;
    exp_33_ram[1819] = 19;
    exp_33_ram[1820] = 239;
    exp_33_ram[1821] = 147;
    exp_33_ram[1822] = 55;
    exp_33_ram[1823] = 19;
    exp_33_ram[1824] = 35;
    exp_33_ram[1825] = 35;
    exp_33_ram[1826] = 147;
    exp_33_ram[1827] = 19;
    exp_33_ram[1828] = 239;
    exp_33_ram[1829] = 147;
    exp_33_ram[1830] = 19;
    exp_33_ram[1831] = 147;
    exp_33_ram[1832] = 179;
    exp_33_ram[1833] = 55;
    exp_33_ram[1834] = 131;
    exp_33_ram[1835] = 147;
    exp_33_ram[1836] = 3;
    exp_33_ram[1837] = 147;
    exp_33_ram[1838] = 131;
    exp_33_ram[1839] = 19;
    exp_33_ram[1840] = 3;
    exp_33_ram[1841] = 35;
    exp_33_ram[1842] = 163;
    exp_33_ram[1843] = 35;
    exp_33_ram[1844] = 163;
    exp_33_ram[1845] = 19;
    exp_33_ram[1846] = 183;
    exp_33_ram[1847] = 147;
    exp_33_ram[1848] = 19;
    exp_33_ram[1849] = 239;
    exp_33_ram[1850] = 147;
    exp_33_ram[1851] = 99;
    exp_33_ram[1852] = 183;
    exp_33_ram[1853] = 19;
    exp_33_ram[1854] = 239;
    exp_33_ram[1855] = 111;
    exp_33_ram[1856] = 35;
    exp_33_ram[1857] = 147;
    exp_33_ram[1858] = 19;
    exp_33_ram[1859] = 239;
    exp_33_ram[1860] = 147;
    exp_33_ram[1861] = 19;
    exp_33_ram[1862] = 147;
    exp_33_ram[1863] = 179;
    exp_33_ram[1864] = 55;
    exp_33_ram[1865] = 131;
    exp_33_ram[1866] = 147;
    exp_33_ram[1867] = 3;
    exp_33_ram[1868] = 147;
    exp_33_ram[1869] = 131;
    exp_33_ram[1870] = 19;
    exp_33_ram[1871] = 3;
    exp_33_ram[1872] = 35;
    exp_33_ram[1873] = 163;
    exp_33_ram[1874] = 35;
    exp_33_ram[1875] = 163;
    exp_33_ram[1876] = 19;
    exp_33_ram[1877] = 183;
    exp_33_ram[1878] = 147;
    exp_33_ram[1879] = 19;
    exp_33_ram[1880] = 239;
    exp_33_ram[1881] = 147;
    exp_33_ram[1882] = 99;
    exp_33_ram[1883] = 183;
    exp_33_ram[1884] = 19;
    exp_33_ram[1885] = 239;
    exp_33_ram[1886] = 111;
    exp_33_ram[1887] = 147;
    exp_33_ram[1888] = 55;
    exp_33_ram[1889] = 19;
    exp_33_ram[1890] = 35;
    exp_33_ram[1891] = 35;
    exp_33_ram[1892] = 19;
    exp_33_ram[1893] = 183;
    exp_33_ram[1894] = 147;
    exp_33_ram[1895] = 19;
    exp_33_ram[1896] = 239;
    exp_33_ram[1897] = 147;
    exp_33_ram[1898] = 99;
    exp_33_ram[1899] = 183;
    exp_33_ram[1900] = 19;
    exp_33_ram[1901] = 239;
    exp_33_ram[1902] = 111;
    exp_33_ram[1903] = 35;
    exp_33_ram[1904] = 147;
    exp_33_ram[1905] = 131;
    exp_33_ram[1906] = 99;
    exp_33_ram[1907] = 183;
    exp_33_ram[1908] = 19;
    exp_33_ram[1909] = 239;
    exp_33_ram[1910] = 111;
    exp_33_ram[1911] = 183;
    exp_33_ram[1912] = 19;
    exp_33_ram[1913] = 239;
    exp_33_ram[1914] = 183;
    exp_33_ram[1915] = 19;
    exp_33_ram[1916] = 239;
    exp_33_ram[1917] = 147;
    exp_33_ram[1918] = 55;
    exp_33_ram[1919] = 19;
    exp_33_ram[1920] = 35;
    exp_33_ram[1921] = 35;
    exp_33_ram[1922] = 19;
    exp_33_ram[1923] = 19;
    exp_33_ram[1924] = 183;
    exp_33_ram[1925] = 147;
    exp_33_ram[1926] = 19;
    exp_33_ram[1927] = 239;
    exp_33_ram[1928] = 19;
    exp_33_ram[1929] = 183;
    exp_33_ram[1930] = 147;
    exp_33_ram[1931] = 19;
    exp_33_ram[1932] = 239;
    exp_33_ram[1933] = 147;
    exp_33_ram[1934] = 99;
    exp_33_ram[1935] = 183;
    exp_33_ram[1936] = 19;
    exp_33_ram[1937] = 239;
    exp_33_ram[1938] = 111;
    exp_33_ram[1939] = 35;
    exp_33_ram[1940] = 19;
    exp_33_ram[1941] = 19;
    exp_33_ram[1942] = 183;
    exp_33_ram[1943] = 147;
    exp_33_ram[1944] = 19;
    exp_33_ram[1945] = 239;
    exp_33_ram[1946] = 19;
    exp_33_ram[1947] = 183;
    exp_33_ram[1948] = 147;
    exp_33_ram[1949] = 19;
    exp_33_ram[1950] = 239;
    exp_33_ram[1951] = 147;
    exp_33_ram[1952] = 99;
    exp_33_ram[1953] = 183;
    exp_33_ram[1954] = 19;
    exp_33_ram[1955] = 239;
    exp_33_ram[1956] = 111;
    exp_33_ram[1957] = 147;
    exp_33_ram[1958] = 55;
    exp_33_ram[1959] = 19;
    exp_33_ram[1960] = 35;
    exp_33_ram[1961] = 35;
    exp_33_ram[1962] = 19;
    exp_33_ram[1963] = 183;
    exp_33_ram[1964] = 147;
    exp_33_ram[1965] = 19;
    exp_33_ram[1966] = 239;
    exp_33_ram[1967] = 147;
    exp_33_ram[1968] = 99;
    exp_33_ram[1969] = 183;
    exp_33_ram[1970] = 19;
    exp_33_ram[1971] = 239;
    exp_33_ram[1972] = 111;
    exp_33_ram[1973] = 35;
    exp_33_ram[1974] = 147;
    exp_33_ram[1975] = 131;
    exp_33_ram[1976] = 99;
    exp_33_ram[1977] = 183;
    exp_33_ram[1978] = 19;
    exp_33_ram[1979] = 239;
    exp_33_ram[1980] = 111;
    exp_33_ram[1981] = 183;
    exp_33_ram[1982] = 19;
    exp_33_ram[1983] = 239;
    exp_33_ram[1984] = 183;
    exp_33_ram[1985] = 19;
    exp_33_ram[1986] = 239;
    exp_33_ram[1987] = 183;
    exp_33_ram[1988] = 19;
    exp_33_ram[1989] = 239;
    exp_33_ram[1990] = 183;
    exp_33_ram[1991] = 19;
    exp_33_ram[1992] = 239;
    exp_33_ram[1993] = 183;
    exp_33_ram[1994] = 19;
    exp_33_ram[1995] = 239;
    exp_33_ram[1996] = 183;
    exp_33_ram[1997] = 19;
    exp_33_ram[1998] = 239;
    exp_33_ram[1999] = 183;
    exp_33_ram[2000] = 19;
    exp_33_ram[2001] = 239;
    exp_33_ram[2002] = 183;
    exp_33_ram[2003] = 19;
    exp_33_ram[2004] = 239;
    exp_33_ram[2005] = 147;
    exp_33_ram[2006] = 55;
    exp_33_ram[2007] = 19;
    exp_33_ram[2008] = 35;
    exp_33_ram[2009] = 35;
    exp_33_ram[2010] = 147;
    exp_33_ram[2011] = 19;
    exp_33_ram[2012] = 147;
    exp_33_ram[2013] = 19;
    exp_33_ram[2014] = 239;
    exp_33_ram[2015] = 19;
    exp_33_ram[2016] = 147;
    exp_33_ram[2017] = 99;
    exp_33_ram[2018] = 183;
    exp_33_ram[2019] = 19;
    exp_33_ram[2020] = 239;
    exp_33_ram[2021] = 111;
    exp_33_ram[2022] = 147;
    exp_33_ram[2023] = 19;
    exp_33_ram[2024] = 147;
    exp_33_ram[2025] = 19;
    exp_33_ram[2026] = 239;
    exp_33_ram[2027] = 19;
    exp_33_ram[2028] = 147;
    exp_33_ram[2029] = 51;
    exp_33_ram[2030] = 147;
    exp_33_ram[2031] = 99;
    exp_33_ram[2032] = 183;
    exp_33_ram[2033] = 19;
    exp_33_ram[2034] = 239;
    exp_33_ram[2035] = 111;
    exp_33_ram[2036] = 147;
    exp_33_ram[2037] = 19;
    exp_33_ram[2038] = 147;
    exp_33_ram[2039] = 19;
    exp_33_ram[2040] = 239;
    exp_33_ram[2041] = 19;
    exp_33_ram[2042] = 147;
    exp_33_ram[2043] = 51;
    exp_33_ram[2044] = 147;
    exp_33_ram[2045] = 99;
    exp_33_ram[2046] = 183;
    exp_33_ram[2047] = 19;
    exp_33_ram[2048] = 239;
    exp_33_ram[2049] = 111;
    exp_33_ram[2050] = 147;
    exp_33_ram[2051] = 19;
    exp_33_ram[2052] = 147;
    exp_33_ram[2053] = 19;
    exp_33_ram[2054] = 239;
    exp_33_ram[2055] = 19;
    exp_33_ram[2056] = 147;
    exp_33_ram[2057] = 51;
    exp_33_ram[2058] = 147;
    exp_33_ram[2059] = 99;
    exp_33_ram[2060] = 183;
    exp_33_ram[2061] = 19;
    exp_33_ram[2062] = 239;
    exp_33_ram[2063] = 111;
    exp_33_ram[2064] = 147;
    exp_33_ram[2065] = 19;
    exp_33_ram[2066] = 147;
    exp_33_ram[2067] = 19;
    exp_33_ram[2068] = 239;
    exp_33_ram[2069] = 147;
    exp_33_ram[2070] = 99;
    exp_33_ram[2071] = 183;
    exp_33_ram[2072] = 19;
    exp_33_ram[2073] = 239;
    exp_33_ram[2074] = 111;
    exp_33_ram[2075] = 183;
    exp_33_ram[2076] = 19;
    exp_33_ram[2077] = 239;
    exp_33_ram[2078] = 183;
    exp_33_ram[2079] = 19;
    exp_33_ram[2080] = 239;
    exp_33_ram[2081] = 147;
    exp_33_ram[2082] = 55;
    exp_33_ram[2083] = 19;
    exp_33_ram[2084] = 35;
    exp_33_ram[2085] = 55;
    exp_33_ram[2086] = 19;
    exp_33_ram[2087] = 35;
    exp_33_ram[2088] = 35;
    exp_33_ram[2089] = 147;
    exp_33_ram[2090] = 147;
    exp_33_ram[2091] = 19;
    exp_33_ram[2092] = 239;
    exp_33_ram[2093] = 19;
    exp_33_ram[2094] = 147;
    exp_33_ram[2095] = 99;
    exp_33_ram[2096] = 183;
    exp_33_ram[2097] = 19;
    exp_33_ram[2098] = 239;
    exp_33_ram[2099] = 111;
    exp_33_ram[2100] = 147;
    exp_33_ram[2101] = 147;
    exp_33_ram[2102] = 19;
    exp_33_ram[2103] = 239;
    exp_33_ram[2104] = 19;
    exp_33_ram[2105] = 147;
    exp_33_ram[2106] = 51;
    exp_33_ram[2107] = 147;
    exp_33_ram[2108] = 99;
    exp_33_ram[2109] = 183;
    exp_33_ram[2110] = 19;
    exp_33_ram[2111] = 239;
    exp_33_ram[2112] = 111;
    exp_33_ram[2113] = 147;
    exp_33_ram[2114] = 147;
    exp_33_ram[2115] = 19;
    exp_33_ram[2116] = 239;
    exp_33_ram[2117] = 19;
    exp_33_ram[2118] = 147;
    exp_33_ram[2119] = 51;
    exp_33_ram[2120] = 147;
    exp_33_ram[2121] = 99;
    exp_33_ram[2122] = 183;
    exp_33_ram[2123] = 19;
    exp_33_ram[2124] = 239;
    exp_33_ram[2125] = 111;
    exp_33_ram[2126] = 147;
    exp_33_ram[2127] = 147;
    exp_33_ram[2128] = 19;
    exp_33_ram[2129] = 239;
    exp_33_ram[2130] = 19;
    exp_33_ram[2131] = 147;
    exp_33_ram[2132] = 51;
    exp_33_ram[2133] = 147;
    exp_33_ram[2134] = 99;
    exp_33_ram[2135] = 183;
    exp_33_ram[2136] = 19;
    exp_33_ram[2137] = 239;
    exp_33_ram[2138] = 111;
    exp_33_ram[2139] = 147;
    exp_33_ram[2140] = 19;
    exp_33_ram[2141] = 239;
    exp_33_ram[2142] = 147;
    exp_33_ram[2143] = 19;
    exp_33_ram[2144] = 147;
    exp_33_ram[2145] = 51;
    exp_33_ram[2146] = 147;
    exp_33_ram[2147] = 51;
    exp_33_ram[2148] = 147;
    exp_33_ram[2149] = 99;
    exp_33_ram[2150] = 183;
    exp_33_ram[2151] = 19;
    exp_33_ram[2152] = 239;
    exp_33_ram[2153] = 111;
    exp_33_ram[2154] = 147;
    exp_33_ram[2155] = 147;
    exp_33_ram[2156] = 19;
    exp_33_ram[2157] = 239;
    exp_33_ram[2158] = 147;
    exp_33_ram[2159] = 99;
    exp_33_ram[2160] = 183;
    exp_33_ram[2161] = 19;
    exp_33_ram[2162] = 239;
    exp_33_ram[2163] = 111;
    exp_33_ram[2164] = 183;
    exp_33_ram[2165] = 19;
    exp_33_ram[2166] = 239;
    exp_33_ram[2167] = 183;
    exp_33_ram[2168] = 19;
    exp_33_ram[2169] = 239;
    exp_33_ram[2170] = 147;
    exp_33_ram[2171] = 55;
    exp_33_ram[2172] = 19;
    exp_33_ram[2173] = 35;
    exp_33_ram[2174] = 35;
    exp_33_ram[2175] = 19;
    exp_33_ram[2176] = 183;
    exp_33_ram[2177] = 147;
    exp_33_ram[2178] = 19;
    exp_33_ram[2179] = 239;
    exp_33_ram[2180] = 147;
    exp_33_ram[2181] = 99;
    exp_33_ram[2182] = 183;
    exp_33_ram[2183] = 19;
    exp_33_ram[2184] = 239;
    exp_33_ram[2185] = 111;
    exp_33_ram[2186] = 19;
    exp_33_ram[2187] = 183;
    exp_33_ram[2188] = 147;
    exp_33_ram[2189] = 19;
    exp_33_ram[2190] = 239;
    exp_33_ram[2191] = 19;
    exp_33_ram[2192] = 147;
    exp_33_ram[2193] = 99;
    exp_33_ram[2194] = 183;
    exp_33_ram[2195] = 19;
    exp_33_ram[2196] = 239;
    exp_33_ram[2197] = 111;
    exp_33_ram[2198] = 19;
    exp_33_ram[2199] = 183;
    exp_33_ram[2200] = 147;
    exp_33_ram[2201] = 19;
    exp_33_ram[2202] = 239;
    exp_33_ram[2203] = 19;
    exp_33_ram[2204] = 147;
    exp_33_ram[2205] = 99;
    exp_33_ram[2206] = 183;
    exp_33_ram[2207] = 19;
    exp_33_ram[2208] = 239;
    exp_33_ram[2209] = 111;
    exp_33_ram[2210] = 19;
    exp_33_ram[2211] = 183;
    exp_33_ram[2212] = 147;
    exp_33_ram[2213] = 19;
    exp_33_ram[2214] = 239;
    exp_33_ram[2215] = 19;
    exp_33_ram[2216] = 147;
    exp_33_ram[2217] = 99;
    exp_33_ram[2218] = 183;
    exp_33_ram[2219] = 19;
    exp_33_ram[2220] = 239;
    exp_33_ram[2221] = 111;
    exp_33_ram[2222] = 19;
    exp_33_ram[2223] = 183;
    exp_33_ram[2224] = 147;
    exp_33_ram[2225] = 19;
    exp_33_ram[2226] = 239;
    exp_33_ram[2227] = 19;
    exp_33_ram[2228] = 147;
    exp_33_ram[2229] = 99;
    exp_33_ram[2230] = 183;
    exp_33_ram[2231] = 19;
    exp_33_ram[2232] = 239;
    exp_33_ram[2233] = 111;
    exp_33_ram[2234] = 183;
    exp_33_ram[2235] = 19;
    exp_33_ram[2236] = 239;
    exp_33_ram[2237] = 183;
    exp_33_ram[2238] = 19;
    exp_33_ram[2239] = 239;
    exp_33_ram[2240] = 147;
    exp_33_ram[2241] = 55;
    exp_33_ram[2242] = 19;
    exp_33_ram[2243] = 35;
    exp_33_ram[2244] = 35;
    exp_33_ram[2245] = 19;
    exp_33_ram[2246] = 183;
    exp_33_ram[2247] = 147;
    exp_33_ram[2248] = 19;
    exp_33_ram[2249] = 239;
    exp_33_ram[2250] = 19;
    exp_33_ram[2251] = 147;
    exp_33_ram[2252] = 99;
    exp_33_ram[2253] = 183;
    exp_33_ram[2254] = 19;
    exp_33_ram[2255] = 239;
    exp_33_ram[2256] = 111;
    exp_33_ram[2257] = 19;
    exp_33_ram[2258] = 183;
    exp_33_ram[2259] = 147;
    exp_33_ram[2260] = 19;
    exp_33_ram[2261] = 239;
    exp_33_ram[2262] = 19;
    exp_33_ram[2263] = 147;
    exp_33_ram[2264] = 51;
    exp_33_ram[2265] = 147;
    exp_33_ram[2266] = 99;
    exp_33_ram[2267] = 183;
    exp_33_ram[2268] = 19;
    exp_33_ram[2269] = 239;
    exp_33_ram[2270] = 111;
    exp_33_ram[2271] = 19;
    exp_33_ram[2272] = 183;
    exp_33_ram[2273] = 147;
    exp_33_ram[2274] = 19;
    exp_33_ram[2275] = 239;
    exp_33_ram[2276] = 19;
    exp_33_ram[2277] = 147;
    exp_33_ram[2278] = 51;
    exp_33_ram[2279] = 147;
    exp_33_ram[2280] = 99;
    exp_33_ram[2281] = 183;
    exp_33_ram[2282] = 19;
    exp_33_ram[2283] = 239;
    exp_33_ram[2284] = 111;
    exp_33_ram[2285] = 19;
    exp_33_ram[2286] = 183;
    exp_33_ram[2287] = 147;
    exp_33_ram[2288] = 19;
    exp_33_ram[2289] = 239;
    exp_33_ram[2290] = 19;
    exp_33_ram[2291] = 147;
    exp_33_ram[2292] = 51;
    exp_33_ram[2293] = 147;
    exp_33_ram[2294] = 99;
    exp_33_ram[2295] = 183;
    exp_33_ram[2296] = 19;
    exp_33_ram[2297] = 239;
    exp_33_ram[2298] = 111;
    exp_33_ram[2299] = 19;
    exp_33_ram[2300] = 183;
    exp_33_ram[2301] = 147;
    exp_33_ram[2302] = 19;
    exp_33_ram[2303] = 239;
    exp_33_ram[2304] = 147;
    exp_33_ram[2305] = 99;
    exp_33_ram[2306] = 183;
    exp_33_ram[2307] = 19;
    exp_33_ram[2308] = 239;
    exp_33_ram[2309] = 111;
    exp_33_ram[2310] = 183;
    exp_33_ram[2311] = 19;
    exp_33_ram[2312] = 239;
    exp_33_ram[2313] = 183;
    exp_33_ram[2314] = 19;
    exp_33_ram[2315] = 239;
    exp_33_ram[2316] = 147;
    exp_33_ram[2317] = 55;
    exp_33_ram[2318] = 19;
    exp_33_ram[2319] = 35;
    exp_33_ram[2320] = 55;
    exp_33_ram[2321] = 19;
    exp_33_ram[2322] = 35;
    exp_33_ram[2323] = 35;
    exp_33_ram[2324] = 147;
    exp_33_ram[2325] = 147;
    exp_33_ram[2326] = 19;
    exp_33_ram[2327] = 239;
    exp_33_ram[2328] = 19;
    exp_33_ram[2329] = 147;
    exp_33_ram[2330] = 51;
    exp_33_ram[2331] = 147;
    exp_33_ram[2332] = 99;
    exp_33_ram[2333] = 183;
    exp_33_ram[2334] = 19;
    exp_33_ram[2335] = 239;
    exp_33_ram[2336] = 111;
    exp_33_ram[2337] = 147;
    exp_33_ram[2338] = 147;
    exp_33_ram[2339] = 19;
    exp_33_ram[2340] = 239;
    exp_33_ram[2341] = 19;
    exp_33_ram[2342] = 147;
    exp_33_ram[2343] = 51;
    exp_33_ram[2344] = 147;
    exp_33_ram[2345] = 99;
    exp_33_ram[2346] = 183;
    exp_33_ram[2347] = 19;
    exp_33_ram[2348] = 239;
    exp_33_ram[2349] = 111;
    exp_33_ram[2350] = 147;
    exp_33_ram[2351] = 147;
    exp_33_ram[2352] = 19;
    exp_33_ram[2353] = 239;
    exp_33_ram[2354] = 19;
    exp_33_ram[2355] = 147;
    exp_33_ram[2356] = 51;
    exp_33_ram[2357] = 147;
    exp_33_ram[2358] = 99;
    exp_33_ram[2359] = 183;
    exp_33_ram[2360] = 19;
    exp_33_ram[2361] = 239;
    exp_33_ram[2362] = 111;
    exp_33_ram[2363] = 147;
    exp_33_ram[2364] = 147;
    exp_33_ram[2365] = 19;
    exp_33_ram[2366] = 239;
    exp_33_ram[2367] = 19;
    exp_33_ram[2368] = 147;
    exp_33_ram[2369] = 51;
    exp_33_ram[2370] = 147;
    exp_33_ram[2371] = 99;
    exp_33_ram[2372] = 183;
    exp_33_ram[2373] = 19;
    exp_33_ram[2374] = 239;
    exp_33_ram[2375] = 111;
    exp_33_ram[2376] = 147;
    exp_33_ram[2377] = 19;
    exp_33_ram[2378] = 239;
    exp_33_ram[2379] = 147;
    exp_33_ram[2380] = 19;
    exp_33_ram[2381] = 147;
    exp_33_ram[2382] = 51;
    exp_33_ram[2383] = 147;
    exp_33_ram[2384] = 51;
    exp_33_ram[2385] = 147;
    exp_33_ram[2386] = 99;
    exp_33_ram[2387] = 183;
    exp_33_ram[2388] = 19;
    exp_33_ram[2389] = 239;
    exp_33_ram[2390] = 111;
    exp_33_ram[2391] = 147;
    exp_33_ram[2392] = 147;
    exp_33_ram[2393] = 19;
    exp_33_ram[2394] = 239;
    exp_33_ram[2395] = 147;
    exp_33_ram[2396] = 99;
    exp_33_ram[2397] = 183;
    exp_33_ram[2398] = 19;
    exp_33_ram[2399] = 239;
    exp_33_ram[2400] = 111;
    exp_33_ram[2401] = 183;
    exp_33_ram[2402] = 19;
    exp_33_ram[2403] = 239;
    exp_33_ram[2404] = 183;
    exp_33_ram[2405] = 19;
    exp_33_ram[2406] = 239;
    exp_33_ram[2407] = 147;
    exp_33_ram[2408] = 55;
    exp_33_ram[2409] = 19;
    exp_33_ram[2410] = 35;
    exp_33_ram[2411] = 35;
    exp_33_ram[2412] = 19;
    exp_33_ram[2413] = 183;
    exp_33_ram[2414] = 147;
    exp_33_ram[2415] = 19;
    exp_33_ram[2416] = 239;
    exp_33_ram[2417] = 19;
    exp_33_ram[2418] = 147;
    exp_33_ram[2419] = 99;
    exp_33_ram[2420] = 183;
    exp_33_ram[2421] = 19;
    exp_33_ram[2422] = 239;
    exp_33_ram[2423] = 111;
    exp_33_ram[2424] = 19;
    exp_33_ram[2425] = 183;
    exp_33_ram[2426] = 147;
    exp_33_ram[2427] = 19;
    exp_33_ram[2428] = 239;
    exp_33_ram[2429] = 19;
    exp_33_ram[2430] = 147;
    exp_33_ram[2431] = 99;
    exp_33_ram[2432] = 183;
    exp_33_ram[2433] = 19;
    exp_33_ram[2434] = 239;
    exp_33_ram[2435] = 111;
    exp_33_ram[2436] = 19;
    exp_33_ram[2437] = 183;
    exp_33_ram[2438] = 147;
    exp_33_ram[2439] = 19;
    exp_33_ram[2440] = 239;
    exp_33_ram[2441] = 19;
    exp_33_ram[2442] = 147;
    exp_33_ram[2443] = 99;
    exp_33_ram[2444] = 183;
    exp_33_ram[2445] = 19;
    exp_33_ram[2446] = 239;
    exp_33_ram[2447] = 111;
    exp_33_ram[2448] = 19;
    exp_33_ram[2449] = 183;
    exp_33_ram[2450] = 147;
    exp_33_ram[2451] = 19;
    exp_33_ram[2452] = 239;
    exp_33_ram[2453] = 147;
    exp_33_ram[2454] = 99;
    exp_33_ram[2455] = 183;
    exp_33_ram[2456] = 19;
    exp_33_ram[2457] = 239;
    exp_33_ram[2458] = 111;
    exp_33_ram[2459] = 19;
    exp_33_ram[2460] = 183;
    exp_33_ram[2461] = 147;
    exp_33_ram[2462] = 19;
    exp_33_ram[2463] = 239;
    exp_33_ram[2464] = 19;
    exp_33_ram[2465] = 147;
    exp_33_ram[2466] = 99;
    exp_33_ram[2467] = 183;
    exp_33_ram[2468] = 19;
    exp_33_ram[2469] = 239;
    exp_33_ram[2470] = 111;
    exp_33_ram[2471] = 183;
    exp_33_ram[2472] = 19;
    exp_33_ram[2473] = 239;
    exp_33_ram[2474] = 183;
    exp_33_ram[2475] = 19;
    exp_33_ram[2476] = 239;
    exp_33_ram[2477] = 147;
    exp_33_ram[2478] = 55;
    exp_33_ram[2479] = 19;
    exp_33_ram[2480] = 35;
    exp_33_ram[2481] = 35;
    exp_33_ram[2482] = 19;
    exp_33_ram[2483] = 183;
    exp_33_ram[2484] = 147;
    exp_33_ram[2485] = 19;
    exp_33_ram[2486] = 239;
    exp_33_ram[2487] = 19;
    exp_33_ram[2488] = 147;
    exp_33_ram[2489] = 99;
    exp_33_ram[2490] = 183;
    exp_33_ram[2491] = 19;
    exp_33_ram[2492] = 239;
    exp_33_ram[2493] = 111;
    exp_33_ram[2494] = 19;
    exp_33_ram[2495] = 183;
    exp_33_ram[2496] = 147;
    exp_33_ram[2497] = 19;
    exp_33_ram[2498] = 239;
    exp_33_ram[2499] = 19;
    exp_33_ram[2500] = 147;
    exp_33_ram[2501] = 51;
    exp_33_ram[2502] = 147;
    exp_33_ram[2503] = 99;
    exp_33_ram[2504] = 183;
    exp_33_ram[2505] = 19;
    exp_33_ram[2506] = 239;
    exp_33_ram[2507] = 111;
    exp_33_ram[2508] = 19;
    exp_33_ram[2509] = 183;
    exp_33_ram[2510] = 147;
    exp_33_ram[2511] = 19;
    exp_33_ram[2512] = 239;
    exp_33_ram[2513] = 19;
    exp_33_ram[2514] = 147;
    exp_33_ram[2515] = 51;
    exp_33_ram[2516] = 147;
    exp_33_ram[2517] = 99;
    exp_33_ram[2518] = 183;
    exp_33_ram[2519] = 19;
    exp_33_ram[2520] = 239;
    exp_33_ram[2521] = 111;
    exp_33_ram[2522] = 147;
    exp_33_ram[2523] = 147;
    exp_33_ram[2524] = 19;
    exp_33_ram[2525] = 239;
    exp_33_ram[2526] = 19;
    exp_33_ram[2527] = 147;
    exp_33_ram[2528] = 51;
    exp_33_ram[2529] = 147;
    exp_33_ram[2530] = 99;
    exp_33_ram[2531] = 183;
    exp_33_ram[2532] = 19;
    exp_33_ram[2533] = 239;
    exp_33_ram[2534] = 111;
    exp_33_ram[2535] = 19;
    exp_33_ram[2536] = 183;
    exp_33_ram[2537] = 147;
    exp_33_ram[2538] = 19;
    exp_33_ram[2539] = 239;
    exp_33_ram[2540] = 147;
    exp_33_ram[2541] = 99;
    exp_33_ram[2542] = 183;
    exp_33_ram[2543] = 19;
    exp_33_ram[2544] = 239;
    exp_33_ram[2545] = 111;
    exp_33_ram[2546] = 183;
    exp_33_ram[2547] = 19;
    exp_33_ram[2548] = 239;
    exp_33_ram[2549] = 183;
    exp_33_ram[2550] = 19;
    exp_33_ram[2551] = 239;
    exp_33_ram[2552] = 147;
    exp_33_ram[2553] = 35;
    exp_33_ram[2554] = 19;
    exp_33_ram[2555] = 183;
    exp_33_ram[2556] = 147;
    exp_33_ram[2557] = 19;
    exp_33_ram[2558] = 239;
    exp_33_ram[2559] = 147;
    exp_33_ram[2560] = 99;
    exp_33_ram[2561] = 183;
    exp_33_ram[2562] = 19;
    exp_33_ram[2563] = 239;
    exp_33_ram[2564] = 111;
    exp_33_ram[2565] = 147;
    exp_33_ram[2566] = 19;
    exp_33_ram[2567] = 147;
    exp_33_ram[2568] = 19;
    exp_33_ram[2569] = 239;
    exp_33_ram[2570] = 19;
    exp_33_ram[2571] = 183;
    exp_33_ram[2572] = 147;
    exp_33_ram[2573] = 19;
    exp_33_ram[2574] = 239;
    exp_33_ram[2575] = 147;
    exp_33_ram[2576] = 99;
    exp_33_ram[2577] = 183;
    exp_33_ram[2578] = 19;
    exp_33_ram[2579] = 239;
    exp_33_ram[2580] = 111;
    exp_33_ram[2581] = 147;
    exp_33_ram[2582] = 19;
    exp_33_ram[2583] = 147;
    exp_33_ram[2584] = 19;
    exp_33_ram[2585] = 239;
    exp_33_ram[2586] = 19;
    exp_33_ram[2587] = 183;
    exp_33_ram[2588] = 147;
    exp_33_ram[2589] = 19;
    exp_33_ram[2590] = 239;
    exp_33_ram[2591] = 147;
    exp_33_ram[2592] = 99;
    exp_33_ram[2593] = 183;
    exp_33_ram[2594] = 19;
    exp_33_ram[2595] = 239;
    exp_33_ram[2596] = 111;
    exp_33_ram[2597] = 147;
    exp_33_ram[2598] = 19;
    exp_33_ram[2599] = 147;
    exp_33_ram[2600] = 19;
    exp_33_ram[2601] = 239;
    exp_33_ram[2602] = 19;
    exp_33_ram[2603] = 183;
    exp_33_ram[2604] = 147;
    exp_33_ram[2605] = 19;
    exp_33_ram[2606] = 239;
    exp_33_ram[2607] = 147;
    exp_33_ram[2608] = 99;
    exp_33_ram[2609] = 183;
    exp_33_ram[2610] = 19;
    exp_33_ram[2611] = 239;
    exp_33_ram[2612] = 111;
    exp_33_ram[2613] = 183;
    exp_33_ram[2614] = 19;
    exp_33_ram[2615] = 239;
    exp_33_ram[2616] = 183;
    exp_33_ram[2617] = 19;
    exp_33_ram[2618] = 239;
    exp_33_ram[2619] = 183;
    exp_33_ram[2620] = 19;
    exp_33_ram[2621] = 239;
    exp_33_ram[2622] = 131;
    exp_33_ram[2623] = 3;
    exp_33_ram[2624] = 19;
    exp_33_ram[2625] = 103;
    exp_33_ram[2626] = 19;
    exp_33_ram[2627] = 35;
    exp_33_ram[2628] = 35;
    exp_33_ram[2629] = 35;
    exp_33_ram[2630] = 35;
    exp_33_ram[2631] = 35;
    exp_33_ram[2632] = 35;
    exp_33_ram[2633] = 35;
    exp_33_ram[2634] = 35;
    exp_33_ram[2635] = 19;
    exp_33_ram[2636] = 183;
    exp_33_ram[2637] = 19;
    exp_33_ram[2638] = 239;
    exp_33_ram[2639] = 147;
    exp_33_ram[2640] = 35;
    exp_33_ram[2641] = 147;
    exp_33_ram[2642] = 35;
    exp_33_ram[2643] = 147;
    exp_33_ram[2644] = 35;
    exp_33_ram[2645] = 147;
    exp_33_ram[2646] = 35;
    exp_33_ram[2647] = 147;
    exp_33_ram[2648] = 35;
    exp_33_ram[2649] = 35;
    exp_33_ram[2650] = 147;
    exp_33_ram[2651] = 35;
    exp_33_ram[2652] = 147;
    exp_33_ram[2653] = 19;
    exp_33_ram[2654] = 239;
    exp_33_ram[2655] = 19;
    exp_33_ram[2656] = 147;
    exp_33_ram[2657] = 35;
    exp_33_ram[2658] = 35;
    exp_33_ram[2659] = 147;
    exp_33_ram[2660] = 19;
    exp_33_ram[2661] = 239;
    exp_33_ram[2662] = 19;
    exp_33_ram[2663] = 183;
    exp_33_ram[2664] = 147;
    exp_33_ram[2665] = 19;
    exp_33_ram[2666] = 239;
    exp_33_ram[2667] = 147;
    exp_33_ram[2668] = 99;
    exp_33_ram[2669] = 183;
    exp_33_ram[2670] = 19;
    exp_33_ram[2671] = 239;
    exp_33_ram[2672] = 111;
    exp_33_ram[2673] = 147;
    exp_33_ram[2674] = 19;
    exp_33_ram[2675] = 239;
    exp_33_ram[2676] = 147;
    exp_33_ram[2677] = 19;
    exp_33_ram[2678] = 239;
    exp_33_ram[2679] = 19;
    exp_33_ram[2680] = 183;
    exp_33_ram[2681] = 147;
    exp_33_ram[2682] = 19;
    exp_33_ram[2683] = 239;
    exp_33_ram[2684] = 147;
    exp_33_ram[2685] = 99;
    exp_33_ram[2686] = 183;
    exp_33_ram[2687] = 19;
    exp_33_ram[2688] = 239;
    exp_33_ram[2689] = 111;
    exp_33_ram[2690] = 147;
    exp_33_ram[2691] = 19;
    exp_33_ram[2692] = 239;
    exp_33_ram[2693] = 147;
    exp_33_ram[2694] = 19;
    exp_33_ram[2695] = 239;
    exp_33_ram[2696] = 19;
    exp_33_ram[2697] = 183;
    exp_33_ram[2698] = 147;
    exp_33_ram[2699] = 19;
    exp_33_ram[2700] = 239;
    exp_33_ram[2701] = 147;
    exp_33_ram[2702] = 99;
    exp_33_ram[2703] = 183;
    exp_33_ram[2704] = 19;
    exp_33_ram[2705] = 239;
    exp_33_ram[2706] = 111;
    exp_33_ram[2707] = 147;
    exp_33_ram[2708] = 19;
    exp_33_ram[2709] = 239;
    exp_33_ram[2710] = 19;
    exp_33_ram[2711] = 183;
    exp_33_ram[2712] = 147;
    exp_33_ram[2713] = 19;
    exp_33_ram[2714] = 239;
    exp_33_ram[2715] = 147;
    exp_33_ram[2716] = 99;
    exp_33_ram[2717] = 183;
    exp_33_ram[2718] = 19;
    exp_33_ram[2719] = 239;
    exp_33_ram[2720] = 111;
    exp_33_ram[2721] = 147;
    exp_33_ram[2722] = 35;
    exp_33_ram[2723] = 147;
    exp_33_ram[2724] = 35;
    exp_33_ram[2725] = 147;
    exp_33_ram[2726] = 35;
    exp_33_ram[2727] = 147;
    exp_33_ram[2728] = 35;
    exp_33_ram[2729] = 147;
    exp_33_ram[2730] = 35;
    exp_33_ram[2731] = 35;
    exp_33_ram[2732] = 147;
    exp_33_ram[2733] = 35;
    exp_33_ram[2734] = 147;
    exp_33_ram[2735] = 19;
    exp_33_ram[2736] = 239;
    exp_33_ram[2737] = 19;
    exp_33_ram[2738] = 147;
    exp_33_ram[2739] = 35;
    exp_33_ram[2740] = 35;
    exp_33_ram[2741] = 147;
    exp_33_ram[2742] = 19;
    exp_33_ram[2743] = 239;
    exp_33_ram[2744] = 19;
    exp_33_ram[2745] = 183;
    exp_33_ram[2746] = 147;
    exp_33_ram[2747] = 19;
    exp_33_ram[2748] = 239;
    exp_33_ram[2749] = 147;
    exp_33_ram[2750] = 99;
    exp_33_ram[2751] = 183;
    exp_33_ram[2752] = 19;
    exp_33_ram[2753] = 239;
    exp_33_ram[2754] = 111;
    exp_33_ram[2755] = 147;
    exp_33_ram[2756] = 19;
    exp_33_ram[2757] = 239;
    exp_33_ram[2758] = 147;
    exp_33_ram[2759] = 19;
    exp_33_ram[2760] = 239;
    exp_33_ram[2761] = 19;
    exp_33_ram[2762] = 183;
    exp_33_ram[2763] = 147;
    exp_33_ram[2764] = 19;
    exp_33_ram[2765] = 239;
    exp_33_ram[2766] = 147;
    exp_33_ram[2767] = 99;
    exp_33_ram[2768] = 183;
    exp_33_ram[2769] = 19;
    exp_33_ram[2770] = 239;
    exp_33_ram[2771] = 111;
    exp_33_ram[2772] = 147;
    exp_33_ram[2773] = 19;
    exp_33_ram[2774] = 239;
    exp_33_ram[2775] = 147;
    exp_33_ram[2776] = 19;
    exp_33_ram[2777] = 239;
    exp_33_ram[2778] = 19;
    exp_33_ram[2779] = 183;
    exp_33_ram[2780] = 147;
    exp_33_ram[2781] = 19;
    exp_33_ram[2782] = 239;
    exp_33_ram[2783] = 147;
    exp_33_ram[2784] = 99;
    exp_33_ram[2785] = 183;
    exp_33_ram[2786] = 19;
    exp_33_ram[2787] = 239;
    exp_33_ram[2788] = 111;
    exp_33_ram[2789] = 147;
    exp_33_ram[2790] = 19;
    exp_33_ram[2791] = 239;
    exp_33_ram[2792] = 19;
    exp_33_ram[2793] = 183;
    exp_33_ram[2794] = 147;
    exp_33_ram[2795] = 19;
    exp_33_ram[2796] = 239;
    exp_33_ram[2797] = 147;
    exp_33_ram[2798] = 99;
    exp_33_ram[2799] = 183;
    exp_33_ram[2800] = 19;
    exp_33_ram[2801] = 239;
    exp_33_ram[2802] = 111;
    exp_33_ram[2803] = 147;
    exp_33_ram[2804] = 35;
    exp_33_ram[2805] = 147;
    exp_33_ram[2806] = 35;
    exp_33_ram[2807] = 147;
    exp_33_ram[2808] = 35;
    exp_33_ram[2809] = 147;
    exp_33_ram[2810] = 35;
    exp_33_ram[2811] = 147;
    exp_33_ram[2812] = 35;
    exp_33_ram[2813] = 35;
    exp_33_ram[2814] = 35;
    exp_33_ram[2815] = 147;
    exp_33_ram[2816] = 19;
    exp_33_ram[2817] = 239;
    exp_33_ram[2818] = 19;
    exp_33_ram[2819] = 147;
    exp_33_ram[2820] = 35;
    exp_33_ram[2821] = 35;
    exp_33_ram[2822] = 147;
    exp_33_ram[2823] = 19;
    exp_33_ram[2824] = 239;
    exp_33_ram[2825] = 19;
    exp_33_ram[2826] = 183;
    exp_33_ram[2827] = 147;
    exp_33_ram[2828] = 19;
    exp_33_ram[2829] = 239;
    exp_33_ram[2830] = 147;
    exp_33_ram[2831] = 99;
    exp_33_ram[2832] = 183;
    exp_33_ram[2833] = 19;
    exp_33_ram[2834] = 239;
    exp_33_ram[2835] = 111;
    exp_33_ram[2836] = 147;
    exp_33_ram[2837] = 19;
    exp_33_ram[2838] = 239;
    exp_33_ram[2839] = 147;
    exp_33_ram[2840] = 19;
    exp_33_ram[2841] = 239;
    exp_33_ram[2842] = 19;
    exp_33_ram[2843] = 183;
    exp_33_ram[2844] = 147;
    exp_33_ram[2845] = 19;
    exp_33_ram[2846] = 239;
    exp_33_ram[2847] = 147;
    exp_33_ram[2848] = 99;
    exp_33_ram[2849] = 183;
    exp_33_ram[2850] = 19;
    exp_33_ram[2851] = 239;
    exp_33_ram[2852] = 111;
    exp_33_ram[2853] = 147;
    exp_33_ram[2854] = 19;
    exp_33_ram[2855] = 239;
    exp_33_ram[2856] = 147;
    exp_33_ram[2857] = 19;
    exp_33_ram[2858] = 239;
    exp_33_ram[2859] = 19;
    exp_33_ram[2860] = 183;
    exp_33_ram[2861] = 147;
    exp_33_ram[2862] = 19;
    exp_33_ram[2863] = 239;
    exp_33_ram[2864] = 147;
    exp_33_ram[2865] = 99;
    exp_33_ram[2866] = 183;
    exp_33_ram[2867] = 19;
    exp_33_ram[2868] = 239;
    exp_33_ram[2869] = 111;
    exp_33_ram[2870] = 147;
    exp_33_ram[2871] = 19;
    exp_33_ram[2872] = 239;
    exp_33_ram[2873] = 19;
    exp_33_ram[2874] = 183;
    exp_33_ram[2875] = 147;
    exp_33_ram[2876] = 19;
    exp_33_ram[2877] = 239;
    exp_33_ram[2878] = 147;
    exp_33_ram[2879] = 99;
    exp_33_ram[2880] = 183;
    exp_33_ram[2881] = 19;
    exp_33_ram[2882] = 239;
    exp_33_ram[2883] = 111;
    exp_33_ram[2884] = 183;
    exp_33_ram[2885] = 19;
    exp_33_ram[2886] = 239;
    exp_33_ram[2887] = 147;
    exp_33_ram[2888] = 35;
    exp_33_ram[2889] = 147;
    exp_33_ram[2890] = 35;
    exp_33_ram[2891] = 147;
    exp_33_ram[2892] = 35;
    exp_33_ram[2893] = 35;
    exp_33_ram[2894] = 147;
    exp_33_ram[2895] = 35;
    exp_33_ram[2896] = 147;
    exp_33_ram[2897] = 35;
    exp_33_ram[2898] = 147;
    exp_33_ram[2899] = 35;
    exp_33_ram[2900] = 147;
    exp_33_ram[2901] = 19;
    exp_33_ram[2902] = 239;
    exp_33_ram[2903] = 19;
    exp_33_ram[2904] = 147;
    exp_33_ram[2905] = 35;
    exp_33_ram[2906] = 35;
    exp_33_ram[2907] = 3;
    exp_33_ram[2908] = 131;
    exp_33_ram[2909] = 19;
    exp_33_ram[2910] = 147;
    exp_33_ram[2911] = 239;
    exp_33_ram[2912] = 239;
    exp_33_ram[2913] = 35;
    exp_33_ram[2914] = 35;
    exp_33_ram[2915] = 35;
    exp_33_ram[2916] = 111;
    exp_33_ram[2917] = 19;
    exp_33_ram[2918] = 239;
    exp_33_ram[2919] = 19;
    exp_33_ram[2920] = 147;
    exp_33_ram[2921] = 3;
    exp_33_ram[2922] = 131;
    exp_33_ram[2923] = 19;
    exp_33_ram[2924] = 147;
    exp_33_ram[2925] = 239;
    exp_33_ram[2926] = 19;
    exp_33_ram[2927] = 147;
    exp_33_ram[2928] = 183;
    exp_33_ram[2929] = 131;
    exp_33_ram[2930] = 19;
    exp_33_ram[2931] = 239;
    exp_33_ram[2932] = 19;
    exp_33_ram[2933] = 147;
    exp_33_ram[2934] = 19;
    exp_33_ram[2935] = 147;
    exp_33_ram[2936] = 19;
    exp_33_ram[2937] = 147;
    exp_33_ram[2938] = 239;
    exp_33_ram[2939] = 147;
    exp_33_ram[2940] = 227;
    exp_33_ram[2941] = 183;
    exp_33_ram[2942] = 131;
    exp_33_ram[2943] = 19;
    exp_33_ram[2944] = 147;
    exp_33_ram[2945] = 3;
    exp_33_ram[2946] = 131;
    exp_33_ram[2947] = 51;
    exp_33_ram[2948] = 147;
    exp_33_ram[2949] = 179;
    exp_33_ram[2950] = 179;
    exp_33_ram[2951] = 179;
    exp_33_ram[2952] = 147;
    exp_33_ram[2953] = 35;
    exp_33_ram[2954] = 35;
    exp_33_ram[2955] = 19;
    exp_33_ram[2956] = 239;
    exp_33_ram[2957] = 19;
    exp_33_ram[2958] = 147;
    exp_33_ram[2959] = 35;
    exp_33_ram[2960] = 35;
    exp_33_ram[2961] = 147;
    exp_33_ram[2962] = 19;
    exp_33_ram[2963] = 239;
    exp_33_ram[2964] = 147;
    exp_33_ram[2965] = 19;
    exp_33_ram[2966] = 239;
    exp_33_ram[2967] = 131;
    exp_33_ram[2968] = 147;
    exp_33_ram[2969] = 35;
    exp_33_ram[2970] = 3;
    exp_33_ram[2971] = 147;
    exp_33_ram[2972] = 227;
    exp_33_ram[2973] = 147;
    exp_33_ram[2974] = 35;
    exp_33_ram[2975] = 147;
    exp_33_ram[2976] = 35;
    exp_33_ram[2977] = 147;
    exp_33_ram[2978] = 35;
    exp_33_ram[2979] = 147;
    exp_33_ram[2980] = 35;
    exp_33_ram[2981] = 147;
    exp_33_ram[2982] = 35;
    exp_33_ram[2983] = 147;
    exp_33_ram[2984] = 35;
    exp_33_ram[2985] = 147;
    exp_33_ram[2986] = 35;
    exp_33_ram[2987] = 147;
    exp_33_ram[2988] = 19;
    exp_33_ram[2989] = 239;
    exp_33_ram[2990] = 19;
    exp_33_ram[2991] = 147;
    exp_33_ram[2992] = 35;
    exp_33_ram[2993] = 35;
    exp_33_ram[2994] = 147;
    exp_33_ram[2995] = 19;
    exp_33_ram[2996] = 239;
    exp_33_ram[2997] = 147;
    exp_33_ram[2998] = 19;
    exp_33_ram[2999] = 239;
    exp_33_ram[3000] = 147;
    exp_33_ram[3001] = 19;
    exp_33_ram[3002] = 239;
    exp_33_ram[3003] = 147;
    exp_33_ram[3004] = 19;
    exp_33_ram[3005] = 239;
    exp_33_ram[3006] = 3;
    exp_33_ram[3007] = 131;
    exp_33_ram[3008] = 19;
    exp_33_ram[3009] = 147;
    exp_33_ram[3010] = 239;
    exp_33_ram[3011] = 19;
    exp_33_ram[3012] = 239;
    exp_33_ram[3013] = 19;
    exp_33_ram[3014] = 147;
    exp_33_ram[3015] = 35;
    exp_33_ram[3016] = 35;
    exp_33_ram[3017] = 147;
    exp_33_ram[3018] = 19;
    exp_33_ram[3019] = 239;
    exp_33_ram[3020] = 147;
    exp_33_ram[3021] = 19;
    exp_33_ram[3022] = 239;
    exp_33_ram[3023] = 239;
    exp_33_ram[3024] = 35;
    exp_33_ram[3025] = 35;
    exp_33_ram[3026] = 35;
    exp_33_ram[3027] = 111;
    exp_33_ram[3028] = 19;
    exp_33_ram[3029] = 239;
    exp_33_ram[3030] = 19;
    exp_33_ram[3031] = 147;
    exp_33_ram[3032] = 3;
    exp_33_ram[3033] = 131;
    exp_33_ram[3034] = 19;
    exp_33_ram[3035] = 147;
    exp_33_ram[3036] = 239;
    exp_33_ram[3037] = 19;
    exp_33_ram[3038] = 147;
    exp_33_ram[3039] = 183;
    exp_33_ram[3040] = 131;
    exp_33_ram[3041] = 19;
    exp_33_ram[3042] = 239;
    exp_33_ram[3043] = 19;
    exp_33_ram[3044] = 147;
    exp_33_ram[3045] = 19;
    exp_33_ram[3046] = 147;
    exp_33_ram[3047] = 19;
    exp_33_ram[3048] = 147;
    exp_33_ram[3049] = 239;
    exp_33_ram[3050] = 147;
    exp_33_ram[3051] = 227;
    exp_33_ram[3052] = 183;
    exp_33_ram[3053] = 131;
    exp_33_ram[3054] = 19;
    exp_33_ram[3055] = 147;
    exp_33_ram[3056] = 3;
    exp_33_ram[3057] = 131;
    exp_33_ram[3058] = 51;
    exp_33_ram[3059] = 147;
    exp_33_ram[3060] = 179;
    exp_33_ram[3061] = 179;
    exp_33_ram[3062] = 179;
    exp_33_ram[3063] = 147;
    exp_33_ram[3064] = 35;
    exp_33_ram[3065] = 35;
    exp_33_ram[3066] = 19;
    exp_33_ram[3067] = 239;
    exp_33_ram[3068] = 19;
    exp_33_ram[3069] = 147;
    exp_33_ram[3070] = 35;
    exp_33_ram[3071] = 35;
    exp_33_ram[3072] = 147;
    exp_33_ram[3073] = 19;
    exp_33_ram[3074] = 239;
    exp_33_ram[3075] = 147;
    exp_33_ram[3076] = 19;
    exp_33_ram[3077] = 239;
    exp_33_ram[3078] = 131;
    exp_33_ram[3079] = 147;
    exp_33_ram[3080] = 35;
    exp_33_ram[3081] = 3;
    exp_33_ram[3082] = 147;
    exp_33_ram[3083] = 227;
    exp_33_ram[3084] = 131;
    exp_33_ram[3085] = 3;
    exp_33_ram[3086] = 3;
    exp_33_ram[3087] = 131;
    exp_33_ram[3088] = 3;
    exp_33_ram[3089] = 131;
    exp_33_ram[3090] = 3;
    exp_33_ram[3091] = 131;
    exp_33_ram[3092] = 19;
    exp_33_ram[3093] = 103;
    exp_33_ram[3094] = 19;
    exp_33_ram[3095] = 35;
    exp_33_ram[3096] = 35;
    exp_33_ram[3097] = 19;
    exp_33_ram[3098] = 239;
    exp_33_ram[3099] = 239;
    exp_33_ram[3100] = 19;
    exp_33_ram[3101] = 131;
    exp_33_ram[3102] = 3;
    exp_33_ram[3103] = 19;
    exp_33_ram[3104] = 103;
    exp_33_ram[3105] = 19;
    exp_33_ram[3106] = 147;
    exp_33_ram[3107] = 51;
    exp_33_ram[3108] = 19;
    exp_33_ram[3109] = 179;
    exp_33_ram[3110] = 99;
    exp_33_ram[3111] = 99;
    exp_33_ram[3112] = 19;
    exp_33_ram[3113] = 179;
    exp_33_ram[3114] = 19;
    exp_33_ram[3115] = 103;
    exp_33_ram[3116] = 227;
    exp_33_ram[3117] = 19;
    exp_33_ram[3118] = 179;
    exp_33_ram[3119] = 111;
    exp_33_ram[3120] = 128;
    exp_33_ram[3121] = 8;
    exp_33_ram[3122] = 83;
    exp_33_ram[3123] = 111;
    exp_33_ram[3124] = 101;
    exp_33_ram[3125] = 84;
    exp_33_ram[3126] = 114;
    exp_33_ram[3127] = 116;
    exp_33_ram[3128] = 74;
    exp_33_ram[3129] = 101;
    exp_33_ram[3130] = 114;
    exp_33_ram[3131] = 77;
    exp_33_ram[3132] = 117;
    exp_33_ram[3133] = 108;
    exp_33_ram[3134] = 83;
    exp_33_ram[3135] = 99;
    exp_33_ram[3136] = 118;
    exp_33_ram[3137] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_179;

  reg [31:0] exp_179_reg;
  always@(*) begin
    case (exp_177)
      0:exp_179_reg <= exp_157;
      1:exp_179_reg <= exp_167;
      default:exp_179_reg <= exp_178;
    endcase
  end
  assign exp_179 = exp_179_reg;
  assign exp_177 = exp_139[2:2];
  assign exp_139 = exp_1;
  assign exp_178 = 0;

      reg [31:0] exp_157_reg = 0;
      always@(posedge clk) begin
        if (exp_156) begin
          exp_157_reg <= exp_164;
        end
      end
      assign exp_157 = exp_157_reg;
    
  reg [31:0] exp_164_reg;
  always@(*) begin
    case (exp_159)
      0:exp_164_reg <= exp_161;
      1:exp_164_reg <= exp_162;
      default:exp_164_reg <= exp_163;
    endcase
  end
  assign exp_164 = exp_164_reg;
  assign exp_159 = exp_157 == exp_158;
  assign exp_158 = 4294967295;
  assign exp_163 = 0;
  assign exp_161 = exp_157 + exp_160;
  assign exp_160 = 1;
  assign exp_162 = 0;
  assign exp_156 = 1;

      reg [31:0] exp_167_reg = 0;
      always@(posedge clk) begin
        if (exp_166) begin
          exp_167_reg <= exp_174;
        end
      end
      assign exp_167 = exp_167_reg;
    
  reg [31:0] exp_174_reg;
  always@(*) begin
    case (exp_169)
      0:exp_174_reg <= exp_171;
      1:exp_174_reg <= exp_172;
      default:exp_174_reg <= exp_173;
    endcase
  end
  assign exp_174 = exp_174_reg;
  assign exp_169 = exp_167 == exp_168;
  assign exp_168 = 4294967295;
  assign exp_173 = 0;
  assign exp_171 = exp_167 + exp_170;
  assign exp_170 = 1;
  assign exp_172 = 0;
  assign exp_166 = exp_159 & exp_165;
  assign exp_165 = 1;
  assign exp_182 = exp_201;
  assign exp_201 = 0;
  assign exp_204 = exp_222;
  assign exp_222 = 0;
  assign exp_226 = exp_241;
  assign exp_241 = stdin_in;
  assign exp_461 = exp_248[15:8];
  assign exp_462 = exp_248[23:16];
  assign exp_463 = exp_248[31:24];
  assign exp_475 = $signed(exp_474);
  assign exp_474 = exp_473 + exp_469;
  assign exp_473 = 0;

  reg [15:0] exp_469_reg;
  always@(*) begin
    case (exp_459)
      0:exp_469_reg <= exp_466;
      1:exp_469_reg <= exp_467;
      default:exp_469_reg <= exp_468;
    endcase
  end
  assign exp_469 = exp_469_reg;
  assign exp_468 = 0;
  assign exp_466 = exp_248[15:0];
  assign exp_467 = exp_248[31:16];
  assign exp_476 = 0;
  assign exp_477 = exp_465;
  assign exp_478 = exp_469;
  assign exp_479 = 0;
  assign exp_480 = 0;

  reg [31:0] exp_839_reg;
  always@(*) begin
    case (exp_629)
      0:exp_839_reg <= exp_835;
      1:exp_839_reg <= exp_837;
      default:exp_839_reg <= exp_838;
    endcase
  end
  assign exp_839 = exp_839_reg;
  assign exp_838 = 0;

  reg [31:0] exp_835_reg;
  always@(*) begin
    case (exp_606)
      0:exp_835_reg <= exp_830;
      1:exp_835_reg <= exp_831;
      default:exp_835_reg <= exp_834;
    endcase
  end
  assign exp_835 = exp_835_reg;
  assign exp_606 = exp_605 & exp_603;
  assign exp_605 = exp_598 == exp_604;
  assign exp_604 = 0;
  assign exp_834 = 0;
  assign exp_830 = exp_829[63:32];

  reg [63:0] exp_829_reg;
  always@(*) begin
    case (exp_826)
      0:exp_829_reg <= exp_825;
      1:exp_829_reg <= exp_827;
      default:exp_829_reg <= exp_828;
    endcase
  end
  assign exp_829 = exp_829_reg;

      reg [0:0] exp_826_reg = 0;
      always@(posedge clk) begin
        if (exp_811) begin
          exp_826_reg <= exp_809;
        end
      end
      assign exp_826 = exp_826_reg;
    
      reg [0:0] exp_809_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_809_reg <= exp_786;
        end
      end
      assign exp_809 = exp_809_reg;
    
      reg [0:0] exp_786_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_786_reg <= exp_783;
        end
      end
      assign exp_786 = exp_786_reg;
      assign exp_783 = exp_781 ^ exp_782;
  assign exp_781 = exp_763 & exp_746;
  assign exp_763 = exp_762 + exp_761;
  assign exp_762 = 0;
  assign exp_761 = exp_759[31:31];

      reg [31:0] exp_759_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_759_reg <= exp_376;
        end
      end
      assign exp_759 = exp_759_reg;
      assign exp_758 = exp_748 == exp_757;
  assign exp_757 = 0;
  assign exp_746 = exp_745 | exp_612;
  assign exp_745 = exp_606 | exp_609;
  assign exp_609 = exp_608 & exp_603;
  assign exp_608 = exp_598 == exp_607;
  assign exp_607 = 1;
  assign exp_612 = exp_611 & exp_603;
  assign exp_611 = exp_598 == exp_610;
  assign exp_610 = 2;
  assign exp_782 = exp_766 & exp_747;
  assign exp_766 = exp_765 + exp_764;
  assign exp_765 = 0;
  assign exp_764 = exp_760[31:31];

      reg [31:0] exp_760_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_760_reg <= exp_377;
        end
      end
      assign exp_760 = exp_760_reg;
      assign exp_747 = exp_606 | exp_609;
  assign exp_768 = exp_748 == exp_767;
  assign exp_767 = 1;
  assign exp_788 = exp_748 == exp_787;
  assign exp_787 = 2;
  assign exp_811 = exp_748 == exp_810;
  assign exp_810 = 3;
  assign exp_828 = 0;

      reg [63:0] exp_825_reg = 0;
      always@(posedge clk) begin
        if (exp_811) begin
          exp_825_reg <= exp_824;
        end
      end
      assign exp_825 = exp_825_reg;
      assign exp_824 = exp_820 + exp_823;
  assign exp_820 = exp_816 + exp_819;
  assign exp_816 = exp_812 + exp_815;
  assign exp_812 = exp_805;

      reg [31:0] exp_805_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_805_reg <= exp_792;
        end
      end
      assign exp_805 = exp_805_reg;
      assign exp_792 = exp_790 * exp_791;
  assign exp_790 = exp_789;
  assign exp_789 = exp_784[15:0];

      reg [31:0] exp_784_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_784_reg <= exp_774;
        end
      end
      assign exp_784 = exp_784_reg;
      assign exp_774 = exp_773 + exp_772;
  assign exp_773 = 0;

  reg [31:0] exp_772_reg;
  always@(*) begin
    case (exp_769)
      0:exp_772_reg <= exp_759;
      1:exp_772_reg <= exp_770;
      default:exp_772_reg <= exp_771;
    endcase
  end
  assign exp_772 = exp_772_reg;
  assign exp_769 = exp_763 & exp_746;
  assign exp_771 = 0;
  assign exp_770 = -exp_759;
  assign exp_791 = exp_785[15:0];

      reg [31:0] exp_785_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_785_reg <= exp_780;
        end
      end
      assign exp_785 = exp_785_reg;
      assign exp_780 = exp_779 + exp_778;
  assign exp_779 = 0;

  reg [31:0] exp_778_reg;
  always@(*) begin
    case (exp_775)
      0:exp_778_reg <= exp_760;
      1:exp_778_reg <= exp_776;
      default:exp_778_reg <= exp_777;
    endcase
  end
  assign exp_778 = exp_778_reg;
  assign exp_775 = exp_766 & exp_747;
  assign exp_777 = 0;
  assign exp_776 = -exp_760;
  assign exp_815 = exp_813 << exp_814;
  assign exp_813 = exp_806;

      reg [31:0] exp_806_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_806_reg <= exp_796;
        end
      end
      assign exp_806 = exp_806_reg;
      assign exp_796 = exp_794 * exp_795;
  assign exp_794 = exp_793;
  assign exp_793 = exp_784[15:0];
  assign exp_795 = exp_785[31:16];
  assign exp_814 = 16;
  assign exp_819 = exp_817 << exp_818;
  assign exp_817 = exp_807;

      reg [31:0] exp_807_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_807_reg <= exp_800;
        end
      end
      assign exp_807 = exp_807_reg;
      assign exp_800 = exp_798 * exp_799;
  assign exp_798 = exp_797;
  assign exp_797 = exp_784[31:16];
  assign exp_799 = exp_785[15:0];
  assign exp_818 = 16;
  assign exp_823 = exp_821 << exp_822;
  assign exp_821 = exp_808;

      reg [31:0] exp_808_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_808_reg <= exp_804;
        end
      end
      assign exp_808 = exp_808_reg;
      assign exp_804 = exp_802 * exp_803;
  assign exp_802 = exp_801;
  assign exp_801 = exp_784[31:16];
  assign exp_803 = exp_785[31:16];
  assign exp_822 = 32;
  assign exp_827 = -exp_825;
  assign exp_831 = exp_829[31:0];

  reg [31:0] exp_837_reg;
  always@(*) begin
    case (exp_630)
      0:exp_837_reg <= exp_740;
      1:exp_837_reg <= exp_741;
      default:exp_837_reg <= exp_836;
    endcase
  end
  assign exp_837 = exp_837_reg;
  assign exp_630 = exp_598[1:1];
  assign exp_836 = 0;

      reg [31:0] exp_740_reg = 0;
      always@(posedge clk) begin
        if (exp_649) begin
          exp_740_reg <= exp_734;
        end
      end
      assign exp_740 = exp_740_reg;
    
  reg [31:0] exp_734_reg;
  always@(*) begin
    case (exp_730)
      0:exp_734_reg <= exp_721;
      1:exp_734_reg <= exp_732;
      default:exp_734_reg <= exp_733;
    endcase
  end
  assign exp_734 = exp_734_reg;
  assign exp_730 = exp_729 & exp_632;
  assign exp_729 = exp_678 == exp_728;

      reg [31:0] exp_678_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_678_reg <= exp_675;
        end
      end
      assign exp_678 = exp_678_reg;
      assign exp_675 = exp_674 + exp_673;
  assign exp_674 = 0;

  reg [31:0] exp_673_reg;
  always@(*) begin
    case (exp_670)
      0:exp_673_reg <= exp_655;
      1:exp_673_reg <= exp_671;
      default:exp_673_reg <= exp_672;
    endcase
  end
  assign exp_673 = exp_673_reg;
  assign exp_670 = exp_661 & exp_632;
  assign exp_661 = exp_660 + exp_659;
  assign exp_660 = 0;
  assign exp_659 = exp_655[31:31];

      reg [31:0] exp_655_reg = 0;
      always@(posedge clk) begin
        if (exp_653) begin
          exp_655_reg <= exp_377;
        end
      end
      assign exp_655 = exp_655_reg;
      assign exp_653 = exp_635 == exp_652;
  assign exp_652 = 0;
  assign exp_632 = ~exp_631;
  assign exp_631 = exp_598[0:0];
  assign exp_672 = 0;
  assign exp_671 = -exp_655;
  assign exp_663 = exp_635 == exp_662;
  assign exp_662 = 1;
  assign exp_728 = 0;
  assign exp_733 = 0;
  assign exp_721 = exp_720 + exp_719;
  assign exp_720 = 0;

  reg [31:0] exp_719_reg;
  always@(*) begin
    case (exp_716)
      0:exp_719_reg <= exp_714;
      1:exp_719_reg <= exp_717;
      default:exp_719_reg <= exp_718;
    endcase
  end
  assign exp_719 = exp_719_reg;
  assign exp_716 = exp_680 & exp_632;

      reg [0:0] exp_680_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_680_reg <= exp_676;
        end
      end
      assign exp_680 = exp_680_reg;
      assign exp_676 = exp_658 ^ exp_661;
  assign exp_658 = exp_657 + exp_656;
  assign exp_657 = 0;
  assign exp_656 = exp_654[31:31];

      reg [31:0] exp_654_reg = 0;
      always@(posedge clk) begin
        if (exp_653) begin
          exp_654_reg <= exp_376;
        end
      end
      assign exp_654 = exp_654_reg;
      assign exp_718 = 0;

      reg [31:0] exp_714_reg = 0;
      always@(posedge clk) begin
        if (exp_647) begin
          exp_714_reg <= exp_684;
        end
      end
      assign exp_714 = exp_714_reg;
    
      reg [31:0] exp_684_reg = 0;
      always@(posedge clk) begin
        if (exp_683) begin
          exp_684_reg <= exp_711;
        end
      end
      assign exp_684 = exp_684_reg;
    
  reg [31:0] exp_711_reg;
  always@(*) begin
    case (exp_645)
      0:exp_711_reg <= exp_703;
      1:exp_711_reg <= exp_709;
      default:exp_711_reg <= exp_710;
    endcase
  end
  assign exp_711 = exp_711_reg;
  assign exp_645 = exp_635 == exp_644;
  assign exp_644 = 2;
  assign exp_710 = 0;

  reg [31:0] exp_703_reg;
  always@(*) begin
    case (exp_693)
      0:exp_703_reg <= exp_697;
      1:exp_703_reg <= exp_701;
      default:exp_703_reg <= exp_702;
    endcase
  end
  assign exp_703 = exp_703_reg;
  assign exp_693 = ~exp_692;
  assign exp_692 = exp_691[32:32];
  assign exp_691 = exp_690 - exp_678;
  assign exp_690 = exp_689;
  assign exp_689 = {exp_687, exp_688};  assign exp_687 = exp_682[31:0];

      reg [31:0] exp_682_reg = 0;
      always@(posedge clk) begin
        if (exp_681) begin
          exp_682_reg <= exp_708;
        end
      end
      assign exp_682 = exp_682_reg;
    
  reg [32:0] exp_708_reg;
  always@(*) begin
    case (exp_645)
      0:exp_708_reg <= exp_695;
      1:exp_708_reg <= exp_706;
      default:exp_708_reg <= exp_707;
    endcase
  end
  assign exp_708 = exp_708_reg;
  assign exp_707 = 0;

  reg [32:0] exp_695_reg;
  always@(*) begin
    case (exp_693)
      0:exp_695_reg <= exp_689;
      1:exp_695_reg <= exp_691;
      default:exp_695_reg <= exp_694;
    endcase
  end
  assign exp_695 = exp_695_reg;
  assign exp_694 = 0;
  assign exp_706 = 0;
  assign exp_681 = 1;
  assign exp_688 = exp_686[31:31];

      reg [31:0] exp_686_reg = 0;
      always@(posedge clk) begin
        if (exp_685) begin
          exp_686_reg <= exp_713;
        end
      end
      assign exp_686 = exp_686_reg;
    
  reg [31:0] exp_713_reg;
  always@(*) begin
    case (exp_645)
      0:exp_713_reg <= exp_705;
      1:exp_713_reg <= exp_677;
      default:exp_713_reg <= exp_712;
    endcase
  end
  assign exp_713 = exp_713_reg;
  assign exp_712 = 0;
  assign exp_705 = exp_686 << exp_704;
  assign exp_704 = 1;

      reg [31:0] exp_677_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_677_reg <= exp_669;
        end
      end
      assign exp_677 = exp_677_reg;
      assign exp_669 = exp_668 + exp_667;
  assign exp_668 = 0;

  reg [31:0] exp_667_reg;
  always@(*) begin
    case (exp_664)
      0:exp_667_reg <= exp_654;
      1:exp_667_reg <= exp_665;
      default:exp_667_reg <= exp_666;
    endcase
  end
  assign exp_667 = exp_667_reg;
  assign exp_664 = exp_658 & exp_632;
  assign exp_666 = 0;
  assign exp_665 = -exp_654;
  assign exp_685 = 1;
  assign exp_702 = 0;
  assign exp_697 = exp_684 << exp_696;
  assign exp_696 = 1;
  assign exp_701 = exp_699 | exp_700;
  assign exp_699 = exp_684 << exp_698;
  assign exp_698 = 1;
  assign exp_700 = 1;
  assign exp_709 = 0;
  assign exp_683 = 1;
  assign exp_647 = exp_635 == exp_646;
  assign exp_646 = 35;
  assign exp_717 = -exp_714;
  assign exp_732 = $signed(exp_731);
  assign exp_731 = -1;
  assign exp_649 = exp_635 == exp_648;
  assign exp_648 = 36;

      reg [31:0] exp_741_reg = 0;
      always@(posedge clk) begin
        if (exp_649) begin
          exp_741_reg <= exp_739;
        end
      end
      assign exp_741 = exp_741_reg;
    
  reg [31:0] exp_739_reg;
  always@(*) begin
    case (exp_737)
      0:exp_739_reg <= exp_727;
      1:exp_739_reg <= exp_654;
      default:exp_739_reg <= exp_738;
    endcase
  end
  assign exp_739 = exp_739_reg;
  assign exp_737 = exp_736 & exp_632;
  assign exp_736 = exp_678 == exp_735;
  assign exp_735 = 0;
  assign exp_738 = 0;
  assign exp_727 = exp_726 + exp_725;
  assign exp_726 = 0;

  reg [31:0] exp_725_reg;
  always@(*) begin
    case (exp_722)
      0:exp_725_reg <= exp_715;
      1:exp_725_reg <= exp_723;
      default:exp_725_reg <= exp_724;
    endcase
  end
  assign exp_725 = exp_725_reg;
  assign exp_722 = exp_679 & exp_632;

      reg [0:0] exp_679_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_679_reg <= exp_658;
        end
      end
      assign exp_679 = exp_679_reg;
      assign exp_724 = 0;

      reg [31:0] exp_715_reg = 0;
      always@(posedge clk) begin
        if (exp_647) begin
          exp_715_reg <= exp_682;
        end
      end
      assign exp_715 = exp_715_reg;
      assign exp_723 = -exp_715;
  assign exp_310 = $signed(exp_309);
  assign exp_309 = 0;
  assign exp_539 = exp_374 != exp_375;
  assign exp_552 = 0;
  assign exp_553 = 0;
  assign exp_540 = $signed(exp_374) < $signed(exp_375);
  assign exp_541 = $signed(exp_374) >= $signed(exp_375);
  assign exp_546 = exp_543 < exp_545;
  assign exp_543 = exp_542 + exp_374;
  assign exp_542 = 0;
  assign exp_545 = exp_544 + exp_375;
  assign exp_544 = 0;
  assign exp_551 = exp_548 >= exp_550;
  assign exp_548 = exp_547 + exp_374;
  assign exp_547 = 0;
  assign exp_550 = exp_549 + exp_375;
  assign exp_549 = 0;
  assign exp_866 = 0;
  assign exp_865 = exp_264 + exp_864;
  assign exp_864 = 4;

  reg [32:0] exp_596_reg;
  always@(*) begin
    case (exp_397)
      0:exp_596_reg <= exp_586;
      1:exp_596_reg <= exp_594;
      default:exp_596_reg <= exp_595;
    endcase
  end
  assign exp_596 = exp_596_reg;
  assign exp_595 = 0;
  assign exp_586 = exp_585 + exp_383;

  reg [31:0] exp_585_reg;
  always@(*) begin
    case (exp_395)
      0:exp_585_reg <= exp_571;
      1:exp_585_reg <= exp_583;
      default:exp_585_reg <= exp_584;
    endcase
  end
  assign exp_585 = exp_585_reg;
  assign exp_584 = 0;
  assign exp_571 = $signed(exp_570);
  assign exp_570 = exp_569 + exp_568;
  assign exp_569 = 0;
  assign exp_568 = {exp_567, exp_564};  assign exp_567 = {exp_566, exp_563};  assign exp_566 = {exp_565, exp_562};  assign exp_565 = {exp_560, exp_561};  assign exp_560 = exp_382[31:31];
  assign exp_561 = exp_382[7:7];
  assign exp_562 = exp_382[30:25];
  assign exp_563 = exp_382[11:8];
  assign exp_564 = 0;
  assign exp_583 = $signed(exp_582);
  assign exp_582 = exp_581 + exp_580;
  assign exp_581 = 0;
  assign exp_580 = {exp_579, exp_576};  assign exp_579 = {exp_578, exp_575};  assign exp_578 = {exp_577, exp_574};  assign exp_577 = {exp_572, exp_573};  assign exp_572 = exp_382[31:31];
  assign exp_573 = exp_382[19:12];
  assign exp_574 = exp_382[20:20];
  assign exp_575 = exp_382[30:21];
  assign exp_576 = 0;

      reg [31:0] exp_383_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_383_reg <= exp_266;
        end
      end
      assign exp_383 = exp_383_reg;
      assign exp_594 = exp_593 & exp_592;
  assign exp_593 = $signed(exp_591);
  assign exp_591 = exp_374 + exp_590;
  assign exp_590 = $signed(exp_589);
  assign exp_589 = exp_588 + exp_587;
  assign exp_588 = 0;
  assign exp_587 = exp_382[31:20];
  assign exp_592 = 4294967294;
  assign exp_263 = exp_256 & exp_254;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_265;
  assign exp_398 = 3;
  assign exp_244 = ~exp_229;
  assign exp_229 = exp_6;
  assign exp_200 = exp_184 & exp_185;
  assign exp_184 = exp_192;
  assign exp_192 = exp_5 & exp_191;
  assign exp_185 = exp_6;
  assign exp_181 = exp_2;

      reg [31:0] exp_221_reg = 0;
      always@(posedge clk) begin
        if (exp_220) begin
          exp_221_reg <= exp_203;
        end
      end
      assign exp_221 = exp_221_reg;
      assign exp_203 = exp_2;
  assign exp_220 = exp_206 & exp_207;
  assign exp_206 = exp_214;
  assign exp_214 = exp_5 & exp_213;
  assign exp_207 = exp_6;
  assign stdin_ready_out = exp_245;
  assign stdout_valid_out = exp_200;
  assign stdout_out = exp_181;
  assign leds_out = exp_221;

endmodule