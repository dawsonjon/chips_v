
module soc(clk, stdin_valid_in, stdin_in, stdout_ready_in, stdin_ready_out, stdout_valid_out, stdout_out, leds_out);
  input [0:0] stdin_valid_in;
  input [31:0] stdin_in;
  input [0:0] stdout_ready_in;
  input [0:0] clk;
  output [0:0] stdin_ready_out;
  output [0:0] stdout_valid_out;
  output [31:0] stdout_out;
  output [31:0] leds_out;
  wire [0:0] exp_245;
  wire [0:0] exp_228;
  wire [0:0] exp_236;
  wire [0:0] exp_5;
  wire [0:0] exp_250;
  wire [0:0] exp_597;
  wire [0:0] exp_534;
  wire [0:0] exp_399;
  wire [6:0] exp_384;
  wire [31:0] exp_382;
  wire [31:0] exp_96;
  wire [31:0] exp_95;
  wire [23:0] exp_94;
  wire [15:0] exp_93;
  wire [7:0] exp_82;
  wire [0:0] exp_81;
  wire [0:0] exp_86;
  wire [11:0] exp_77;
  wire [29:0] exp_85;
  wire [31:0] exp_8;
  wire [31:0] exp_264;
  wire [32:0] exp_867;
  wire [0:0] exp_863;
  wire [0:0] exp_559;
  wire [0:0] exp_537;
  wire [0:0] exp_395;
  wire [6:0] exp_394;
  wire [0:0] exp_397;
  wire [6:0] exp_396;
  wire [0:0] exp_558;
  wire [0:0] exp_403;
  wire [6:0] exp_402;
  wire [0:0] exp_557;
  wire [0:0] exp_556;
  wire [0:0] exp_555;
  wire [2:0] exp_385;
  wire [0:0] exp_554;
  wire [0:0] exp_538;
  wire [31:0] exp_374;
  wire [31:0] exp_312;
  wire [0:0] exp_308;
  wire [4:0] exp_288;
  wire [0:0] exp_307;
  wire [0:0] exp_311;
  wire [31:0] exp_304;
  wire [0:0] exp_285;
  wire [0:0] exp_858;
  wire [0:0] exp_857;
  wire [0:0] exp_856;
  wire [0:0] exp_855;
  wire [4:0] exp_267;
  wire [4:0] exp_850;
  wire [0:0] exp_849;
  wire [0:0] exp_441;
  wire [0:0] exp_440;
  wire [0:0] exp_439;
  wire [0:0] exp_438;
  wire [0:0] exp_437;
  wire [0:0] exp_436;
  wire [0:0] exp_387;
  wire [4:0] exp_386;
  wire [0:0] exp_389;
  wire [5:0] exp_388;
  wire [0:0] exp_391;
  wire [5:0] exp_390;
  wire [0:0] exp_393;
  wire [4:0] exp_392;
  wire [0:0] exp_844;
  wire [0:0] exp_843;
  wire [0:0] exp_629;
  wire [0:0] exp_603;
  wire [0:0] exp_601;
  wire [6:0] exp_599;
  wire [5:0] exp_600;
  wire [0:0] exp_602;
  wire [0:0] exp_628;
  wire [2:0] exp_598;
  wire [0:0] exp_842;
  wire [0:0] exp_840;
  wire [0:0] exp_833;
  wire [2:0] exp_748;
  wire [2:0] exp_755;
  wire [0:0] exp_750;
  wire [2:0] exp_749;
  wire [0:0] exp_754;
  wire [2:0] exp_752;
  wire [0:0] exp_751;
  wire [0:0] exp_753;
  wire [0:0] exp_744;
  wire [0:0] exp_743;
  wire [0:0] exp_742;
  wire [2:0] exp_832;
  wire [0:0] exp_841;
  wire [0:0] exp_651;
  wire [5:0] exp_635;
  wire [5:0] exp_642;
  wire [0:0] exp_637;
  wire [5:0] exp_636;
  wire [0:0] exp_641;
  wire [5:0] exp_639;
  wire [0:0] exp_638;
  wire [0:0] exp_640;
  wire [5:0] exp_650;
  wire [0:0] exp_262;
  wire [0:0] exp_261;
  wire [0:0] exp_259;
  wire [0:0] exp_258;
  wire [0:0] exp_256;
  wire [0:0] exp_257;
  wire [0:0] exp_255;
  wire [0:0] exp_868;
  wire [0:0] exp_254;
  wire [0:0] exp_253;
  wire [0:0] exp_872;
  wire [0:0] exp_871;
  wire [0:0] exp_870;
  wire [0:0] exp_869;
  wire [0:0] exp_249;
  wire [0:0] exp_240;
  wire [0:0] exp_235;
  wire [0:0] exp_232;
  wire [31:0] exp_1;
  wire [31:0] exp_246;
  wire [31:0] exp_453;
  wire [31:0] exp_452;
  wire [31:0] exp_451;
  wire [31:0] exp_450;
  wire [11:0] exp_449;
  wire [11:0] exp_448;
  wire [11:0] exp_447;
  wire [0:0] exp_401;
  wire [5:0] exp_400;
  wire [0:0] exp_446;
  wire [11:0] exp_442;
  wire [11:0] exp_445;
  wire [6:0] exp_443;
  wire [4:0] exp_444;
  wire [31:0] exp_231;
  wire [0:0] exp_234;
  wire [31:0] exp_233;
  wire [0:0] exp_239;
  wire [0:0] exp_218;
  wire [0:0] exp_213;
  wire [0:0] exp_210;
  wire [31:0] exp_209;
  wire [0:0] exp_212;
  wire [31:0] exp_211;
  wire [0:0] exp_217;
  wire [0:0] exp_196;
  wire [0:0] exp_191;
  wire [0:0] exp_188;
  wire [31:0] exp_187;
  wire [0:0] exp_190;
  wire [31:0] exp_189;
  wire [0:0] exp_195;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_147;
  wire [31:0] exp_146;
  wire [0:0] exp_149;
  wire [31:0] exp_148;
  wire [0:0] exp_154;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_18;
  wire [0:0] exp_17;
  wire [0:0] exp_20;
  wire [13:0] exp_19;
  wire [0:0] exp_25;
  wire [0:0] exp_4;
  wire [0:0] exp_13;
  wire [0:0] exp_138;
  wire [0:0] exp_15;
  wire [0:0] exp_6;
  wire [0:0] exp_251;
  wire [0:0] exp_536;
  wire [0:0] exp_535;
  wire [0:0] exp_137;
  wire [0:0] exp_132;
  wire [0:0] exp_136;
  wire [0:0] exp_134;
  wire [0:0] exp_14;
  wire [0:0] exp_22;
  wire [0:0] exp_133;
  wire [0:0] exp_135;
  wire [0:0] exp_131;
  wire [0:0] exp_117;
  wire [0:0] exp_142;
  wire [0:0] exp_176;
  wire [0:0] exp_183;
  wire [0:0] exp_198;
  wire [0:0] exp_205;
  wire [0:0] exp_223;
  wire [0:0] exp_227;
  wire [0:0] exp_243;
  wire [0:0] exp_846;
  wire [0:0] exp_845;
  wire [0:0] exp_260;
  wire [0:0] exp_303;
  wire [31:0] exp_275;
  wire [0:0] exp_274;
  wire [1:0] exp_283;
  wire [4:0] exp_270;
  wire [0:0] exp_273;
  wire [0:0] exp_852;
  wire [0:0] exp_851;
  wire [4:0] exp_269;
  wire [31:0] exp_271;
  wire [31:0] exp_848;
  wire [0:0] exp_847;
  wire [31:0] exp_484;
  wire [0:0] exp_483;
  wire [31:0] exp_435;
  wire [2:0] exp_378;
  wire [2:0] exp_369;
  wire [0:0] exp_366;
  wire [0:0] exp_300;
  wire [6:0] exp_290;
  wire [6:0] exp_299;
  wire [0:0] exp_302;
  wire [6:0] exp_301;
  wire [0:0] exp_368;
  wire [2:0] exp_356;
  wire [0:0] exp_298;
  wire [4:0] exp_297;
  wire [0:0] exp_355;
  wire [2:0] exp_343;
  wire [0:0] exp_296;
  wire [5:0] exp_295;
  wire [0:0] exp_342;
  wire [2:0] exp_292;
  wire [0:0] exp_341;
  wire [0:0] exp_354;
  wire [0:0] exp_367;
  wire [0:0] exp_373;
  wire [0:0] exp_434;
  wire [31:0] exp_414;
  wire [0:0] exp_380;
  wire [0:0] exp_372;
  wire [0:0] exp_358;
  wire [0:0] exp_345;
  wire [0:0] exp_331;
  wire [0:0] exp_329;
  wire [0:0] exp_330;
  wire [0:0] exp_294;
  wire [4:0] exp_293;
  wire [0:0] exp_344;
  wire [0:0] exp_357;
  wire [0:0] exp_371;
  wire [0:0] exp_370;
  wire [0:0] exp_413;
  wire [31:0] exp_411;
  wire [31:0] exp_376;
  wire [31:0] exp_362;
  wire [0:0] exp_359;
  wire [0:0] exp_361;
  wire [31:0] exp_351;
  wire [0:0] exp_350;
  wire [31:0] exp_337;
  wire [0:0] exp_336;
  wire [31:0] exp_335;
  wire [31:0] exp_333;
  wire [19:0] exp_332;
  wire [3:0] exp_334;
  wire [31:0] exp_349;
  wire [31:0] exp_347;
  wire [19:0] exp_346;
  wire [3:0] exp_348;
  wire [31:0] exp_360;
  wire [31:0] exp_377;
  wire [31:0] exp_365;
  wire [0:0] exp_363;
  wire [0:0] exp_364;
  wire [31:0] exp_353;
  wire [0:0] exp_352;
  wire [31:0] exp_340;
  wire [0:0] exp_339;
  wire [31:0] exp_324;
  wire [0:0] exp_323;
  wire [31:0] exp_318;
  wire [0:0] exp_314;
  wire [4:0] exp_289;
  wire [0:0] exp_313;
  wire [0:0] exp_317;
  wire [31:0] exp_306;
  wire [0:0] exp_286;
  wire [0:0] exp_862;
  wire [0:0] exp_861;
  wire [0:0] exp_860;
  wire [0:0] exp_859;
  wire [4:0] exp_268;
  wire [0:0] exp_305;
  wire [31:0] exp_282;
  wire [0:0] exp_281;
  wire [1:0] exp_284;
  wire [4:0] exp_277;
  wire [0:0] exp_280;
  wire [0:0] exp_854;
  wire [0:0] exp_853;
  wire [4:0] exp_276;
  wire [31:0] exp_278;
  wire [31:0] exp_287;
  wire [31:0] exp_316;
  wire [0:0] exp_315;
  wire [31:0] exp_322;
  wire [31:0] exp_319;
  wire [31:0] exp_321;
  wire [11:0] exp_320;
  wire [31:0] exp_338;
  wire [31:0] exp_266;
  wire [0:0] exp_265;
  wire [31:0] exp_412;
  wire [31:0] exp_416;
  wire [31:0] exp_415;
  wire [5:0] exp_410;
  wire [5:0] exp_409;
  wire [5:0] exp_408;
  wire [4:0] exp_379;
  wire [4:0] exp_328;
  wire [0:0] exp_327;
  wire [4:0] exp_326;
  wire [4:0] exp_291;
  wire [31:0] exp_432;
  wire [1:0] exp_418;
  wire [0:0] exp_417;
  wire [31:0] exp_433;
  wire [1:0] exp_424;
  wire [0:0] exp_423;
  wire [31:0] exp_420;
  wire [31:0] exp_419;
  wire [31:0] exp_422;
  wire [31:0] exp_421;
  wire [31:0] exp_425;
  wire [31:0] exp_429;
  wire [32:0] exp_428;
  wire [32:0] exp_426;
  wire [0:0] exp_407;
  wire [0:0] exp_381;
  wire [0:0] exp_325;
  wire [0:0] exp_406;
  wire [0:0] exp_405;
  wire [0:0] exp_404;
  wire [32:0] exp_427;
  wire [31:0] exp_430;
  wire [31:0] exp_431;
  wire [31:0] exp_482;
  wire [0:0] exp_481;
  wire [31:0] exp_472;
  wire [7:0] exp_471;
  wire [7:0] exp_470;
  wire [7:0] exp_465;
  wire [1:0] exp_456;
  wire [1:0] exp_455;
  wire [1:0] exp_454;
  wire [0:0] exp_464;
  wire [7:0] exp_460;
  wire [31:0] exp_248;
  wire [31:0] exp_238;
  wire [0:0] exp_237;
  wire [31:0] exp_216;
  wire [0:0] exp_215;
  wire [31:0] exp_194;
  wire [0:0] exp_193;
  wire [31:0] exp_153;
  wire [0:0] exp_152;
  wire [31:0] exp_24;
  wire [0:0] exp_23;
  wire [31:0] exp_3;
  wire [31:0] exp_12;
  wire [31:0] exp_119;
  wire [31:0] exp_130;
  wire [23:0] exp_129;
  wire [15:0] exp_128;
  wire [7:0] exp_54;
  wire [0:0] exp_53;
  wire [0:0] exp_121;
  wire [11:0] exp_49;
  wire [29:0] exp_120;
  wire [31:0] exp_10;
  wire [0:0] exp_52;
  wire [0:0] exp_116;
  wire [0:0] exp_114;
  wire [0:0] exp_115;
  wire [3:0] exp_16;
  wire [3:0] exp_7;
  wire [3:0] exp_252;
  wire [3:0] exp_533;
  wire [0:0] exp_532;
  wire [3:0] exp_520;
  wire [3:0] exp_516;
  wire [1:0] exp_519;
  wire [1:0] exp_518;
  wire [1:0] exp_517;
  wire [3:0] exp_525;
  wire [3:0] exp_521;
  wire [0:0] exp_524;
  wire [0:0] exp_523;
  wire [0:0] exp_522;
  wire [3:0] exp_526;
  wire [3:0] exp_527;
  wire [3:0] exp_528;
  wire [3:0] exp_529;
  wire [3:0] exp_530;
  wire [3:0] exp_531;
  wire [11:0] exp_48;
  wire [29:0] exp_112;
  wire [7:0] exp_50;
  wire [7:0] exp_113;
  wire [31:0] exp_11;
  wire [31:0] exp_2;
  wire [31:0] exp_247;
  wire [31:0] exp_515;
  wire [0:0] exp_514;
  wire [31:0] exp_502;
  wire [0:0] exp_501;
  wire [31:0] exp_488;
  wire [7:0] exp_487;
  wire [7:0] exp_486;
  wire [7:0] exp_485;
  wire [31:0] exp_375;
  wire [31:0] exp_496;
  wire [3:0] exp_495;
  wire [31:0] exp_498;
  wire [4:0] exp_497;
  wire [31:0] exp_500;
  wire [4:0] exp_499;
  wire [31:0] exp_506;
  wire [0:0] exp_459;
  wire [0:0] exp_458;
  wire [0:0] exp_457;
  wire [0:0] exp_505;
  wire [31:0] exp_492;
  wire [15:0] exp_491;
  wire [15:0] exp_490;
  wire [15:0] exp_489;
  wire [31:0] exp_504;
  wire [4:0] exp_503;
  wire [31:0] exp_508;
  wire [31:0] exp_507;
  wire [31:0] exp_494;
  wire [31:0] exp_493;
  wire [31:0] exp_509;
  wire [31:0] exp_510;
  wire [31:0] exp_511;
  wire [31:0] exp_512;
  wire [31:0] exp_513;
  wire [7:0] exp_47;
  wire [7:0] exp_75;
  wire [0:0] exp_74;
  wire [0:0] exp_88;
  wire [11:0] exp_70;
  wire [29:0] exp_87;
  wire [0:0] exp_73;
  wire [0:0] exp_84;
  wire [11:0] exp_69;
  wire [31:0] exp_83;
  wire [7:0] exp_71;
  wire [0:0] exp_46;
  wire [0:0] exp_123;
  wire [11:0] exp_42;
  wire [29:0] exp_122;
  wire [0:0] exp_45;
  wire [0:0] exp_111;
  wire [0:0] exp_109;
  wire [0:0] exp_110;
  wire [11:0] exp_41;
  wire [29:0] exp_107;
  wire [7:0] exp_43;
  wire [7:0] exp_108;
  wire [7:0] exp_40;
  wire [7:0] exp_68;
  wire [0:0] exp_67;
  wire [0:0] exp_90;
  wire [11:0] exp_63;
  wire [29:0] exp_89;
  wire [0:0] exp_66;
  wire [11:0] exp_62;
  wire [7:0] exp_64;
  wire [0:0] exp_39;
  wire [0:0] exp_125;
  wire [11:0] exp_35;
  wire [29:0] exp_124;
  wire [0:0] exp_38;
  wire [0:0] exp_106;
  wire [0:0] exp_104;
  wire [0:0] exp_105;
  wire [11:0] exp_34;
  wire [29:0] exp_102;
  wire [7:0] exp_36;
  wire [7:0] exp_103;
  wire [7:0] exp_33;
  wire [7:0] exp_61;
  wire [0:0] exp_60;
  wire [0:0] exp_92;
  wire [11:0] exp_56;
  wire [29:0] exp_91;
  wire [0:0] exp_59;
  wire [11:0] exp_55;
  wire [7:0] exp_57;
  wire [0:0] exp_32;
  wire [0:0] exp_127;
  wire [11:0] exp_28;
  wire [29:0] exp_126;
  wire [0:0] exp_31;
  wire [0:0] exp_101;
  wire [0:0] exp_99;
  wire [0:0] exp_100;
  wire [11:0] exp_27;
  wire [29:0] exp_97;
  wire [7:0] exp_29;
  wire [7:0] exp_98;
  wire [0:0] exp_118;
  wire [31:0] exp_141;
  wire [31:0] exp_179;
  wire [0:0] exp_177;
  wire [31:0] exp_139;
  wire [0:0] exp_178;
  wire [31:0] exp_157;
  wire [31:0] exp_164;
  wire [0:0] exp_159;
  wire [31:0] exp_158;
  wire [0:0] exp_163;
  wire [31:0] exp_161;
  wire [0:0] exp_160;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [31:0] exp_167;
  wire [31:0] exp_174;
  wire [0:0] exp_169;
  wire [31:0] exp_168;
  wire [0:0] exp_173;
  wire [31:0] exp_171;
  wire [0:0] exp_170;
  wire [0:0] exp_172;
  wire [0:0] exp_166;
  wire [0:0] exp_165;
  wire [31:0] exp_182;
  wire [31:0] exp_201;
  wire [31:0] exp_204;
  wire [31:0] exp_222;
  wire [31:0] exp_226;
  wire [31:0] exp_241;
  wire [7:0] exp_461;
  wire [7:0] exp_462;
  wire [7:0] exp_463;
  wire [31:0] exp_475;
  wire [15:0] exp_474;
  wire [15:0] exp_473;
  wire [15:0] exp_469;
  wire [0:0] exp_468;
  wire [15:0] exp_466;
  wire [15:0] exp_467;
  wire [31:0] exp_476;
  wire [31:0] exp_477;
  wire [31:0] exp_478;
  wire [31:0] exp_479;
  wire [31:0] exp_480;
  wire [31:0] exp_839;
  wire [0:0] exp_838;
  wire [31:0] exp_835;
  wire [0:0] exp_606;
  wire [0:0] exp_605;
  wire [0:0] exp_604;
  wire [0:0] exp_834;
  wire [31:0] exp_830;
  wire [63:0] exp_829;
  wire [0:0] exp_826;
  wire [0:0] exp_809;
  wire [0:0] exp_786;
  wire [0:0] exp_783;
  wire [0:0] exp_781;
  wire [0:0] exp_763;
  wire [0:0] exp_762;
  wire [0:0] exp_761;
  wire [31:0] exp_759;
  wire [0:0] exp_758;
  wire [0:0] exp_757;
  wire [0:0] exp_746;
  wire [0:0] exp_745;
  wire [0:0] exp_609;
  wire [0:0] exp_608;
  wire [0:0] exp_607;
  wire [0:0] exp_612;
  wire [0:0] exp_611;
  wire [1:0] exp_610;
  wire [0:0] exp_782;
  wire [0:0] exp_766;
  wire [0:0] exp_765;
  wire [0:0] exp_764;
  wire [31:0] exp_760;
  wire [0:0] exp_747;
  wire [0:0] exp_768;
  wire [0:0] exp_767;
  wire [0:0] exp_788;
  wire [1:0] exp_787;
  wire [0:0] exp_811;
  wire [1:0] exp_810;
  wire [0:0] exp_828;
  wire [63:0] exp_825;
  wire [63:0] exp_824;
  wire [63:0] exp_820;
  wire [63:0] exp_816;
  wire [63:0] exp_812;
  wire [31:0] exp_805;
  wire [31:0] exp_792;
  wire [31:0] exp_790;
  wire [15:0] exp_789;
  wire [31:0] exp_784;
  wire [31:0] exp_774;
  wire [31:0] exp_773;
  wire [31:0] exp_772;
  wire [0:0] exp_769;
  wire [0:0] exp_771;
  wire [31:0] exp_770;
  wire [15:0] exp_791;
  wire [31:0] exp_785;
  wire [31:0] exp_780;
  wire [31:0] exp_779;
  wire [31:0] exp_778;
  wire [0:0] exp_775;
  wire [0:0] exp_777;
  wire [31:0] exp_776;
  wire [63:0] exp_815;
  wire [63:0] exp_813;
  wire [31:0] exp_806;
  wire [31:0] exp_796;
  wire [31:0] exp_794;
  wire [15:0] exp_793;
  wire [15:0] exp_795;
  wire [4:0] exp_814;
  wire [63:0] exp_819;
  wire [63:0] exp_817;
  wire [31:0] exp_807;
  wire [31:0] exp_800;
  wire [31:0] exp_798;
  wire [15:0] exp_797;
  wire [15:0] exp_799;
  wire [4:0] exp_818;
  wire [63:0] exp_823;
  wire [63:0] exp_821;
  wire [31:0] exp_808;
  wire [31:0] exp_804;
  wire [31:0] exp_802;
  wire [15:0] exp_801;
  wire [15:0] exp_803;
  wire [5:0] exp_822;
  wire [63:0] exp_827;
  wire [31:0] exp_831;
  wire [31:0] exp_837;
  wire [0:0] exp_630;
  wire [0:0] exp_836;
  wire [31:0] exp_740;
  wire [31:0] exp_734;
  wire [0:0] exp_730;
  wire [0:0] exp_729;
  wire [31:0] exp_678;
  wire [31:0] exp_675;
  wire [31:0] exp_674;
  wire [31:0] exp_673;
  wire [0:0] exp_670;
  wire [0:0] exp_661;
  wire [0:0] exp_660;
  wire [0:0] exp_659;
  wire [31:0] exp_655;
  wire [0:0] exp_653;
  wire [0:0] exp_652;
  wire [0:0] exp_632;
  wire [0:0] exp_631;
  wire [0:0] exp_672;
  wire [31:0] exp_671;
  wire [0:0] exp_663;
  wire [0:0] exp_662;
  wire [0:0] exp_728;
  wire [0:0] exp_733;
  wire [31:0] exp_721;
  wire [31:0] exp_720;
  wire [31:0] exp_719;
  wire [0:0] exp_716;
  wire [0:0] exp_680;
  wire [0:0] exp_676;
  wire [0:0] exp_658;
  wire [0:0] exp_657;
  wire [0:0] exp_656;
  wire [31:0] exp_654;
  wire [0:0] exp_718;
  wire [31:0] exp_714;
  wire [31:0] exp_684;
  wire [31:0] exp_711;
  wire [0:0] exp_645;
  wire [1:0] exp_644;
  wire [0:0] exp_710;
  wire [31:0] exp_703;
  wire [0:0] exp_693;
  wire [0:0] exp_692;
  wire [32:0] exp_691;
  wire [32:0] exp_690;
  wire [32:0] exp_689;
  wire [31:0] exp_687;
  wire [31:0] exp_682;
  wire [32:0] exp_708;
  wire [0:0] exp_707;
  wire [32:0] exp_695;
  wire [0:0] exp_694;
  wire [0:0] exp_706;
  wire [0:0] exp_681;
  wire [0:0] exp_688;
  wire [31:0] exp_686;
  wire [31:0] exp_713;
  wire [0:0] exp_712;
  wire [31:0] exp_705;
  wire [0:0] exp_704;
  wire [31:0] exp_677;
  wire [31:0] exp_669;
  wire [31:0] exp_668;
  wire [31:0] exp_667;
  wire [0:0] exp_664;
  wire [0:0] exp_666;
  wire [31:0] exp_665;
  wire [0:0] exp_685;
  wire [0:0] exp_702;
  wire [31:0] exp_697;
  wire [0:0] exp_696;
  wire [31:0] exp_701;
  wire [31:0] exp_699;
  wire [0:0] exp_698;
  wire [0:0] exp_700;
  wire [0:0] exp_709;
  wire [0:0] exp_683;
  wire [0:0] exp_647;
  wire [5:0] exp_646;
  wire [31:0] exp_717;
  wire [31:0] exp_732;
  wire [0:0] exp_731;
  wire [0:0] exp_649;
  wire [5:0] exp_648;
  wire [31:0] exp_741;
  wire [31:0] exp_739;
  wire [0:0] exp_737;
  wire [0:0] exp_736;
  wire [0:0] exp_735;
  wire [0:0] exp_738;
  wire [31:0] exp_727;
  wire [31:0] exp_726;
  wire [31:0] exp_725;
  wire [0:0] exp_722;
  wire [0:0] exp_679;
  wire [0:0] exp_724;
  wire [31:0] exp_715;
  wire [31:0] exp_723;
  wire [31:0] exp_310;
  wire [0:0] exp_309;
  wire [0:0] exp_539;
  wire [0:0] exp_552;
  wire [0:0] exp_553;
  wire [0:0] exp_540;
  wire [0:0] exp_541;
  wire [0:0] exp_546;
  wire [31:0] exp_543;
  wire [31:0] exp_542;
  wire [31:0] exp_545;
  wire [31:0] exp_544;
  wire [0:0] exp_551;
  wire [31:0] exp_548;
  wire [31:0] exp_547;
  wire [31:0] exp_550;
  wire [31:0] exp_549;
  wire [0:0] exp_866;
  wire [31:0] exp_865;
  wire [2:0] exp_864;
  wire [32:0] exp_596;
  wire [0:0] exp_595;
  wire [31:0] exp_586;
  wire [31:0] exp_585;
  wire [0:0] exp_584;
  wire [31:0] exp_571;
  wire [12:0] exp_570;
  wire [12:0] exp_569;
  wire [12:0] exp_568;
  wire [11:0] exp_567;
  wire [7:0] exp_566;
  wire [1:0] exp_565;
  wire [0:0] exp_560;
  wire [0:0] exp_561;
  wire [5:0] exp_562;
  wire [3:0] exp_563;
  wire [0:0] exp_564;
  wire [31:0] exp_583;
  wire [20:0] exp_582;
  wire [20:0] exp_581;
  wire [20:0] exp_580;
  wire [19:0] exp_579;
  wire [9:0] exp_578;
  wire [8:0] exp_577;
  wire [0:0] exp_572;
  wire [7:0] exp_573;
  wire [0:0] exp_574;
  wire [9:0] exp_575;
  wire [0:0] exp_576;
  wire [31:0] exp_383;
  wire [32:0] exp_594;
  wire [32:0] exp_593;
  wire [31:0] exp_591;
  wire [31:0] exp_590;
  wire [11:0] exp_589;
  wire [11:0] exp_588;
  wire [11:0] exp_587;
  wire [32:0] exp_592;
  wire [0:0] exp_263;
  wire [0:0] exp_80;
  wire [11:0] exp_76;
  wire [7:0] exp_78;
  wire [0:0] exp_9;
  wire [1:0] exp_398;
  wire [0:0] exp_244;
  wire [0:0] exp_229;
  wire [0:0] exp_200;
  wire [0:0] exp_184;
  wire [0:0] exp_192;
  wire [0:0] exp_185;
  wire [31:0] exp_181;
  wire [31:0] exp_221;
  wire [31:0] exp_203;
  wire [0:0] exp_220;
  wire [0:0] exp_206;
  wire [0:0] exp_214;
  wire [0:0] exp_207;

  assign exp_245 = exp_228 & exp_244;
  assign exp_228 = exp_236;
  assign exp_236 = exp_5 & exp_235;
  assign exp_5 = exp_250;
  assign exp_250 = exp_597;
  assign exp_597 = exp_534 & exp_262;
  assign exp_534 = exp_399 | exp_401;
  assign exp_399 = exp_384 == exp_398;
  assign exp_384 = exp_382[6:0];

      reg [31:0] exp_382_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_382_reg <= exp_96;
        end
      end
      assign exp_382 = exp_382_reg;
    
      reg [31:0] exp_96_reg = 0;
      always@(posedge clk) begin
        if (exp_9) begin
          exp_96_reg <= exp_95;
        end
      end
      assign exp_96 = exp_96_reg;
      assign exp_95 = {exp_94, exp_61};  assign exp_94 = {exp_93, exp_68};  assign exp_93 = {exp_82, exp_75};  assign exp_81 = exp_86;
  assign exp_86 = 1;
  assign exp_77 = exp_85;
  assign exp_85 = exp_8[31:2];
  assign exp_8 = exp_264;

      reg [31:0] exp_264_reg = 0;
      always@(posedge clk) begin
        if (exp_263) begin
          exp_264_reg <= exp_867;
        end
      end
      assign exp_264 = exp_264_reg;
    
  reg [32:0] exp_867_reg;
  always@(*) begin
    case (exp_863)
      0:exp_867_reg <= exp_865;
      1:exp_867_reg <= exp_596;
      default:exp_867_reg <= exp_866;
    endcase
  end
  assign exp_867 = exp_867_reg;
  assign exp_863 = exp_559 & exp_262;
  assign exp_559 = exp_537 | exp_558;
  assign exp_537 = exp_395 | exp_397;
  assign exp_395 = exp_384 == exp_394;
  assign exp_394 = 111;
  assign exp_397 = exp_384 == exp_396;
  assign exp_396 = 103;

  reg [0:0] exp_558_reg;
  always@(*) begin
    case (exp_403)
      0:exp_558_reg <= exp_556;
      1:exp_558_reg <= exp_555;
      default:exp_558_reg <= exp_557;
    endcase
  end
  assign exp_558 = exp_558_reg;
  assign exp_403 = exp_384 == exp_402;
  assign exp_402 = 99;
  assign exp_557 = 0;
  assign exp_556 = 0;

  reg [0:0] exp_555_reg;
  always@(*) begin
    case (exp_385)
      0:exp_555_reg <= exp_538;
      1:exp_555_reg <= exp_539;
      2:exp_555_reg <= exp_552;
      3:exp_555_reg <= exp_553;
      4:exp_555_reg <= exp_540;
      5:exp_555_reg <= exp_541;
      6:exp_555_reg <= exp_546;
      7:exp_555_reg <= exp_551;
      default:exp_555_reg <= exp_554;
    endcase
  end
  assign exp_555 = exp_555_reg;
  assign exp_385 = exp_382[14:12];
  assign exp_554 = 0;
  assign exp_538 = exp_374 == exp_375;

      reg [31:0] exp_374_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_374_reg <= exp_312;
        end
      end
      assign exp_374 = exp_374_reg;
    
  reg [31:0] exp_312_reg;
  always@(*) begin
    case (exp_308)
      0:exp_312_reg <= exp_304;
      1:exp_312_reg <= exp_310;
      default:exp_312_reg <= exp_311;
    endcase
  end
  assign exp_312 = exp_312_reg;
  assign exp_308 = exp_288 == exp_307;
  assign exp_288 = exp_96[19:15];
  assign exp_307 = 0;
  assign exp_311 = 0;

  reg [31:0] exp_304_reg;
  always@(*) begin
    case (exp_285)
      0:exp_304_reg <= exp_275;
      1:exp_304_reg <= exp_287;
      default:exp_304_reg <= exp_303;
    endcase
  end
  assign exp_304 = exp_304_reg;
  assign exp_285 = exp_858;
  assign exp_858 = exp_857 & exp_254;
  assign exp_857 = exp_856 & exp_262;
  assign exp_856 = exp_855 & exp_849;
  assign exp_855 = exp_267 == exp_850;
  assign exp_267 = exp_96[19:15];
  assign exp_850 = exp_382[11:7];
  assign exp_849 = exp_441 | exp_844;
  assign exp_441 = exp_440 | exp_399;
  assign exp_440 = exp_439 | exp_393;
  assign exp_439 = exp_438 | exp_391;
  assign exp_438 = exp_437 | exp_397;
  assign exp_437 = exp_436 | exp_395;
  assign exp_436 = exp_387 | exp_389;
  assign exp_387 = exp_384 == exp_386;
  assign exp_386 = 19;
  assign exp_389 = exp_384 == exp_388;
  assign exp_388 = 51;
  assign exp_391 = exp_384 == exp_390;
  assign exp_390 = 55;
  assign exp_393 = exp_384 == exp_392;
  assign exp_392 = 23;
  assign exp_844 = exp_843 & exp_603;

  reg [0:0] exp_843_reg;
  always@(*) begin
    case (exp_629)
      0:exp_843_reg <= exp_840;
      1:exp_843_reg <= exp_841;
      default:exp_843_reg <= exp_842;
    endcase
  end
  assign exp_843 = exp_843_reg;
  assign exp_629 = exp_603 & exp_628;
  assign exp_603 = exp_601 & exp_602;
  assign exp_601 = exp_599 == exp_600;
  assign exp_599 = exp_382[6:0];
  assign exp_600 = 51;
  assign exp_602 = exp_382[25:25];
  assign exp_628 = exp_598[2:2];
  assign exp_598 = exp_382[14:12];
  assign exp_842 = 0;
  assign exp_840 = exp_833 & exp_603;
  assign exp_833 = exp_748 == exp_832;

      reg [2:0] exp_748_reg = 0;
      always@(posedge clk) begin
        if (exp_744) begin
          exp_748_reg <= exp_755;
        end
      end
      assign exp_748 = exp_748_reg;
    
  reg [2:0] exp_755_reg;
  always@(*) begin
    case (exp_750)
      0:exp_755_reg <= exp_752;
      1:exp_755_reg <= exp_753;
      default:exp_755_reg <= exp_754;
    endcase
  end
  assign exp_755 = exp_755_reg;
  assign exp_750 = exp_748 == exp_749;
  assign exp_749 = 4;
  assign exp_754 = 0;
  assign exp_752 = exp_748 + exp_751;
  assign exp_751 = 1;
  assign exp_753 = 0;
  assign exp_744 = exp_603 & exp_743;
  assign exp_743 = ~exp_742;
  assign exp_742 = exp_598[2:2];
  assign exp_832 = 4;
  assign exp_841 = exp_651 & exp_603;
  assign exp_651 = exp_635 == exp_650;

      reg [5:0] exp_635_reg = 0;
      always@(posedge clk) begin
        if (exp_629) begin
          exp_635_reg <= exp_642;
        end
      end
      assign exp_635 = exp_635_reg;
    
  reg [5:0] exp_642_reg;
  always@(*) begin
    case (exp_637)
      0:exp_642_reg <= exp_639;
      1:exp_642_reg <= exp_640;
      default:exp_642_reg <= exp_641;
    endcase
  end
  assign exp_642 = exp_642_reg;
  assign exp_637 = exp_635 == exp_636;
  assign exp_636 = 37;
  assign exp_641 = 0;
  assign exp_639 = exp_635 + exp_638;
  assign exp_638 = 1;
  assign exp_640 = 0;
  assign exp_650 = 37;

      reg [0:0] exp_262_reg = 0;
      always@(posedge clk) begin
        if (exp_254) begin
          exp_262_reg <= exp_261;
        end
      end
      assign exp_262 = exp_262_reg;
      assign exp_261 = exp_259 & exp_260;

      reg [0:0] exp_259_reg = 0;
      always@(posedge clk) begin
        if (exp_254) begin
          exp_259_reg <= exp_258;
        end
      end
      assign exp_259 = exp_259_reg;
      assign exp_258 = exp_256 & exp_257;
  assign exp_256 = 1;
  assign exp_257 = ~exp_255;
  assign exp_255 = exp_868;
  assign exp_868 = exp_262 & exp_559;
  assign exp_254 = ~exp_253;
  assign exp_253 = exp_872;
  assign exp_872 = exp_262 & exp_871;
  assign exp_871 = exp_870 | exp_846;
  assign exp_870 = exp_250 & exp_869;
  assign exp_869 = ~exp_249;
  assign exp_249 = exp_240;

  reg [0:0] exp_240_reg;
  always@(*) begin
    case (exp_235)
      0:exp_240_reg <= exp_218;
      1:exp_240_reg <= exp_227;
      default:exp_240_reg <= exp_239;
    endcase
  end
  assign exp_240 = exp_240_reg;
  assign exp_235 = exp_232 & exp_234;
  assign exp_232 = exp_1 >= exp_231;
  assign exp_1 = exp_246;
  assign exp_246 = exp_453;
  assign exp_453 = exp_452 + exp_451;
  assign exp_452 = 0;
  assign exp_451 = exp_374 + exp_450;
  assign exp_450 = $signed(exp_449);
  assign exp_449 = exp_448 + exp_447;
  assign exp_448 = 0;

  reg [11:0] exp_447_reg;
  always@(*) begin
    case (exp_401)
      0:exp_447_reg <= exp_442;
      1:exp_447_reg <= exp_445;
      default:exp_447_reg <= exp_446;
    endcase
  end
  assign exp_447 = exp_447_reg;
  assign exp_401 = exp_384 == exp_400;
  assign exp_400 = 35;
  assign exp_446 = 0;
  assign exp_442 = exp_382[31:20];
  assign exp_445 = {exp_443, exp_444};  assign exp_443 = exp_382[31:25];
  assign exp_444 = exp_382[11:7];
  assign exp_231 = 2147483664;
  assign exp_234 = exp_1 <= exp_233;
  assign exp_233 = 2147483664;
  assign exp_239 = 0;

  reg [0:0] exp_218_reg;
  always@(*) begin
    case (exp_213)
      0:exp_218_reg <= exp_196;
      1:exp_218_reg <= exp_205;
      default:exp_218_reg <= exp_217;
    endcase
  end
  assign exp_218 = exp_218_reg;
  assign exp_213 = exp_210 & exp_212;
  assign exp_210 = exp_1 >= exp_209;
  assign exp_209 = 2147483660;
  assign exp_212 = exp_1 <= exp_211;
  assign exp_211 = 2147483660;
  assign exp_217 = 0;

  reg [0:0] exp_196_reg;
  always@(*) begin
    case (exp_191)
      0:exp_196_reg <= exp_155;
      1:exp_196_reg <= exp_183;
      default:exp_196_reg <= exp_195;
    endcase
  end
  assign exp_196 = exp_196_reg;
  assign exp_191 = exp_188 & exp_190;
  assign exp_188 = exp_1 >= exp_187;
  assign exp_187 = 2147483656;
  assign exp_190 = exp_1 <= exp_189;
  assign exp_189 = 2147483656;
  assign exp_195 = 0;

  reg [0:0] exp_155_reg;
  always@(*) begin
    case (exp_150)
      0:exp_155_reg <= exp_26;
      1:exp_155_reg <= exp_142;
      default:exp_155_reg <= exp_154;
    endcase
  end
  assign exp_155 = exp_155_reg;
  assign exp_150 = exp_147 & exp_149;
  assign exp_147 = exp_1 >= exp_146;
  assign exp_146 = 2147483648;
  assign exp_149 = exp_1 <= exp_148;
  assign exp_148 = 2147483652;
  assign exp_154 = 0;

  reg [0:0] exp_26_reg;
  always@(*) begin
    case (exp_21)
      0:exp_26_reg <= exp_4;
      1:exp_26_reg <= exp_13;
      default:exp_26_reg <= exp_25;
    endcase
  end
  assign exp_26 = exp_26_reg;
  assign exp_21 = exp_18 & exp_20;
  assign exp_18 = exp_1 >= exp_17;
  assign exp_17 = 0;
  assign exp_20 = exp_1 <= exp_19;
  assign exp_19 = 16380;
  assign exp_25 = 0;
  assign exp_4 = 0;
  assign exp_13 = exp_138;

  reg [0:0] exp_138_reg;
  always@(*) begin
    case (exp_15)
      0:exp_138_reg <= exp_132;
      1:exp_138_reg <= exp_117;
      default:exp_138_reg <= exp_137;
    endcase
  end
  assign exp_138 = exp_138_reg;
  assign exp_15 = exp_6;
  assign exp_6 = exp_251;
  assign exp_251 = exp_536;
  assign exp_536 = exp_535 + exp_401;
  assign exp_535 = 0;
  assign exp_137 = 0;

      reg [0:0] exp_132_reg = 0;
      always@(posedge clk) begin
        if (exp_131) begin
          exp_132_reg <= exp_136;
        end
      end
      assign exp_132 = exp_132_reg;
      assign exp_136 = exp_134 & exp_135;
  assign exp_134 = exp_14 & exp_133;
  assign exp_14 = exp_22;
  assign exp_22 = exp_5 & exp_21;
  assign exp_133 = ~exp_15;
  assign exp_135 = ~exp_132;
  assign exp_131 = 1;
  assign exp_117 = 1;
  assign exp_142 = exp_176;
  assign exp_176 = 1;
  assign exp_183 = exp_198;
  assign exp_198 = stdout_ready_in;
  assign exp_205 = exp_223;
  assign exp_223 = 1;
  assign exp_227 = exp_243;
  assign exp_243 = stdin_valid_in;
  assign exp_846 = exp_603 & exp_845;
  assign exp_845 = ~exp_843;
  assign exp_260 = ~exp_255;
  assign exp_303 = 0;

  //Create RAM
  reg [31:0] exp_275_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_273) begin
      exp_275_ram[exp_269] <= exp_271;
    end
  end
  assign exp_275 = exp_275_ram[exp_270];
  assign exp_274 = exp_283;
  assign exp_283 = 1;
  assign exp_270 = exp_267;
  assign exp_273 = exp_852;
  assign exp_852 = exp_851 & exp_254;
  assign exp_851 = exp_849 & exp_262;
  assign exp_269 = exp_850;
  assign exp_271 = exp_848;

  reg [31:0] exp_848_reg;
  always@(*) begin
    case (exp_844)
      0:exp_848_reg <= exp_484;
      1:exp_848_reg <= exp_839;
      default:exp_848_reg <= exp_847;
    endcase
  end
  assign exp_848 = exp_848_reg;
  assign exp_847 = 0;

  reg [31:0] exp_484_reg;
  always@(*) begin
    case (exp_399)
      0:exp_484_reg <= exp_435;
      1:exp_484_reg <= exp_482;
      default:exp_484_reg <= exp_483;
    endcase
  end
  assign exp_484 = exp_484_reg;
  assign exp_483 = 0;

  reg [31:0] exp_435_reg;
  always@(*) begin
    case (exp_378)
      0:exp_435_reg <= exp_414;
      1:exp_435_reg <= exp_416;
      2:exp_435_reg <= exp_432;
      3:exp_435_reg <= exp_433;
      4:exp_435_reg <= exp_425;
      5:exp_435_reg <= exp_429;
      6:exp_435_reg <= exp_430;
      7:exp_435_reg <= exp_431;
      default:exp_435_reg <= exp_434;
    endcase
  end
  assign exp_435 = exp_435_reg;

      reg [2:0] exp_378_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_378_reg <= exp_369;
        end
      end
      assign exp_378 = exp_378_reg;
    
  reg [2:0] exp_369_reg;
  always@(*) begin
    case (exp_366)
      0:exp_369_reg <= exp_356;
      1:exp_369_reg <= exp_367;
      default:exp_369_reg <= exp_368;
    endcase
  end
  assign exp_369 = exp_369_reg;
  assign exp_366 = exp_300 | exp_302;
  assign exp_300 = exp_290 == exp_299;
  assign exp_290 = exp_96[6:0];
  assign exp_299 = 111;
  assign exp_302 = exp_290 == exp_301;
  assign exp_301 = 103;
  assign exp_368 = 0;

  reg [2:0] exp_356_reg;
  always@(*) begin
    case (exp_298)
      0:exp_356_reg <= exp_343;
      1:exp_356_reg <= exp_354;
      default:exp_356_reg <= exp_355;
    endcase
  end
  assign exp_356 = exp_356_reg;
  assign exp_298 = exp_290 == exp_297;
  assign exp_297 = 23;
  assign exp_355 = 0;

  reg [2:0] exp_343_reg;
  always@(*) begin
    case (exp_296)
      0:exp_343_reg <= exp_292;
      1:exp_343_reg <= exp_341;
      default:exp_343_reg <= exp_342;
    endcase
  end
  assign exp_343 = exp_343_reg;
  assign exp_296 = exp_290 == exp_295;
  assign exp_295 = 55;
  assign exp_342 = 0;
  assign exp_292 = exp_96[14:12];
  assign exp_341 = 0;
  assign exp_354 = 0;
  assign exp_367 = 0;
  assign exp_373 = exp_254 & exp_259;
  assign exp_434 = 0;

  reg [31:0] exp_414_reg;
  always@(*) begin
    case (exp_380)
      0:exp_414_reg <= exp_411;
      1:exp_414_reg <= exp_412;
      default:exp_414_reg <= exp_413;
    endcase
  end
  assign exp_414 = exp_414_reg;

      reg [0:0] exp_380_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_380_reg <= exp_372;
        end
      end
      assign exp_380 = exp_380_reg;
      assign exp_372 = exp_358 & exp_371;
  assign exp_358 = exp_345 & exp_357;
  assign exp_345 = exp_331 & exp_344;
  assign exp_331 = exp_329 & exp_330;
  assign exp_329 = exp_96[30:30];
  assign exp_330 = ~exp_294;
  assign exp_294 = exp_290 == exp_293;
  assign exp_293 = 19;
  assign exp_344 = ~exp_296;
  assign exp_357 = ~exp_298;
  assign exp_371 = ~exp_370;
  assign exp_370 = exp_300 | exp_302;
  assign exp_413 = 0;
  assign exp_411 = exp_376 + exp_377;

      reg [31:0] exp_376_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_376_reg <= exp_362;
        end
      end
      assign exp_376 = exp_376_reg;
    
  reg [31:0] exp_362_reg;
  always@(*) begin
    case (exp_359)
      0:exp_362_reg <= exp_351;
      1:exp_362_reg <= exp_360;
      default:exp_362_reg <= exp_361;
    endcase
  end
  assign exp_362 = exp_362_reg;
  assign exp_359 = exp_300 | exp_302;
  assign exp_361 = 0;

  reg [31:0] exp_351_reg;
  always@(*) begin
    case (exp_298)
      0:exp_351_reg <= exp_337;
      1:exp_351_reg <= exp_349;
      default:exp_351_reg <= exp_350;
    endcase
  end
  assign exp_351 = exp_351_reg;
  assign exp_350 = 0;

  reg [31:0] exp_337_reg;
  always@(*) begin
    case (exp_296)
      0:exp_337_reg <= exp_312;
      1:exp_337_reg <= exp_335;
      default:exp_337_reg <= exp_336;
    endcase
  end
  assign exp_337 = exp_337_reg;
  assign exp_336 = 0;
  assign exp_335 = exp_333 << exp_334;
  assign exp_333 = exp_332;
  assign exp_332 = exp_96[31:12];
  assign exp_334 = 12;
  assign exp_349 = exp_347 << exp_348;
  assign exp_347 = exp_346;
  assign exp_346 = exp_96[31:12];
  assign exp_348 = 12;
  assign exp_360 = 4;

      reg [31:0] exp_377_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_377_reg <= exp_365;
        end
      end
      assign exp_377 = exp_377_reg;
    
  reg [31:0] exp_365_reg;
  always@(*) begin
    case (exp_363)
      0:exp_365_reg <= exp_353;
      1:exp_365_reg <= exp_266;
      default:exp_365_reg <= exp_364;
    endcase
  end
  assign exp_365 = exp_365_reg;
  assign exp_363 = exp_300 | exp_302;
  assign exp_364 = 0;

  reg [31:0] exp_353_reg;
  always@(*) begin
    case (exp_298)
      0:exp_353_reg <= exp_340;
      1:exp_353_reg <= exp_266;
      default:exp_353_reg <= exp_352;
    endcase
  end
  assign exp_353 = exp_353_reg;
  assign exp_352 = 0;

  reg [31:0] exp_340_reg;
  always@(*) begin
    case (exp_296)
      0:exp_340_reg <= exp_324;
      1:exp_340_reg <= exp_338;
      default:exp_340_reg <= exp_339;
    endcase
  end
  assign exp_340 = exp_340_reg;
  assign exp_339 = 0;

  reg [31:0] exp_324_reg;
  always@(*) begin
    case (exp_294)
      0:exp_324_reg <= exp_318;
      1:exp_324_reg <= exp_322;
      default:exp_324_reg <= exp_323;
    endcase
  end
  assign exp_324 = exp_324_reg;
  assign exp_323 = 0;

  reg [31:0] exp_318_reg;
  always@(*) begin
    case (exp_314)
      0:exp_318_reg <= exp_306;
      1:exp_318_reg <= exp_316;
      default:exp_318_reg <= exp_317;
    endcase
  end
  assign exp_318 = exp_318_reg;
  assign exp_314 = exp_289 == exp_313;
  assign exp_289 = exp_96[24:20];
  assign exp_313 = 0;
  assign exp_317 = 0;

  reg [31:0] exp_306_reg;
  always@(*) begin
    case (exp_286)
      0:exp_306_reg <= exp_282;
      1:exp_306_reg <= exp_287;
      default:exp_306_reg <= exp_305;
    endcase
  end
  assign exp_306 = exp_306_reg;
  assign exp_286 = exp_862;
  assign exp_862 = exp_861 & exp_254;
  assign exp_861 = exp_860 & exp_262;
  assign exp_860 = exp_859 & exp_849;
  assign exp_859 = exp_268 == exp_850;
  assign exp_268 = exp_96[24:20];
  assign exp_305 = 0;

  //Create RAM
  reg [31:0] exp_282_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_280) begin
      exp_282_ram[exp_276] <= exp_278;
    end
  end
  assign exp_282 = exp_282_ram[exp_277];
  assign exp_281 = exp_284;
  assign exp_284 = 1;
  assign exp_277 = exp_268;
  assign exp_280 = exp_854;
  assign exp_854 = exp_853 & exp_254;
  assign exp_853 = exp_849 & exp_262;
  assign exp_276 = exp_850;
  assign exp_278 = exp_848;
  assign exp_287 = exp_848;
  assign exp_316 = $signed(exp_315);
  assign exp_315 = 0;
  assign exp_322 = exp_319 + exp_321;
  assign exp_319 = 0;
  assign exp_321 = $signed(exp_320);
  assign exp_320 = exp_96[31:20];
  assign exp_338 = 0;

      reg [31:0] exp_266_reg = 0;
      always@(posedge clk) begin
        if (exp_265) begin
          exp_266_reg <= exp_264;
        end
      end
      assign exp_266 = exp_266_reg;
      assign exp_265 = exp_256 & exp_254;
  assign exp_412 = exp_376 - exp_377;
  assign exp_416 = exp_376 << exp_415;
  assign exp_415 = $signed(exp_410);
  assign exp_410 = exp_409 + exp_408;
  assign exp_409 = 0;
  assign exp_408 = exp_379;

      reg [4:0] exp_379_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_379_reg <= exp_328;
        end
      end
      assign exp_379 = exp_379_reg;
    
  reg [4:0] exp_328_reg;
  always@(*) begin
    case (exp_294)
      0:exp_328_reg <= exp_326;
      1:exp_328_reg <= exp_291;
      default:exp_328_reg <= exp_327;
    endcase
  end
  assign exp_328 = exp_328_reg;
  assign exp_327 = 0;
  assign exp_326 = exp_324[4:0];
  assign exp_291 = exp_96[24:20];
  assign exp_432 = $signed(exp_418);
  assign exp_418 = exp_417;
  assign exp_417 = $signed(exp_376) < $signed(exp_377);
  assign exp_433 = $signed(exp_424);
  assign exp_424 = exp_423;
  assign exp_423 = exp_420 < exp_422;
  assign exp_420 = exp_419 + exp_376;
  assign exp_419 = 0;
  assign exp_422 = exp_421 + exp_377;
  assign exp_421 = 0;
  assign exp_425 = exp_376 ^ exp_377;
  assign exp_429 = exp_428[31:0];
  assign exp_428 = $signed(exp_426) >>> $signed(exp_427);
  assign exp_426 = {exp_407, exp_376};
  reg [0:0] exp_407_reg;
  always@(*) begin
    case (exp_381)
      0:exp_407_reg <= exp_405;
      1:exp_407_reg <= exp_404;
      default:exp_407_reg <= exp_406;
    endcase
  end
  assign exp_407 = exp_407_reg;

      reg [0:0] exp_381_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_381_reg <= exp_325;
        end
      end
      assign exp_381 = exp_381_reg;
      assign exp_325 = exp_96[30:30];
  assign exp_406 = 0;
  assign exp_405 = 0;
  assign exp_404 = exp_376[31:31];
  assign exp_427 = $signed(exp_410);
  assign exp_430 = exp_376 | exp_377;
  assign exp_431 = exp_376 & exp_377;

  reg [31:0] exp_482_reg;
  always@(*) begin
    case (exp_385)
      0:exp_482_reg <= exp_472;
      1:exp_482_reg <= exp_475;
      2:exp_482_reg <= exp_248;
      3:exp_482_reg <= exp_476;
      4:exp_482_reg <= exp_477;
      5:exp_482_reg <= exp_478;
      6:exp_482_reg <= exp_479;
      7:exp_482_reg <= exp_480;
      default:exp_482_reg <= exp_481;
    endcase
  end
  assign exp_482 = exp_482_reg;
  assign exp_481 = 0;
  assign exp_472 = $signed(exp_471);
  assign exp_471 = exp_470 + exp_465;
  assign exp_470 = 0;

  reg [7:0] exp_465_reg;
  always@(*) begin
    case (exp_456)
      0:exp_465_reg <= exp_460;
      1:exp_465_reg <= exp_461;
      2:exp_465_reg <= exp_462;
      3:exp_465_reg <= exp_463;
      default:exp_465_reg <= exp_464;
    endcase
  end
  assign exp_465 = exp_465_reg;
  assign exp_456 = exp_455 + exp_454;
  assign exp_455 = 0;
  assign exp_454 = exp_453[1:0];
  assign exp_464 = 0;
  assign exp_460 = exp_248[7:0];
  assign exp_248 = exp_238;

  reg [31:0] exp_238_reg;
  always@(*) begin
    case (exp_235)
      0:exp_238_reg <= exp_216;
      1:exp_238_reg <= exp_226;
      default:exp_238_reg <= exp_237;
    endcase
  end
  assign exp_238 = exp_238_reg;
  assign exp_237 = 0;

  reg [31:0] exp_216_reg;
  always@(*) begin
    case (exp_213)
      0:exp_216_reg <= exp_194;
      1:exp_216_reg <= exp_204;
      default:exp_216_reg <= exp_215;
    endcase
  end
  assign exp_216 = exp_216_reg;
  assign exp_215 = 0;

  reg [31:0] exp_194_reg;
  always@(*) begin
    case (exp_191)
      0:exp_194_reg <= exp_153;
      1:exp_194_reg <= exp_182;
      default:exp_194_reg <= exp_193;
    endcase
  end
  assign exp_194 = exp_194_reg;
  assign exp_193 = 0;

  reg [31:0] exp_153_reg;
  always@(*) begin
    case (exp_150)
      0:exp_153_reg <= exp_24;
      1:exp_153_reg <= exp_141;
      default:exp_153_reg <= exp_152;
    endcase
  end
  assign exp_153 = exp_153_reg;
  assign exp_152 = 0;

  reg [31:0] exp_24_reg;
  always@(*) begin
    case (exp_21)
      0:exp_24_reg <= exp_3;
      1:exp_24_reg <= exp_12;
      default:exp_24_reg <= exp_23;
    endcase
  end
  assign exp_24 = exp_24_reg;
  assign exp_23 = 0;
  assign exp_3 = 0;
  assign exp_12 = exp_119;

      reg [31:0] exp_119_reg = 0;
      always@(posedge clk) begin
        if (exp_118) begin
          exp_119_reg <= exp_130;
        end
      end
      assign exp_119 = exp_119_reg;
      assign exp_130 = {exp_129, exp_33};  assign exp_129 = {exp_128, exp_40};  assign exp_128 = {exp_54, exp_47};
  //Create RAM
  reg [7:0] exp_54_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_54_ram[0] = 0;
    exp_54_ram[1] = 0;
    exp_54_ram[2] = 0;
    exp_54_ram[3] = 0;
    exp_54_ram[4] = 0;
    exp_54_ram[5] = 0;
    exp_54_ram[6] = 0;
    exp_54_ram[7] = 0;
    exp_54_ram[8] = 0;
    exp_54_ram[9] = 0;
    exp_54_ram[10] = 0;
    exp_54_ram[11] = 0;
    exp_54_ram[12] = 0;
    exp_54_ram[13] = 0;
    exp_54_ram[14] = 0;
    exp_54_ram[15] = 0;
    exp_54_ram[16] = 0;
    exp_54_ram[17] = 0;
    exp_54_ram[18] = 0;
    exp_54_ram[19] = 0;
    exp_54_ram[20] = 0;
    exp_54_ram[21] = 0;
    exp_54_ram[22] = 0;
    exp_54_ram[23] = 0;
    exp_54_ram[24] = 0;
    exp_54_ram[25] = 0;
    exp_54_ram[26] = 0;
    exp_54_ram[27] = 0;
    exp_54_ram[28] = 0;
    exp_54_ram[29] = 0;
    exp_54_ram[30] = 0;
    exp_54_ram[31] = 0;
    exp_54_ram[32] = 255;
    exp_54_ram[33] = 104;
    exp_54_ram[34] = 0;
    exp_54_ram[35] = 0;
    exp_54_ram[36] = 0;
    exp_54_ram[37] = 0;
    exp_54_ram[38] = 0;
    exp_54_ram[39] = 0;
    exp_54_ram[40] = 40;
    exp_54_ram[41] = 0;
    exp_54_ram[42] = 165;
    exp_54_ram[43] = 14;
    exp_54_ram[44] = 0;
    exp_54_ram[45] = 12;
    exp_54_ram[46] = 15;
    exp_54_ram[47] = 0;
    exp_54_ram[48] = 0;
    exp_54_ram[49] = 0;
    exp_54_ram[50] = 0;
    exp_54_ram[51] = 0;
    exp_54_ram[52] = 2;
    exp_54_ram[53] = 0;
    exp_54_ram[54] = 64;
    exp_54_ram[55] = 0;
    exp_54_ram[56] = 0;
    exp_54_ram[57] = 0;
    exp_54_ram[58] = 0;
    exp_54_ram[59] = 0;
    exp_54_ram[60] = 0;
    exp_54_ram[61] = 1;
    exp_54_ram[62] = 3;
    exp_54_ram[63] = 1;
    exp_54_ram[64] = 1;
    exp_54_ram[65] = 1;
    exp_54_ram[66] = 3;
    exp_54_ram[67] = 0;
    exp_54_ram[68] = 2;
    exp_54_ram[69] = 1;
    exp_54_ram[70] = 0;
    exp_54_ram[71] = 0;
    exp_54_ram[72] = 1;
    exp_54_ram[73] = 255;
    exp_54_ram[74] = 1;
    exp_54_ram[75] = 0;
    exp_54_ram[76] = 255;
    exp_54_ram[77] = 1;
    exp_54_ram[78] = 64;
    exp_54_ram[79] = 3;
    exp_54_ram[80] = 1;
    exp_54_ram[81] = 1;
    exp_54_ram[82] = 3;
    exp_54_ram[83] = 1;
    exp_54_ram[84] = 0;
    exp_54_ram[85] = 2;
    exp_54_ram[86] = 0;
    exp_54_ram[87] = 0;
    exp_54_ram[88] = 0;
    exp_54_ram[89] = 255;
    exp_54_ram[90] = 1;
    exp_54_ram[91] = 0;
    exp_54_ram[92] = 255;
    exp_54_ram[93] = 1;
    exp_54_ram[94] = 0;
    exp_54_ram[95] = 0;
    exp_54_ram[96] = 14;
    exp_54_ram[97] = 1;
    exp_54_ram[98] = 1;
    exp_54_ram[99] = 242;
    exp_54_ram[100] = 1;
    exp_54_ram[101] = 243;
    exp_54_ram[102] = 0;
    exp_54_ram[103] = 0;
    exp_54_ram[104] = 2;
    exp_54_ram[105] = 0;
    exp_54_ram[106] = 12;
    exp_54_ram[107] = 15;
    exp_54_ram[108] = 1;
    exp_54_ram[109] = 0;
    exp_54_ram[110] = 0;
    exp_54_ram[111] = 0;
    exp_54_ram[112] = 0;
    exp_54_ram[113] = 2;
    exp_54_ram[114] = 0;
    exp_54_ram[115] = 64;
    exp_54_ram[116] = 10;
    exp_54_ram[117] = 65;
    exp_54_ram[118] = 0;
    exp_54_ram[119] = 1;
    exp_54_ram[120] = 1;
    exp_54_ram[121] = 1;
    exp_54_ram[122] = 1;
    exp_54_ram[123] = 3;
    exp_54_ram[124] = 3;
    exp_54_ram[125] = 1;
    exp_54_ram[126] = 0;
    exp_54_ram[127] = 2;
    exp_54_ram[128] = 0;
    exp_54_ram[129] = 1;
    exp_54_ram[130] = 1;
    exp_54_ram[131] = 255;
    exp_54_ram[132] = 1;
    exp_54_ram[133] = 1;
    exp_54_ram[134] = 255;
    exp_54_ram[135] = 1;
    exp_54_ram[136] = 65;
    exp_54_ram[137] = 3;
    exp_54_ram[138] = 1;
    exp_54_ram[139] = 1;
    exp_54_ram[140] = 3;
    exp_54_ram[141] = 1;
    exp_54_ram[142] = 0;
    exp_54_ram[143] = 2;
    exp_54_ram[144] = 0;
    exp_54_ram[145] = 0;
    exp_54_ram[146] = 0;
    exp_54_ram[147] = 255;
    exp_54_ram[148] = 1;
    exp_54_ram[149] = 0;
    exp_54_ram[150] = 255;
    exp_54_ram[151] = 1;
    exp_54_ram[152] = 0;
    exp_54_ram[153] = 0;
    exp_54_ram[154] = 1;
    exp_54_ram[155] = 1;
    exp_54_ram[156] = 244;
    exp_54_ram[157] = 1;
    exp_54_ram[158] = 244;
    exp_54_ram[159] = 0;
    exp_54_ram[160] = 0;
    exp_54_ram[161] = 0;
    exp_54_ram[162] = 0;
    exp_54_ram[163] = 0;
    exp_54_ram[164] = 1;
    exp_54_ram[165] = 0;
    exp_54_ram[166] = 3;
    exp_54_ram[167] = 1;
    exp_54_ram[168] = 1;
    exp_54_ram[169] = 1;
    exp_54_ram[170] = 3;
    exp_54_ram[171] = 1;
    exp_54_ram[172] = 0;
    exp_54_ram[173] = 2;
    exp_54_ram[174] = 0;
    exp_54_ram[175] = 0;
    exp_54_ram[176] = 1;
    exp_54_ram[177] = 255;
    exp_54_ram[178] = 1;
    exp_54_ram[179] = 0;
    exp_54_ram[180] = 255;
    exp_54_ram[181] = 1;
    exp_54_ram[182] = 64;
    exp_54_ram[183] = 3;
    exp_54_ram[184] = 1;
    exp_54_ram[185] = 1;
    exp_54_ram[186] = 3;
    exp_54_ram[187] = 1;
    exp_54_ram[188] = 2;
    exp_54_ram[189] = 0;
    exp_54_ram[190] = 0;
    exp_54_ram[191] = 0;
    exp_54_ram[192] = 1;
    exp_54_ram[193] = 255;
    exp_54_ram[194] = 1;
    exp_54_ram[195] = 0;
    exp_54_ram[196] = 255;
    exp_54_ram[197] = 1;
    exp_54_ram[198] = 1;
    exp_54_ram[199] = 64;
    exp_54_ram[200] = 0;
    exp_54_ram[201] = 235;
    exp_54_ram[202] = 24;
    exp_54_ram[203] = 0;
    exp_54_ram[204] = 4;
    exp_54_ram[205] = 15;
    exp_54_ram[206] = 0;
    exp_54_ram[207] = 0;
    exp_54_ram[208] = 0;
    exp_54_ram[209] = 0;
    exp_54_ram[210] = 165;
    exp_54_ram[211] = 0;
    exp_54_ram[212] = 0;
    exp_54_ram[213] = 2;
    exp_54_ram[214] = 0;
    exp_54_ram[215] = 64;
    exp_54_ram[216] = 2;
    exp_54_ram[217] = 0;
    exp_54_ram[218] = 238;
    exp_54_ram[219] = 0;
    exp_54_ram[220] = 0;
    exp_54_ram[221] = 239;
    exp_54_ram[222] = 1;
    exp_54_ram[223] = 1;
    exp_54_ram[224] = 252;
    exp_54_ram[225] = 1;
    exp_54_ram[226] = 251;
    exp_54_ram[227] = 0;
    exp_54_ram[228] = 0;
    exp_54_ram[229] = 0;
    exp_54_ram[230] = 0;
    exp_54_ram[231] = 1;
    exp_54_ram[232] = 3;
    exp_54_ram[233] = 0;
    exp_54_ram[234] = 0;
    exp_54_ram[235] = 0;
    exp_54_ram[236] = 0;
    exp_54_ram[237] = 1;
    exp_54_ram[238] = 1;
    exp_54_ram[239] = 1;
    exp_54_ram[240] = 3;
    exp_54_ram[241] = 1;
    exp_54_ram[242] = 0;
    exp_54_ram[243] = 3;
    exp_54_ram[244] = 0;
    exp_54_ram[245] = 1;
    exp_54_ram[246] = 1;
    exp_54_ram[247] = 255;
    exp_54_ram[248] = 1;
    exp_54_ram[249] = 1;
    exp_54_ram[250] = 255;
    exp_54_ram[251] = 1;
    exp_54_ram[252] = 65;
    exp_54_ram[253] = 3;
    exp_54_ram[254] = 3;
    exp_54_ram[255] = 1;
    exp_54_ram[256] = 2;
    exp_54_ram[257] = 1;
    exp_54_ram[258] = 1;
    exp_54_ram[259] = 0;
    exp_54_ram[260] = 0;
    exp_54_ram[261] = 1;
    exp_54_ram[262] = 1;
    exp_54_ram[263] = 255;
    exp_54_ram[264] = 1;
    exp_54_ram[265] = 1;
    exp_54_ram[266] = 255;
    exp_54_ram[267] = 1;
    exp_54_ram[268] = 1;
    exp_54_ram[269] = 0;
    exp_54_ram[270] = 0;
    exp_54_ram[271] = 255;
    exp_54_ram[272] = 0;
    exp_54_ram[273] = 1;
    exp_54_ram[274] = 0;
    exp_54_ram[275] = 1;
    exp_54_ram[276] = 65;
    exp_54_ram[277] = 2;
    exp_54_ram[278] = 2;
    exp_54_ram[279] = 1;
    exp_54_ram[280] = 2;
    exp_54_ram[281] = 0;
    exp_54_ram[282] = 1;
    exp_54_ram[283] = 2;
    exp_54_ram[284] = 0;
    exp_54_ram[285] = 1;
    exp_54_ram[286] = 1;
    exp_54_ram[287] = 0;
    exp_54_ram[288] = 2;
    exp_54_ram[289] = 206;
    exp_54_ram[290] = 0;
    exp_54_ram[291] = 255;
    exp_54_ram[292] = 0;
    exp_54_ram[293] = 1;
    exp_54_ram[294] = 0;
    exp_54_ram[295] = 0;
    exp_54_ram[296] = 1;
    exp_54_ram[297] = 0;
    exp_54_ram[298] = 218;
    exp_54_ram[299] = 255;
    exp_54_ram[300] = 204;
    exp_54_ram[301] = 0;
    exp_54_ram[302] = 0;
    exp_54_ram[303] = 218;
    exp_54_ram[304] = 0;
    exp_54_ram[305] = 255;
    exp_54_ram[306] = 1;
    exp_54_ram[307] = 0;
    exp_54_ram[308] = 0;
    exp_54_ram[309] = 0;
    exp_54_ram[310] = 127;
    exp_54_ram[311] = 1;
    exp_54_ram[312] = 127;
    exp_54_ram[313] = 1;
    exp_54_ram[314] = 0;
    exp_54_ram[315] = 0;
    exp_54_ram[316] = 127;
    exp_54_ram[317] = 1;
    exp_54_ram[318] = 1;
    exp_54_ram[319] = 0;
    exp_54_ram[320] = 8;
    exp_54_ram[321] = 0;
    exp_54_ram[322] = 0;
    exp_54_ram[323] = 1;
    exp_54_ram[324] = 0;
    exp_54_ram[325] = 254;
    exp_54_ram[326] = 8;
    exp_54_ram[327] = 0;
    exp_54_ram[328] = 0;
    exp_54_ram[329] = 0;
    exp_54_ram[330] = 0;
    exp_54_ram[331] = 4;
    exp_54_ram[332] = 0;
    exp_54_ram[333] = 0;
    exp_54_ram[334] = 3;
    exp_54_ram[335] = 4;
    exp_54_ram[336] = 255;
    exp_54_ram[337] = 0;
    exp_54_ram[338] = 255;
    exp_54_ram[339] = 0;
    exp_54_ram[340] = 0;
    exp_54_ram[341] = 0;
    exp_54_ram[342] = 0;
    exp_54_ram[343] = 254;
    exp_54_ram[344] = 0;
    exp_54_ram[345] = 253;
    exp_54_ram[346] = 2;
    exp_54_ram[347] = 252;
    exp_54_ram[348] = 255;
    exp_54_ram[349] = 0;
    exp_54_ram[350] = 0;
    exp_54_ram[351] = 0;
    exp_54_ram[352] = 0;
    exp_54_ram[353] = 254;
    exp_54_ram[354] = 251;
    exp_54_ram[355] = 252;
    exp_54_ram[356] = 254;
    exp_54_ram[357] = 247;
    exp_54_ram[358] = 248;
    exp_54_ram[359] = 0;
    exp_54_ram[360] = 248;
    exp_54_ram[361] = 255;
    exp_54_ram[362] = 0;
    exp_54_ram[363] = 0;
    exp_54_ram[364] = 0;
    exp_54_ram[365] = 6;
    exp_54_ram[366] = 55;
    exp_54_ram[367] = 65;
    exp_54_ram[368] = 0;
    exp_54_ram[369] = 64;
    exp_54_ram[370] = 4;
    exp_54_ram[371] = 0;
    exp_54_ram[372] = 64;
    exp_54_ram[373] = 1;
    exp_54_ram[374] = 0;
    exp_54_ram[375] = 0;
    exp_54_ram[376] = 0;
    exp_54_ram[377] = 0;
    exp_54_ram[378] = 0;
    exp_54_ram[379] = 0;
    exp_54_ram[380] = 1;
    exp_54_ram[381] = 0;
    exp_54_ram[382] = 0;
    exp_54_ram[383] = 0;
    exp_54_ram[384] = 1;
    exp_54_ram[385] = 0;
    exp_54_ram[386] = 255;
    exp_54_ram[387] = 0;
    exp_54_ram[388] = 0;
    exp_54_ram[389] = 252;
    exp_54_ram[390] = 0;
    exp_54_ram[391] = 0;
    exp_54_ram[392] = 252;
    exp_54_ram[393] = 254;
    exp_54_ram[394] = 0;
    exp_54_ram[395] = 0;
    exp_54_ram[396] = 0;
    exp_54_ram[397] = 1;
    exp_54_ram[398] = 1;
    exp_54_ram[399] = 1;
    exp_54_ram[400] = 0;
    exp_54_ram[401] = 24;
    exp_54_ram[402] = 0;
    exp_54_ram[403] = 0;
    exp_54_ram[404] = 0;
    exp_54_ram[405] = 8;
    exp_54_ram[406] = 0;
    exp_54_ram[407] = 45;
    exp_54_ram[408] = 0;
    exp_54_ram[409] = 67;
    exp_54_ram[410] = 65;
    exp_54_ram[411] = 67;
    exp_54_ram[412] = 9;
    exp_54_ram[413] = 0;
    exp_54_ram[414] = 0;
    exp_54_ram[415] = 3;
    exp_54_ram[416] = 2;
    exp_54_ram[417] = 7;
    exp_54_ram[418] = 2;
    exp_54_ram[419] = 255;
    exp_54_ram[420] = 65;
    exp_54_ram[421] = 0;
    exp_54_ram[422] = 0;
    exp_54_ram[423] = 0;
    exp_54_ram[424] = 0;
    exp_54_ram[425] = 1;
    exp_54_ram[426] = 1;
    exp_54_ram[427] = 0;
    exp_54_ram[428] = 1;
    exp_54_ram[429] = 0;
    exp_54_ram[430] = 0;
    exp_54_ram[431] = 1;
    exp_54_ram[432] = 1;
    exp_54_ram[433] = 0;
    exp_54_ram[434] = 0;
    exp_54_ram[435] = 0;
    exp_54_ram[436] = 0;
    exp_54_ram[437] = 2;
    exp_54_ram[438] = 0;
    exp_54_ram[439] = 37;
    exp_54_ram[440] = 2;
    exp_54_ram[441] = 248;
    exp_54_ram[442] = 253;
    exp_54_ram[443] = 0;
    exp_54_ram[444] = 0;
    exp_54_ram[445] = 251;
    exp_54_ram[446] = 67;
    exp_54_ram[447] = 3;
    exp_54_ram[448] = 3;
    exp_54_ram[449] = 0;
    exp_54_ram[450] = 0;
    exp_54_ram[451] = 31;
    exp_54_ram[452] = 0;
    exp_54_ram[453] = 0;
    exp_54_ram[454] = 0;
    exp_54_ram[455] = 0;
    exp_54_ram[456] = 0;
    exp_54_ram[457] = 65;
    exp_54_ram[458] = 25;
    exp_54_ram[459] = 0;
    exp_54_ram[460] = 0;
    exp_54_ram[461] = 0;
    exp_54_ram[462] = 0;
    exp_54_ram[463] = 0;
    exp_54_ram[464] = 3;
    exp_54_ram[465] = 2;
    exp_54_ram[466] = 9;
    exp_54_ram[467] = 255;
    exp_54_ram[468] = 0;
    exp_54_ram[469] = 2;
    exp_54_ram[470] = 65;
    exp_54_ram[471] = 1;
    exp_54_ram[472] = 0;
    exp_54_ram[473] = 0;
    exp_54_ram[474] = 255;
    exp_54_ram[475] = 255;
    exp_54_ram[476] = 0;
    exp_54_ram[477] = 0;
    exp_54_ram[478] = 2;
    exp_54_ram[479] = 0;
    exp_54_ram[480] = 0;
    exp_54_ram[481] = 0;
    exp_54_ram[482] = 0;
    exp_54_ram[483] = 0;
    exp_54_ram[484] = 0;
    exp_54_ram[485] = 0;
    exp_54_ram[486] = 0;
    exp_54_ram[487] = 0;
    exp_54_ram[488] = 0;
    exp_54_ram[489] = 255;
    exp_54_ram[490] = 255;
    exp_54_ram[491] = 67;
    exp_54_ram[492] = 0;
    exp_54_ram[493] = 65;
    exp_54_ram[494] = 0;
    exp_54_ram[495] = 1;
    exp_54_ram[496] = 0;
    exp_54_ram[497] = 0;
    exp_54_ram[498] = 237;
    exp_54_ram[499] = 253;
    exp_54_ram[500] = 0;
    exp_54_ram[501] = 0;
    exp_54_ram[502] = 249;
    exp_54_ram[503] = 0;
    exp_54_ram[504] = 0;
    exp_54_ram[505] = 0;
    exp_54_ram[506] = 235;
    exp_54_ram[507] = 0;
    exp_54_ram[508] = 0;
    exp_54_ram[509] = 0;
    exp_54_ram[510] = 0;
    exp_54_ram[511] = 0;
    exp_54_ram[512] = 0;
    exp_54_ram[513] = 0;
    exp_54_ram[514] = 254;
    exp_54_ram[515] = 0;
    exp_54_ram[516] = 6;
    exp_54_ram[517] = 6;
    exp_54_ram[518] = 0;
    exp_54_ram[519] = 0;
    exp_54_ram[520] = 255;
    exp_54_ram[521] = 2;
    exp_54_ram[522] = 0;
    exp_54_ram[523] = 0;
    exp_54_ram[524] = 0;
    exp_54_ram[525] = 0;
    exp_54_ram[526] = 0;
    exp_54_ram[527] = 254;
    exp_54_ram[528] = 0;
    exp_54_ram[529] = 0;
    exp_54_ram[530] = 64;
    exp_54_ram[531] = 0;
    exp_54_ram[532] = 0;
    exp_54_ram[533] = 0;
    exp_54_ram[534] = 254;
    exp_54_ram[535] = 0;
    exp_54_ram[536] = 0;
    exp_54_ram[537] = 251;
    exp_54_ram[538] = 0;
    exp_54_ram[539] = 0;
    exp_54_ram[540] = 64;
    exp_54_ram[541] = 0;
    exp_54_ram[542] = 64;
    exp_54_ram[543] = 249;
    exp_54_ram[544] = 64;
    exp_54_ram[545] = 0;
    exp_54_ram[546] = 249;
    exp_54_ram[547] = 64;
    exp_54_ram[548] = 0;
    exp_54_ram[549] = 0;
    exp_54_ram[550] = 0;
    exp_54_ram[551] = 0;
    exp_54_ram[552] = 247;
    exp_54_ram[553] = 0;
    exp_54_ram[554] = 0;
    exp_54_ram[555] = 64;
    exp_54_ram[556] = 254;
    exp_54_ram[557] = 64;
    exp_54_ram[558] = 246;
    exp_54_ram[559] = 64;
    exp_54_ram[560] = 0;
    exp_54_ram[561] = 2;
    exp_54_ram[562] = 2;
    exp_54_ram[563] = 64;
    exp_54_ram[564] = 0;
    exp_54_ram[565] = 254;
    exp_54_ram[566] = 0;
    exp_54_ram[567] = 0;
    exp_54_ram[568] = 0;
    exp_54_ram[569] = 0;
    exp_54_ram[570] = 0;
    exp_54_ram[571] = 0;
    exp_54_ram[572] = 0;
    exp_54_ram[573] = 0;
    exp_54_ram[574] = 254;
    exp_54_ram[575] = 2;
    exp_54_ram[576] = 2;
    exp_54_ram[577] = 64;
    exp_54_ram[578] = 0;
    exp_54_ram[579] = 254;
    exp_54_ram[580] = 0;
    exp_54_ram[581] = 0;
    exp_54_ram[582] = 0;
    exp_54_ram[583] = 0;
    exp_54_ram[584] = 0;
    exp_54_ram[585] = 0;
    exp_54_ram[586] = 0;
    exp_54_ram[587] = 0;
    exp_54_ram[588] = 254;
    exp_54_ram[589] = 0;
    exp_54_ram[590] = 2;
    exp_54_ram[591] = 15;
    exp_54_ram[592] = 0;
    exp_54_ram[593] = 0;
    exp_54_ram[594] = 0;
    exp_54_ram[595] = 2;
    exp_54_ram[596] = 64;
    exp_54_ram[597] = 0;
    exp_54_ram[598] = 165;
    exp_54_ram[599] = 0;
    exp_54_ram[600] = 0;
    exp_54_ram[601] = 64;
    exp_54_ram[602] = 0;
    exp_54_ram[603] = 1;
    exp_54_ram[604] = 1;
    exp_54_ram[605] = 252;
    exp_54_ram[606] = 1;
    exp_54_ram[607] = 252;
    exp_54_ram[608] = 99;
    exp_54_ram[609] = 46;
    exp_54_ram[610] = 0;
    exp_54_ram[611] = 115;
    exp_54_ram[612] = 0;
    exp_54_ram[613] = 101;
    exp_54_ram[614] = 0;
    exp_54_ram[615] = 32;
    exp_54_ram[616] = 32;
    exp_54_ram[617] = 48;
    exp_54_ram[618] = 49;
    exp_54_ram[619] = 32;
    exp_54_ram[620] = 48;
    exp_54_ram[621] = 0;
    exp_54_ram[622] = 97;
    exp_54_ram[623] = 0;
    exp_54_ram[624] = 32;
    exp_54_ram[625] = 32;
    exp_54_ram[626] = 48;
    exp_54_ram[627] = 49;
    exp_54_ram[628] = 32;
    exp_54_ram[629] = 48;
    exp_54_ram[630] = 0;
    exp_54_ram[631] = 97;
    exp_54_ram[632] = 0;
    exp_54_ram[633] = 97;
    exp_54_ram[634] = 0;
    exp_54_ram[635] = 97;
    exp_54_ram[636] = 0;
    exp_54_ram[637] = 97;
    exp_54_ram[638] = 0;
    exp_54_ram[639] = 97;
    exp_54_ram[640] = 0;
    exp_54_ram[641] = 97;
    exp_54_ram[642] = 0;
    exp_54_ram[643] = 97;
    exp_54_ram[644] = 0;
    exp_54_ram[645] = 97;
    exp_54_ram[646] = 0;
    exp_54_ram[647] = 32;
    exp_54_ram[648] = 32;
    exp_54_ram[649] = 48;
    exp_54_ram[650] = 49;
    exp_54_ram[651] = 32;
    exp_54_ram[652] = 48;
    exp_54_ram[653] = 0;
    exp_54_ram[654] = 102;
    exp_54_ram[655] = 0;
    exp_54_ram[656] = 102;
    exp_54_ram[657] = 0;
    exp_54_ram[658] = 102;
    exp_54_ram[659] = 0;
    exp_54_ram[660] = 115;
    exp_54_ram[661] = 0;
    exp_54_ram[662] = 2;
    exp_54_ram[663] = 3;
    exp_54_ram[664] = 4;
    exp_54_ram[665] = 4;
    exp_54_ram[666] = 5;
    exp_54_ram[667] = 5;
    exp_54_ram[668] = 5;
    exp_54_ram[669] = 5;
    exp_54_ram[670] = 6;
    exp_54_ram[671] = 6;
    exp_54_ram[672] = 6;
    exp_54_ram[673] = 6;
    exp_54_ram[674] = 6;
    exp_54_ram[675] = 6;
    exp_54_ram[676] = 6;
    exp_54_ram[677] = 6;
    exp_54_ram[678] = 7;
    exp_54_ram[679] = 7;
    exp_54_ram[680] = 7;
    exp_54_ram[681] = 7;
    exp_54_ram[682] = 7;
    exp_54_ram[683] = 7;
    exp_54_ram[684] = 7;
    exp_54_ram[685] = 7;
    exp_54_ram[686] = 7;
    exp_54_ram[687] = 7;
    exp_54_ram[688] = 7;
    exp_54_ram[689] = 7;
    exp_54_ram[690] = 7;
    exp_54_ram[691] = 7;
    exp_54_ram[692] = 7;
    exp_54_ram[693] = 7;
    exp_54_ram[694] = 8;
    exp_54_ram[695] = 8;
    exp_54_ram[696] = 8;
    exp_54_ram[697] = 8;
    exp_54_ram[698] = 8;
    exp_54_ram[699] = 8;
    exp_54_ram[700] = 8;
    exp_54_ram[701] = 8;
    exp_54_ram[702] = 8;
    exp_54_ram[703] = 8;
    exp_54_ram[704] = 8;
    exp_54_ram[705] = 8;
    exp_54_ram[706] = 8;
    exp_54_ram[707] = 8;
    exp_54_ram[708] = 8;
    exp_54_ram[709] = 8;
    exp_54_ram[710] = 8;
    exp_54_ram[711] = 8;
    exp_54_ram[712] = 8;
    exp_54_ram[713] = 8;
    exp_54_ram[714] = 8;
    exp_54_ram[715] = 8;
    exp_54_ram[716] = 8;
    exp_54_ram[717] = 8;
    exp_54_ram[718] = 8;
    exp_54_ram[719] = 8;
    exp_54_ram[720] = 8;
    exp_54_ram[721] = 8;
    exp_54_ram[722] = 8;
    exp_54_ram[723] = 8;
    exp_54_ram[724] = 8;
    exp_54_ram[725] = 8;
    exp_54_ram[726] = 0;
    exp_54_ram[727] = 0;
    exp_54_ram[728] = 0;
    exp_54_ram[729] = 0;
    exp_54_ram[730] = 0;
    exp_54_ram[731] = 0;
    exp_54_ram[732] = 0;
    exp_54_ram[733] = 0;
    exp_54_ram[734] = 254;
    exp_54_ram[735] = 255;
    exp_54_ram[736] = 0;
    exp_54_ram[737] = 0;
    exp_54_ram[738] = 247;
    exp_54_ram[739] = 0;
    exp_54_ram[740] = 0;
    exp_54_ram[741] = 252;
    exp_54_ram[742] = 0;
    exp_54_ram[743] = 0;
    exp_54_ram[744] = 0;
    exp_54_ram[745] = 0;
    exp_54_ram[746] = 0;
    exp_54_ram[747] = 1;
    exp_54_ram[748] = 0;
    exp_54_ram[749] = 0;
    exp_54_ram[750] = 0;
    exp_54_ram[751] = 0;
    exp_54_ram[752] = 6;
    exp_54_ram[753] = 0;
    exp_54_ram[754] = 0;
    exp_54_ram[755] = 0;
    exp_54_ram[756] = 2;
    exp_54_ram[757] = 0;
    exp_54_ram[758] = 1;
    exp_54_ram[759] = 1;
    exp_54_ram[760] = 255;
    exp_54_ram[761] = 255;
    exp_54_ram[762] = 255;
    exp_54_ram[763] = 255;
    exp_54_ram[764] = 255;
    exp_54_ram[765] = 255;
    exp_54_ram[766] = 255;
    exp_54_ram[767] = 64;
    exp_54_ram[768] = 253;
    exp_54_ram[769] = 0;
    exp_54_ram[770] = 255;
    exp_54_ram[771] = 0;
    exp_54_ram[772] = 0;
    exp_54_ram[773] = 0;
    exp_54_ram[774] = 64;
    exp_54_ram[775] = 3;
    exp_54_ram[776] = 0;
    exp_54_ram[777] = 0;
    exp_54_ram[778] = 0;
    exp_54_ram[779] = 0;
    exp_54_ram[780] = 0;
    exp_54_ram[781] = 2;
    exp_54_ram[782] = 0;
    exp_54_ram[783] = 0;
    exp_54_ram[784] = 0;
    exp_54_ram[785] = 0;
    exp_54_ram[786] = 0;
    exp_54_ram[787] = 1;
    exp_54_ram[788] = 252;
    exp_54_ram[789] = 0;
    exp_54_ram[790] = 0;
    exp_54_ram[791] = 0;
    exp_54_ram[792] = 0;
    exp_54_ram[793] = 1;
    exp_54_ram[794] = 252;
    exp_54_ram[795] = 0;
    exp_54_ram[796] = 0;
    exp_54_ram[797] = 2;
    exp_54_ram[798] = 254;
    exp_54_ram[799] = 128;
    exp_54_ram[800] = 239;
    exp_54_ram[801] = 8;
    exp_54_ram[802] = 0;
    exp_54_ram[803] = 0;
    exp_54_ram[804] = 0;
    exp_54_ram[805] = 0;
    exp_54_ram[806] = 0;
    exp_54_ram[807] = 0;
    exp_54_ram[808] = 2;
    exp_54_ram[809] = 64;
    exp_54_ram[810] = 0;
    exp_54_ram[811] = 0;
    exp_54_ram[812] = 255;
    exp_54_ram[813] = 0;
    exp_54_ram[814] = 0;
    exp_54_ram[815] = 0;
    exp_54_ram[816] = 0;
    exp_54_ram[817] = 0;
    exp_54_ram[818] = 252;
    exp_54_ram[819] = 0;
    exp_54_ram[820] = 0;
    exp_54_ram[821] = 252;
    exp_54_ram[822] = 0;
    exp_54_ram[823] = 0;
    exp_54_ram[824] = 0;
    exp_54_ram[825] = 4;
    exp_54_ram[826] = 255;
    exp_54_ram[827] = 6;
    exp_54_ram[828] = 0;
    exp_54_ram[829] = 0;
    exp_54_ram[830] = 0;
    exp_54_ram[831] = 182;
    exp_54_ram[832] = 0;
    exp_54_ram[833] = 0;
    exp_54_ram[834] = 25;
    exp_54_ram[835] = 0;
    exp_54_ram[836] = 181;
    exp_54_ram[837] = 0;
    exp_54_ram[838] = 0;
    exp_54_ram[839] = 0;
    exp_54_ram[840] = 0;
    exp_54_ram[841] = 1;
    exp_54_ram[842] = 0;
    exp_54_ram[843] = 0;
    exp_54_ram[844] = 0;
    exp_54_ram[845] = 0;
    exp_54_ram[846] = 255;
    exp_54_ram[847] = 255;
    exp_54_ram[848] = 4;
    exp_54_ram[849] = 255;
    exp_54_ram[850] = 0;
    exp_54_ram[851] = 1;
    exp_54_ram[852] = 2;
    exp_54_ram[853] = 0;
    exp_54_ram[854] = 1;
    exp_54_ram[855] = 2;
    exp_54_ram[856] = 255;
    exp_54_ram[857] = 0;
    exp_54_ram[858] = 247;
    exp_54_ram[859] = 0;
    exp_54_ram[860] = 0;
    exp_54_ram[861] = 1;
    exp_54_ram[862] = 0;
    exp_54_ram[863] = 1;
    exp_54_ram[864] = 0;
    exp_54_ram[865] = 1;
    exp_54_ram[866] = 0;
    exp_54_ram[867] = 0;
    exp_54_ram[868] = 128;
    exp_54_ram[869] = 0;
    exp_54_ram[870] = 0;
    exp_54_ram[871] = 0;
    exp_54_ram[872] = 0;
    exp_54_ram[873] = 0;
    exp_54_ram[874] = 0;
    exp_54_ram[875] = 0;
    exp_54_ram[876] = 0;
    exp_54_ram[877] = 64;
    exp_54_ram[878] = 0;
    exp_54_ram[879] = 64;
    exp_54_ram[880] = 255;
    exp_54_ram[881] = 64;
    exp_54_ram[882] = 0;
    exp_54_ram[883] = 133;
    exp_54_ram[884] = 0;
    exp_54_ram[885] = 1;
    exp_54_ram[886] = 0;
    exp_54_ram[887] = 254;
    exp_54_ram[888] = 1;
    exp_54_ram[889] = 1;
    exp_54_ram[890] = 0;
    exp_54_ram[891] = 0;
    exp_54_ram[892] = 0;
    exp_54_ram[893] = 1;
    exp_54_ram[894] = 1;
    exp_54_ram[895] = 1;
    exp_54_ram[896] = 0;
    exp_54_ram[897] = 1;
    exp_54_ram[898] = 0;
    exp_54_ram[899] = 123;
    exp_54_ram[900] = 0;
    exp_54_ram[901] = 0;
    exp_54_ram[902] = 118;
    exp_54_ram[903] = 24;
    exp_54_ram[904] = 4;
    exp_54_ram[905] = 1;
    exp_54_ram[906] = 0;
    exp_54_ram[907] = 0;
    exp_54_ram[908] = 24;
    exp_54_ram[909] = 6;
    exp_54_ram[910] = 0;
    exp_54_ram[911] = 0;
    exp_54_ram[912] = 239;
    exp_54_ram[913] = 0;
    exp_54_ram[914] = 154;
    exp_54_ram[915] = 0;
    exp_54_ram[916] = 1;
    exp_54_ram[917] = 1;
    exp_54_ram[918] = 0;
    exp_54_ram[919] = 0;
    exp_54_ram[920] = 253;
    exp_54_ram[921] = 0;
    exp_54_ram[922] = 231;
    exp_54_ram[923] = 0;
    exp_54_ram[924] = 0;
    exp_54_ram[925] = 22;
    exp_54_ram[926] = 151;
    exp_54_ram[927] = 0;
    exp_54_ram[928] = 1;
    exp_54_ram[929] = 1;
    exp_54_ram[930] = 0;
    exp_54_ram[931] = 0;
    exp_54_ram[932] = 249;
    exp_54_ram[933] = 0;
    exp_54_ram[934] = 0;
    exp_54_ram[935] = 0;
    exp_54_ram[936] = 0;
    exp_54_ram[937] = 64;
    exp_54_ram[938] = 0;
    exp_54_ram[939] = 0;
    exp_54_ram[940] = 0;
    exp_54_ram[941] = 64;
    exp_54_ram[942] = 0;
    exp_54_ram[943] = 0;
    exp_54_ram[944] = 0;
    exp_54_ram[945] = 65;
    exp_54_ram[946] = 65;
    exp_54_ram[947] = 0;
    exp_54_ram[948] = 0;
    exp_54_ram[949] = 0;
    exp_54_ram[950] = 0;
    exp_54_ram[951] = 0;
    exp_54_ram[952] = 65;
    exp_54_ram[953] = 0;
    exp_54_ram[954] = 0;
    exp_54_ram[955] = 0;
    exp_54_ram[956] = 24;
    exp_54_ram[957] = 255;
    exp_54_ram[958] = 0;
    exp_54_ram[959] = 143;
    exp_54_ram[960] = 0;
    exp_54_ram[961] = 65;
    exp_54_ram[962] = 0;
    exp_54_ram[963] = 0;
    exp_54_ram[964] = 1;
    exp_54_ram[965] = 0;
    exp_54_ram[966] = 1;
    exp_54_ram[967] = 0;
    exp_54_ram[968] = 1;
    exp_54_ram[969] = 0;
    exp_54_ram[970] = 1;
    exp_54_ram[971] = 1;
    exp_54_ram[972] = 1;
    exp_54_ram[973] = 0;
    exp_54_ram[974] = 0;
    exp_54_ram[975] = 0;
    exp_54_ram[976] = 0;
    exp_54_ram[977] = 2;
    exp_54_ram[978] = 0;
    exp_54_ram[979] = 255;
    exp_54_ram[980] = 0;
    exp_54_ram[981] = 0;
    exp_54_ram[982] = 0;
    exp_54_ram[983] = 227;
    exp_54_ram[984] = 0;
    exp_54_ram[985] = 246;
    exp_54_ram[986] = 0;
    exp_54_ram[987] = 146;
    exp_54_ram[988] = 0;
    exp_54_ram[989] = 255;
    exp_54_ram[990] = 0;
    exp_54_ram[991] = 0;
    exp_54_ram[992] = 0;
    exp_54_ram[993] = 0;
    exp_54_ram[994] = 0;
    exp_54_ram[995] = 0;
    exp_54_ram[996] = 0;
    exp_54_ram[997] = 1;
    exp_54_ram[998] = 0;
    exp_54_ram[999] = 255;
    exp_54_ram[1000] = 0;
    exp_54_ram[1001] = 0;
    exp_54_ram[1002] = 0;
    exp_54_ram[1003] = 1;
    exp_54_ram[1004] = 0;
    exp_54_ram[1005] = 0;
    exp_54_ram[1006] = 221;
    exp_54_ram[1007] = 0;
    exp_54_ram[1008] = 246;
    exp_54_ram[1009] = 0;
    exp_54_ram[1010] = 0;
    exp_54_ram[1011] = 140;
    exp_54_ram[1012] = 64;
    exp_54_ram[1013] = 0;
    exp_54_ram[1014] = 64;
    exp_54_ram[1015] = 255;
    exp_54_ram[1016] = 64;
    exp_54_ram[1017] = 0;
    exp_54_ram[1018] = 0;
    exp_54_ram[1019] = 0;
    exp_54_ram[1020] = 0;
    exp_54_ram[1021] = 0;
    exp_54_ram[1022] = 0;
    exp_54_ram[1023] = 1;
    exp_54_ram[1024] = 0;
    exp_54_ram[1025] = 249;
    exp_54_ram[1026] = 0;
    exp_54_ram[1027] = 6;
    exp_54_ram[1028] = 1;
    exp_54_ram[1029] = 0;
    exp_54_ram[1030] = 247;
    exp_54_ram[1031] = 1;
    exp_54_ram[1032] = 6;
    exp_54_ram[1033] = 6;
    exp_54_ram[1034] = 7;
    exp_54_ram[1035] = 5;
    exp_54_ram[1036] = 5;
    exp_54_ram[1037] = 184;
    exp_54_ram[1038] = 0;
    exp_54_ram[1039] = 2;
    exp_54_ram[1040] = 248;
    exp_54_ram[1041] = 2;
    exp_54_ram[1042] = 182;
    exp_54_ram[1043] = 1;
    exp_54_ram[1044] = 0;
    exp_54_ram[1045] = 251;
    exp_54_ram[1046] = 0;
    exp_54_ram[1047] = 0;
    exp_54_ram[1048] = 1;
    exp_54_ram[1049] = 2;
    exp_54_ram[1050] = 0;
    exp_54_ram[1051] = 0;
    exp_54_ram[1052] = 251;
    exp_54_ram[1053] = 180;
    exp_54_ram[1054] = 1;
    exp_54_ram[1055] = 1;
    exp_54_ram[1056] = 0;
    exp_54_ram[1057] = 0;
    exp_54_ram[1058] = 0;
    exp_54_ram[1059] = 0;
    exp_54_ram[1060] = 2;
    exp_54_ram[1061] = 0;
    exp_54_ram[1062] = 177;
    exp_54_ram[1063] = 1;
    exp_54_ram[1064] = 0;
    exp_54_ram[1065] = 0;
    exp_54_ram[1066] = 3;
    exp_54_ram[1067] = 104;
    exp_54_ram[1068] = 0;
    exp_54_ram[1069] = 0;
    exp_54_ram[1070] = 0;
    exp_54_ram[1071] = 1;
    exp_54_ram[1072] = 3;
    exp_54_ram[1073] = 0;
    exp_54_ram[1074] = 0;
    exp_54_ram[1075] = 0;
    exp_54_ram[1076] = 3;
    exp_54_ram[1077] = 0;
    exp_54_ram[1078] = 0;
    exp_54_ram[1079] = 101;
    exp_54_ram[1080] = 0;
    exp_54_ram[1081] = 0;
    exp_54_ram[1082] = 0;
    exp_54_ram[1083] = 1;
    exp_54_ram[1084] = 3;
    exp_54_ram[1085] = 0;
    exp_54_ram[1086] = 0;
    exp_54_ram[1087] = 0;
    exp_54_ram[1088] = 3;
    exp_54_ram[1089] = 0;
    exp_54_ram[1090] = 0;
    exp_54_ram[1091] = 98;
    exp_54_ram[1092] = 0;
    exp_54_ram[1093] = 0;
    exp_54_ram[1094] = 0;
    exp_54_ram[1095] = 1;
    exp_54_ram[1096] = 3;
    exp_54_ram[1097] = 0;
    exp_54_ram[1098] = 0;
    exp_54_ram[1099] = 0;
    exp_54_ram[1100] = 3;
    exp_54_ram[1101] = 0;
    exp_54_ram[1102] = 0;
    exp_54_ram[1103] = 95;
    exp_54_ram[1104] = 0;
    exp_54_ram[1105] = 0;
    exp_54_ram[1106] = 0;
    exp_54_ram[1107] = 1;
    exp_54_ram[1108] = 3;
    exp_54_ram[1109] = 0;
    exp_54_ram[1110] = 0;
    exp_54_ram[1111] = 62;
    exp_54_ram[1112] = 3;
    exp_54_ram[1113] = 0;
    exp_54_ram[1114] = 1;
    exp_54_ram[1115] = 118;
    exp_54_ram[1116] = 92;
    exp_54_ram[1117] = 0;
    exp_54_ram[1118] = 0;
    exp_54_ram[1119] = 0;
    exp_54_ram[1120] = 0;
    exp_54_ram[1121] = 6;
    exp_54_ram[1122] = 3;
    exp_54_ram[1123] = 0;
    exp_54_ram[1124] = 90;
    exp_54_ram[1125] = 0;
    exp_54_ram[1126] = 0;
    exp_54_ram[1127] = 0;
    exp_54_ram[1128] = 0;
    exp_54_ram[1129] = 0;
    exp_54_ram[1130] = 3;
    exp_54_ram[1131] = 0;
    exp_54_ram[1132] = 88;
    exp_54_ram[1133] = 0;
    exp_54_ram[1134] = 0;
    exp_54_ram[1135] = 0;
    exp_54_ram[1136] = 6;
    exp_54_ram[1137] = 3;
    exp_54_ram[1138] = 0;
    exp_54_ram[1139] = 0;
    exp_54_ram[1140] = 6;
    exp_54_ram[1141] = 6;
    exp_54_ram[1142] = 3;
    exp_54_ram[1143] = 0;
    exp_54_ram[1144] = 0;
    exp_54_ram[1145] = 0;
    exp_54_ram[1146] = 6;
    exp_54_ram[1147] = 5;
    exp_54_ram[1148] = 251;
    exp_54_ram[1149] = 5;
    exp_54_ram[1150] = 7;
    exp_54_ram[1151] = 0;
    exp_54_ram[1152] = 252;
    exp_54_ram[1153] = 3;
    exp_54_ram[1154] = 0;
    exp_54_ram[1155] = 2;
    exp_54_ram[1156] = 2;
    exp_54_ram[1157] = 3;
    exp_54_ram[1158] = 3;
    exp_54_ram[1159] = 3;
    exp_54_ram[1160] = 2;
    exp_54_ram[1161] = 3;
    exp_54_ram[1162] = 1;
    exp_54_ram[1163] = 1;
    exp_54_ram[1164] = 1;
    exp_54_ram[1165] = 0;
    exp_54_ram[1166] = 0;
    exp_54_ram[1167] = 0;
    exp_54_ram[1168] = 123;
    exp_54_ram[1169] = 0;
    exp_54_ram[1170] = 24;
    exp_54_ram[1171] = 0;
    exp_54_ram[1172] = 169;
    exp_54_ram[1173] = 0;
    exp_54_ram[1174] = 22;
    exp_54_ram[1175] = 0;
    exp_54_ram[1176] = 0;
    exp_54_ram[1177] = 216;
    exp_54_ram[1178] = 0;
    exp_54_ram[1179] = 0;
    exp_54_ram[1180] = 2;
    exp_54_ram[1181] = 64;
    exp_54_ram[1182] = 0;
    exp_54_ram[1183] = 1;
    exp_54_ram[1184] = 0;
    exp_54_ram[1185] = 64;
    exp_54_ram[1186] = 0;
    exp_54_ram[1187] = 252;
    exp_54_ram[1188] = 0;
    exp_54_ram[1189] = 0;
    exp_54_ram[1190] = 0;
    exp_54_ram[1191] = 24;
    exp_54_ram[1192] = 0;
    exp_54_ram[1193] = 0;
    exp_54_ram[1194] = 169;
    exp_54_ram[1195] = 0;
    exp_54_ram[1196] = 0;
    exp_54_ram[1197] = 0;
    exp_54_ram[1198] = 0;
    exp_54_ram[1199] = 211;
    exp_54_ram[1200] = 0;
    exp_54_ram[1201] = 2;
    exp_54_ram[1202] = 64;
    exp_54_ram[1203] = 0;
    exp_54_ram[1204] = 1;
    exp_54_ram[1205] = 1;
    exp_54_ram[1206] = 0;
    exp_54_ram[1207] = 64;
    exp_54_ram[1208] = 252;
    exp_54_ram[1209] = 0;
    exp_54_ram[1210] = 0;
    exp_54_ram[1211] = 24;
    exp_54_ram[1212] = 68;
    exp_54_ram[1213] = 0;
    exp_54_ram[1214] = 0;
    exp_54_ram[1215] = 0;
    exp_54_ram[1216] = 0;
    exp_54_ram[1217] = 0;
    exp_54_ram[1218] = 0;
    exp_54_ram[1219] = 225;
    exp_54_ram[1220] = 66;
    exp_54_ram[1221] = 0;
    exp_54_ram[1222] = 0;
    exp_54_ram[1223] = 0;
    exp_54_ram[1224] = 0;
    exp_54_ram[1225] = 3;
    exp_54_ram[1226] = 137;
    exp_54_ram[1227] = 64;
    exp_54_ram[1228] = 0;
    exp_54_ram[1229] = 0;
    exp_54_ram[1230] = 0;
    exp_54_ram[1231] = 0;
    exp_54_ram[1232] = 0;
    exp_54_ram[1233] = 1;
    exp_54_ram[1234] = 1;
    exp_54_ram[1235] = 1;
    exp_54_ram[1236] = 0;
    exp_54_ram[1237] = 0;
    exp_54_ram[1238] = 0;
    exp_54_ram[1239] = 211;
    exp_54_ram[1240] = 0;
    exp_54_ram[1241] = 1;
    exp_54_ram[1242] = 3;
    exp_54_ram[1243] = 0;
    exp_54_ram[1244] = 3;
    exp_54_ram[1245] = 3;
    exp_54_ram[1246] = 3;
    exp_54_ram[1247] = 2;
    exp_54_ram[1248] = 2;
    exp_54_ram[1249] = 2;
    exp_54_ram[1250] = 2;
    exp_54_ram[1251] = 1;
    exp_54_ram[1252] = 1;
    exp_54_ram[1253] = 1;
    exp_54_ram[1254] = 4;
    exp_54_ram[1255] = 0;
    exp_54_ram[1256] = 246;
    exp_54_ram[1257] = 9;
    exp_54_ram[1258] = 1;
    exp_54_ram[1259] = 0;
    exp_54_ram[1260] = 8;
    exp_54_ram[1261] = 9;
    exp_54_ram[1262] = 9;
    exp_54_ram[1263] = 1;
    exp_54_ram[1264] = 0;
    exp_54_ram[1265] = 2;
    exp_54_ram[1266] = 0;
    exp_54_ram[1267] = 3;
    exp_54_ram[1268] = 0;
    exp_54_ram[1269] = 8;
    exp_54_ram[1270] = 4;
    exp_54_ram[1271] = 8;
    exp_54_ram[1272] = 9;
    exp_54_ram[1273] = 5;
    exp_54_ram[1274] = 4;
    exp_54_ram[1275] = 5;
    exp_54_ram[1276] = 2;
    exp_54_ram[1277] = 2;
    exp_54_ram[1278] = 4;
    exp_54_ram[1279] = 251;
    exp_54_ram[1280] = 0;
    exp_54_ram[1281] = 157;
    exp_54_ram[1282] = 0;
    exp_54_ram[1283] = 0;
    exp_54_ram[1284] = 3;
    exp_54_ram[1285] = 222;
    exp_54_ram[1286] = 5;
    exp_54_ram[1287] = 4;
    exp_54_ram[1288] = 2;
    exp_54_ram[1289] = 3;
    exp_54_ram[1290] = 64;
    exp_54_ram[1291] = 0;
    exp_54_ram[1292] = 4;
    exp_54_ram[1293] = 248;
    exp_54_ram[1294] = 0;
    exp_54_ram[1295] = 154;
    exp_54_ram[1296] = 0;
    exp_54_ram[1297] = 2;
    exp_54_ram[1298] = 0;
    exp_54_ram[1299] = 0;
    exp_54_ram[1300] = 0;
    exp_54_ram[1301] = 5;
    exp_54_ram[1302] = 6;
    exp_54_ram[1303] = 7;
    exp_54_ram[1304] = 6;
    exp_54_ram[1305] = 7;
    exp_54_ram[1306] = 6;
    exp_54_ram[1307] = 4;
    exp_54_ram[1308] = 244;
    exp_54_ram[1309] = 0;
    exp_54_ram[1310] = 150;
    exp_54_ram[1311] = 0;
    exp_54_ram[1312] = 0;
    exp_54_ram[1313] = 5;
    exp_54_ram[1314] = 215;
    exp_54_ram[1315] = 7;
    exp_54_ram[1316] = 6;
    exp_54_ram[1317] = 2;
    exp_54_ram[1318] = 5;
    exp_54_ram[1319] = 64;
    exp_54_ram[1320] = 0;
    exp_54_ram[1321] = 6;
    exp_54_ram[1322] = 240;
    exp_54_ram[1323] = 0;
    exp_54_ram[1324] = 146;
    exp_54_ram[1325] = 0;
    exp_54_ram[1326] = 0;
    exp_54_ram[1327] = 2;
    exp_54_ram[1328] = 0;
    exp_54_ram[1329] = 0;
    exp_54_ram[1330] = 238;
    exp_54_ram[1331] = 0;
    exp_54_ram[1332] = 144;
    exp_54_ram[1333] = 2;
    exp_54_ram[1334] = 0;
    exp_54_ram[1335] = 0;
    exp_54_ram[1336] = 0;
    exp_54_ram[1337] = 1;
    exp_54_ram[1338] = 0;
    exp_54_ram[1339] = 0;
    exp_54_ram[1340] = 0;
    exp_54_ram[1341] = 0;
    exp_54_ram[1342] = 0;
    exp_54_ram[1343] = 9;
    exp_54_ram[1344] = 9;
    exp_54_ram[1345] = 9;
    exp_54_ram[1346] = 9;
    exp_54_ram[1347] = 8;
    exp_54_ram[1348] = 8;
    exp_54_ram[1349] = 8;
    exp_54_ram[1350] = 10;
    exp_54_ram[1351] = 0;
    exp_54_ram[1352] = 248;
    exp_54_ram[1353] = 0;
    exp_54_ram[1354] = 7;
    exp_54_ram[1355] = 2;
    exp_54_ram[1356] = 0;
    exp_54_ram[1357] = 3;
    exp_54_ram[1358] = 6;
    exp_54_ram[1359] = 6;
    exp_54_ram[1360] = 6;
    exp_54_ram[1361] = 7;
    exp_54_ram[1362] = 230;
    exp_54_ram[1363] = 2;
    exp_54_ram[1364] = 3;
    exp_54_ram[1365] = 0;
    exp_54_ram[1366] = 2;
    exp_54_ram[1367] = 229;
    exp_54_ram[1368] = 0;
    exp_54_ram[1369] = 135;
    exp_54_ram[1370] = 0;
    exp_54_ram[1371] = 0;
    exp_54_ram[1372] = 7;
    exp_54_ram[1373] = 255;
    exp_54_ram[1374] = 31;
    exp_54_ram[1375] = 0;
    exp_54_ram[1376] = 0;
    exp_54_ram[1377] = 255;
    exp_54_ram[1378] = 0;
    exp_54_ram[1379] = 0;
    exp_54_ram[1380] = 0;
    exp_54_ram[1381] = 0;
    exp_54_ram[1382] = 0;
    exp_54_ram[1383] = 198;
    exp_54_ram[1384] = 2;
    exp_54_ram[1385] = 0;
    exp_54_ram[1386] = 0;
    exp_54_ram[1387] = 224;
    exp_54_ram[1388] = 7;
    exp_54_ram[1389] = 0;
    exp_54_ram[1390] = 2;
    exp_54_ram[1391] = 7;
    exp_54_ram[1392] = 0;
    exp_54_ram[1393] = 7;
    exp_54_ram[1394] = 7;
    exp_54_ram[1395] = 6;
    exp_54_ram[1396] = 0;
    exp_54_ram[1397] = 7;
    exp_54_ram[1398] = 8;
    exp_54_ram[1399] = 0;
    exp_54_ram[1400] = 250;
    exp_54_ram[1401] = 2;
    exp_54_ram[1402] = 3;
    exp_54_ram[1403] = 0;
    exp_54_ram[1404] = 220;
    exp_54_ram[1405] = 0;
    exp_54_ram[1406] = 218;
    exp_54_ram[1407] = 0;
    exp_54_ram[1408] = 0;
    exp_54_ram[1409] = 0;
    exp_54_ram[1410] = 225;
    exp_54_ram[1411] = 64;
    exp_54_ram[1412] = 0;
    exp_54_ram[1413] = 64;
    exp_54_ram[1414] = 0;
    exp_54_ram[1415] = 247;
    exp_54_ram[1416] = 2;
    exp_54_ram[1417] = 2;
    exp_54_ram[1418] = 3;
    exp_54_ram[1419] = 0;
    exp_54_ram[1420] = 216;
    exp_54_ram[1421] = 0;
    exp_54_ram[1422] = 214;
    exp_54_ram[1423] = 2;
    exp_54_ram[1424] = 247;
    exp_54_ram[1425] = 2;
    exp_54_ram[1426] = 247;
    exp_54_ram[1427] = 249;
    exp_54_ram[1428] = 0;
    exp_54_ram[1429] = 0;
    exp_54_ram[1430] = 3;
    exp_54_ram[1431] = 6;
    exp_54_ram[1432] = 186;
    exp_54_ram[1433] = 3;
    exp_54_ram[1434] = 2;
    exp_54_ram[1435] = 0;
    exp_54_ram[1436] = 212;
    exp_54_ram[1437] = 0;
    exp_54_ram[1438] = 210;
    exp_54_ram[1439] = 6;
    exp_54_ram[1440] = 7;
    exp_54_ram[1441] = 0;
    exp_54_ram[1442] = 0;
    exp_54_ram[1443] = 0;
    exp_54_ram[1444] = 252;
    exp_54_ram[1445] = 0;
    exp_54_ram[1446] = 2;
    exp_54_ram[1447] = 2;
    exp_54_ram[1448] = 182;
    exp_54_ram[1449] = 0;
    exp_54_ram[1450] = 0;
    exp_54_ram[1451] = 253;
    exp_54_ram[1452] = 2;
    exp_54_ram[1453] = 208;
    exp_54_ram[1454] = 3;
    exp_54_ram[1455] = 253;
    exp_54_ram[1456] = 3;
    exp_54_ram[1457] = 4;
    exp_54_ram[1458] = 0;
    exp_54_ram[1459] = 251;
    exp_54_ram[1460] = 4;
    exp_54_ram[1461] = 5;
    exp_54_ram[1462] = 0;
    exp_54_ram[1463] = 0;
    exp_54_ram[1464] = 4;
    exp_54_ram[1465] = 0;
    exp_54_ram[1466] = 0;
    exp_54_ram[1467] = 4;
    exp_54_ram[1468] = 3;
    exp_54_ram[1469] = 245;
    exp_54_ram[1470] = 0;
    exp_54_ram[1471] = 0;
    exp_54_ram[1472] = 0;
    exp_54_ram[1473] = 225;
    exp_54_ram[1474] = 1;
    exp_54_ram[1475] = 0;
    exp_54_ram[1476] = 0;
    exp_54_ram[1477] = 0;
    exp_54_ram[1478] = 174;
    exp_54_ram[1479] = 0;
    exp_54_ram[1480] = 0;
    exp_54_ram[1481] = 2;
    exp_54_ram[1482] = 253;
    exp_54_ram[1483] = 200;
    exp_54_ram[1484] = 0;
    exp_54_ram[1485] = 0;
    exp_54_ram[1486] = 241;
    exp_54_ram[1487] = 253;
    exp_54_ram[1488] = 2;
    exp_54_ram[1489] = 4;
    exp_54_ram[1490] = 253;
    exp_54_ram[1491] = 4;
    exp_54_ram[1492] = 4;
    exp_54_ram[1493] = 4;
    exp_54_ram[1494] = 3;
    exp_54_ram[1495] = 5;
    exp_54_ram[1496] = 0;
    exp_54_ram[1497] = 255;
    exp_54_ram[1498] = 0;
    exp_54_ram[1499] = 246;
    exp_54_ram[1500] = 0;
    exp_54_ram[1501] = 1;
    exp_54_ram[1502] = 136;
    exp_54_ram[1503] = 255;
    exp_54_ram[1504] = 0;
    exp_54_ram[1505] = 0;
    exp_54_ram[1506] = 1;
    exp_54_ram[1507] = 0;
    exp_54_ram[1508] = 152;
    exp_54_ram[1509] = 190;
    exp_54_ram[1510] = 0;
    exp_54_ram[1511] = 152;
    exp_54_ram[1512] = 189;
    exp_54_ram[1513] = 0;
    exp_54_ram[1514] = 0;
    exp_54_ram[1515] = 1;
    exp_54_ram[1516] = 0;
    exp_54_ram[1517] = 250;
    exp_54_ram[1518] = 4;
    exp_54_ram[1519] = 4;
    exp_54_ram[1520] = 5;
    exp_54_ram[1521] = 5;
    exp_54_ram[1522] = 5;
    exp_54_ram[1523] = 5;
    exp_54_ram[1524] = 5;
    exp_54_ram[1525] = 5;
    exp_54_ram[1526] = 6;
    exp_54_ram[1527] = 0;
    exp_54_ram[1528] = 153;
    exp_54_ram[1529] = 185;
    exp_54_ram[1530] = 7;
    exp_54_ram[1531] = 252;
    exp_54_ram[1532] = 0;
    exp_54_ram[1533] = 250;
    exp_54_ram[1534] = 1;
    exp_54_ram[1535] = 250;
    exp_54_ram[1536] = 0;
    exp_54_ram[1537] = 250;
    exp_54_ram[1538] = 1;
    exp_54_ram[1539] = 250;
    exp_54_ram[1540] = 250;
    exp_54_ram[1541] = 255;
    exp_54_ram[1542] = 252;
    exp_54_ram[1543] = 250;
    exp_54_ram[1544] = 0;
    exp_54_ram[1545] = 207;
    exp_54_ram[1546] = 0;
    exp_54_ram[1547] = 0;
    exp_54_ram[1548] = 250;
    exp_54_ram[1549] = 250;
    exp_54_ram[1550] = 250;
    exp_54_ram[1551] = 0;
    exp_54_ram[1552] = 252;
    exp_54_ram[1553] = 0;
    exp_54_ram[1554] = 0;
    exp_54_ram[1555] = 153;
    exp_54_ram[1556] = 0;
    exp_54_ram[1557] = 193;
    exp_54_ram[1558] = 0;
    exp_54_ram[1559] = 0;
    exp_54_ram[1560] = 0;
    exp_54_ram[1561] = 155;
    exp_54_ram[1562] = 177;
    exp_54_ram[1563] = 103;
    exp_54_ram[1564] = 250;
    exp_54_ram[1565] = 0;
    exp_54_ram[1566] = 229;
    exp_54_ram[1567] = 0;
    exp_54_ram[1568] = 0;
    exp_54_ram[1569] = 248;
    exp_54_ram[1570] = 0;
    exp_54_ram[1571] = 0;
    exp_54_ram[1572] = 156;
    exp_54_ram[1573] = 0;
    exp_54_ram[1574] = 189;
    exp_54_ram[1575] = 0;
    exp_54_ram[1576] = 0;
    exp_54_ram[1577] = 0;
    exp_54_ram[1578] = 157;
    exp_54_ram[1579] = 173;
    exp_54_ram[1580] = 98;
    exp_54_ram[1581] = 250;
    exp_54_ram[1582] = 0;
    exp_54_ram[1583] = 220;
    exp_54_ram[1584] = 0;
    exp_54_ram[1585] = 0;
    exp_54_ram[1586] = 243;
    exp_54_ram[1587] = 0;
    exp_54_ram[1588] = 0;
    exp_54_ram[1589] = 153;
    exp_54_ram[1590] = 0;
    exp_54_ram[1591] = 185;
    exp_54_ram[1592] = 0;
    exp_54_ram[1593] = 0;
    exp_54_ram[1594] = 0;
    exp_54_ram[1595] = 158;
    exp_54_ram[1596] = 168;
    exp_54_ram[1597] = 94;
    exp_54_ram[1598] = 250;
    exp_54_ram[1599] = 0;
    exp_54_ram[1600] = 230;
    exp_54_ram[1601] = 0;
    exp_54_ram[1602] = 0;
    exp_54_ram[1603] = 156;
    exp_54_ram[1604] = 0;
    exp_54_ram[1605] = 181;
    exp_54_ram[1606] = 0;
    exp_54_ram[1607] = 0;
    exp_54_ram[1608] = 0;
    exp_54_ram[1609] = 158;
    exp_54_ram[1610] = 165;
    exp_54_ram[1611] = 91;
    exp_54_ram[1612] = 7;
    exp_54_ram[1613] = 252;
    exp_54_ram[1614] = 0;
    exp_54_ram[1615] = 250;
    exp_54_ram[1616] = 1;
    exp_54_ram[1617] = 250;
    exp_54_ram[1618] = 0;
    exp_54_ram[1619] = 250;
    exp_54_ram[1620] = 1;
    exp_54_ram[1621] = 250;
    exp_54_ram[1622] = 250;
    exp_54_ram[1623] = 0;
    exp_54_ram[1624] = 252;
    exp_54_ram[1625] = 250;
    exp_54_ram[1626] = 0;
    exp_54_ram[1627] = 187;
    exp_54_ram[1628] = 0;
    exp_54_ram[1629] = 0;
    exp_54_ram[1630] = 250;
    exp_54_ram[1631] = 250;
    exp_54_ram[1632] = 250;
    exp_54_ram[1633] = 0;
    exp_54_ram[1634] = 231;
    exp_54_ram[1635] = 0;
    exp_54_ram[1636] = 0;
    exp_54_ram[1637] = 153;
    exp_54_ram[1638] = 0;
    exp_54_ram[1639] = 173;
    exp_54_ram[1640] = 0;
    exp_54_ram[1641] = 0;
    exp_54_ram[1642] = 0;
    exp_54_ram[1643] = 159;
    exp_54_ram[1644] = 156;
    exp_54_ram[1645] = 82;
    exp_54_ram[1646] = 250;
    exp_54_ram[1647] = 0;
    exp_54_ram[1648] = 208;
    exp_54_ram[1649] = 0;
    exp_54_ram[1650] = 0;
    exp_54_ram[1651] = 227;
    exp_54_ram[1652] = 0;
    exp_54_ram[1653] = 0;
    exp_54_ram[1654] = 156;
    exp_54_ram[1655] = 0;
    exp_54_ram[1656] = 168;
    exp_54_ram[1657] = 0;
    exp_54_ram[1658] = 0;
    exp_54_ram[1659] = 0;
    exp_54_ram[1660] = 159;
    exp_54_ram[1661] = 152;
    exp_54_ram[1662] = 78;
    exp_54_ram[1663] = 250;
    exp_54_ram[1664] = 0;
    exp_54_ram[1665] = 200;
    exp_54_ram[1666] = 0;
    exp_54_ram[1667] = 0;
    exp_54_ram[1668] = 223;
    exp_54_ram[1669] = 0;
    exp_54_ram[1670] = 0;
    exp_54_ram[1671] = 153;
    exp_54_ram[1672] = 0;
    exp_54_ram[1673] = 164;
    exp_54_ram[1674] = 0;
    exp_54_ram[1675] = 0;
    exp_54_ram[1676] = 0;
    exp_54_ram[1677] = 160;
    exp_54_ram[1678] = 148;
    exp_54_ram[1679] = 74;
    exp_54_ram[1680] = 250;
    exp_54_ram[1681] = 0;
    exp_54_ram[1682] = 209;
    exp_54_ram[1683] = 0;
    exp_54_ram[1684] = 0;
    exp_54_ram[1685] = 156;
    exp_54_ram[1686] = 0;
    exp_54_ram[1687] = 161;
    exp_54_ram[1688] = 0;
    exp_54_ram[1689] = 0;
    exp_54_ram[1690] = 0;
    exp_54_ram[1691] = 160;
    exp_54_ram[1692] = 144;
    exp_54_ram[1693] = 70;
    exp_54_ram[1694] = 7;
    exp_54_ram[1695] = 252;
    exp_54_ram[1696] = 0;
    exp_54_ram[1697] = 250;
    exp_54_ram[1698] = 1;
    exp_54_ram[1699] = 250;
    exp_54_ram[1700] = 0;
    exp_54_ram[1701] = 250;
    exp_54_ram[1702] = 1;
    exp_54_ram[1703] = 250;
    exp_54_ram[1704] = 250;
    exp_54_ram[1705] = 252;
    exp_54_ram[1706] = 250;
    exp_54_ram[1707] = 0;
    exp_54_ram[1708] = 167;
    exp_54_ram[1709] = 0;
    exp_54_ram[1710] = 0;
    exp_54_ram[1711] = 250;
    exp_54_ram[1712] = 250;
    exp_54_ram[1713] = 250;
    exp_54_ram[1714] = 0;
    exp_54_ram[1715] = 211;
    exp_54_ram[1716] = 0;
    exp_54_ram[1717] = 0;
    exp_54_ram[1718] = 156;
    exp_54_ram[1719] = 0;
    exp_54_ram[1720] = 152;
    exp_54_ram[1721] = 0;
    exp_54_ram[1722] = 0;
    exp_54_ram[1723] = 0;
    exp_54_ram[1724] = 161;
    exp_54_ram[1725] = 136;
    exp_54_ram[1726] = 62;
    exp_54_ram[1727] = 250;
    exp_54_ram[1728] = 0;
    exp_54_ram[1729] = 188;
    exp_54_ram[1730] = 0;
    exp_54_ram[1731] = 0;
    exp_54_ram[1732] = 207;
    exp_54_ram[1733] = 0;
    exp_54_ram[1734] = 0;
    exp_54_ram[1735] = 161;
    exp_54_ram[1736] = 0;
    exp_54_ram[1737] = 148;
    exp_54_ram[1738] = 0;
    exp_54_ram[1739] = 0;
    exp_54_ram[1740] = 0;
    exp_54_ram[1741] = 163;
    exp_54_ram[1742] = 132;
    exp_54_ram[1743] = 58;
    exp_54_ram[1744] = 250;
    exp_54_ram[1745] = 0;
    exp_54_ram[1746] = 180;
    exp_54_ram[1747] = 0;
    exp_54_ram[1748] = 0;
    exp_54_ram[1749] = 203;
    exp_54_ram[1750] = 0;
    exp_54_ram[1751] = 0;
    exp_54_ram[1752] = 156;
    exp_54_ram[1753] = 0;
    exp_54_ram[1754] = 144;
    exp_54_ram[1755] = 0;
    exp_54_ram[1756] = 0;
    exp_54_ram[1757] = 0;
    exp_54_ram[1758] = 164;
    exp_54_ram[1759] = 128;
    exp_54_ram[1760] = 53;
    exp_54_ram[1761] = 250;
    exp_54_ram[1762] = 0;
    exp_54_ram[1763] = 189;
    exp_54_ram[1764] = 0;
    exp_54_ram[1765] = 0;
    exp_54_ram[1766] = 161;
    exp_54_ram[1767] = 0;
    exp_54_ram[1768] = 140;
    exp_54_ram[1769] = 0;
    exp_54_ram[1770] = 0;
    exp_54_ram[1771] = 0;
    exp_54_ram[1772] = 164;
    exp_54_ram[1773] = 252;
    exp_54_ram[1774] = 50;
    exp_54_ram[1775] = 0;
    exp_54_ram[1776] = 165;
    exp_54_ram[1777] = 251;
    exp_54_ram[1778] = 7;
    exp_54_ram[1779] = 252;
    exp_54_ram[1780] = 0;
    exp_54_ram[1781] = 250;
    exp_54_ram[1782] = 1;
    exp_54_ram[1783] = 250;
    exp_54_ram[1784] = 250;
    exp_54_ram[1785] = 3;
    exp_54_ram[1786] = 250;
    exp_54_ram[1787] = 3;
    exp_54_ram[1788] = 250;
    exp_54_ram[1789] = 255;
    exp_54_ram[1790] = 252;
    exp_54_ram[1791] = 250;
    exp_54_ram[1792] = 0;
    exp_54_ram[1793] = 145;
    exp_54_ram[1794] = 0;
    exp_54_ram[1795] = 0;
    exp_54_ram[1796] = 250;
    exp_54_ram[1797] = 250;
    exp_54_ram[1798] = 250;
    exp_54_ram[1799] = 250;
    exp_54_ram[1800] = 0;
    exp_54_ram[1801] = 0;
    exp_54_ram[1802] = 183;
    exp_54_ram[1803] = 150;
    exp_54_ram[1804] = 252;
    exp_54_ram[1805] = 252;
    exp_54_ram[1806] = 252;
    exp_54_ram[1807] = 13;
    exp_54_ram[1808] = 0;
    exp_54_ram[1809] = 148;
    exp_54_ram[1810] = 0;
    exp_54_ram[1811] = 0;
    exp_54_ram[1812] = 253;
    exp_54_ram[1813] = 253;
    exp_54_ram[1814] = 0;
    exp_54_ram[1815] = 0;
    exp_54_ram[1816] = 149;
    exp_54_ram[1817] = 0;
    exp_54_ram[1818] = 0;
    exp_54_ram[1819] = 0;
    exp_54_ram[1820] = 246;
    exp_54_ram[1821] = 0;
    exp_54_ram[1822] = 146;
    exp_54_ram[1823] = 0;
    exp_54_ram[1824] = 0;
    exp_54_ram[1825] = 0;
    exp_54_ram[1826] = 0;
    exp_54_ram[1827] = 0;
    exp_54_ram[1828] = 0;
    exp_54_ram[1829] = 130;
    exp_54_ram[1830] = 0;
    exp_54_ram[1831] = 250;
    exp_54_ram[1832] = 0;
    exp_54_ram[1833] = 246;
    exp_54_ram[1834] = 0;
    exp_54_ram[1835] = 0;
    exp_54_ram[1836] = 253;
    exp_54_ram[1837] = 253;
    exp_54_ram[1838] = 1;
    exp_54_ram[1839] = 0;
    exp_54_ram[1840] = 0;
    exp_54_ram[1841] = 1;
    exp_54_ram[1842] = 0;
    exp_54_ram[1843] = 0;
    exp_54_ram[1844] = 252;
    exp_54_ram[1845] = 252;
    exp_54_ram[1846] = 0;
    exp_54_ram[1847] = 167;
    exp_54_ram[1848] = 0;
    exp_54_ram[1849] = 0;
    exp_54_ram[1850] = 250;
    exp_54_ram[1851] = 250;
    exp_54_ram[1852] = 250;
    exp_54_ram[1853] = 0;
    exp_54_ram[1854] = 166;
    exp_54_ram[1855] = 0;
    exp_54_ram[1856] = 0;
    exp_54_ram[1857] = 231;
    exp_54_ram[1858] = 253;
    exp_54_ram[1859] = 0;
    exp_54_ram[1860] = 252;
    exp_54_ram[1861] = 253;
    exp_54_ram[1862] = 0;
    exp_54_ram[1863] = 242;
    exp_54_ram[1864] = 7;
    exp_54_ram[1865] = 252;
    exp_54_ram[1866] = 0;
    exp_54_ram[1867] = 250;
    exp_54_ram[1868] = 1;
    exp_54_ram[1869] = 250;
    exp_54_ram[1870] = 0;
    exp_54_ram[1871] = 250;
    exp_54_ram[1872] = 3;
    exp_54_ram[1873] = 250;
    exp_54_ram[1874] = 3;
    exp_54_ram[1875] = 250;
    exp_54_ram[1876] = 0;
    exp_54_ram[1877] = 252;
    exp_54_ram[1878] = 250;
    exp_54_ram[1879] = 0;
    exp_54_ram[1880] = 252;
    exp_54_ram[1881] = 0;
    exp_54_ram[1882] = 0;
    exp_54_ram[1883] = 250;
    exp_54_ram[1884] = 250;
    exp_54_ram[1885] = 250;
    exp_54_ram[1886] = 0;
    exp_54_ram[1887] = 168;
    exp_54_ram[1888] = 0;
    exp_54_ram[1889] = 0;
    exp_54_ram[1890] = 223;
    exp_54_ram[1891] = 250;
    exp_54_ram[1892] = 0;
    exp_54_ram[1893] = 157;
    exp_54_ram[1894] = 0;
    exp_54_ram[1895] = 0;
    exp_54_ram[1896] = 221;
    exp_54_ram[1897] = 250;
    exp_54_ram[1898] = 250;
    exp_54_ram[1899] = 0;
    exp_54_ram[1900] = 0;
    exp_54_ram[1901] = 158;
    exp_54_ram[1902] = 0;
    exp_54_ram[1903] = 153;
    exp_54_ram[1904] = 0;
    exp_54_ram[1905] = 0;
    exp_54_ram[1906] = 250;
    exp_54_ram[1907] = 250;
    exp_54_ram[1908] = 250;
    exp_54_ram[1909] = 0;
    exp_54_ram[1910] = 152;
    exp_54_ram[1911] = 0;
    exp_54_ram[1912] = 0;
    exp_54_ram[1913] = 217;
    exp_54_ram[1914] = 250;
    exp_54_ram[1915] = 252;
    exp_54_ram[1916] = 252;
    exp_54_ram[1917] = 252;
    exp_54_ram[1918] = 13;
    exp_54_ram[1919] = 0;
    exp_54_ram[1920] = 249;
    exp_54_ram[1921] = 0;
    exp_54_ram[1922] = 0;
    exp_54_ram[1923] = 253;
    exp_54_ram[1924] = 253;
    exp_54_ram[1925] = 0;
    exp_54_ram[1926] = 0;
    exp_54_ram[1927] = 249;
    exp_54_ram[1928] = 0;
    exp_54_ram[1929] = 0;
    exp_54_ram[1930] = 0;
    exp_54_ram[1931] = 246;
    exp_54_ram[1932] = 0;
    exp_54_ram[1933] = 247;
    exp_54_ram[1934] = 0;
    exp_54_ram[1935] = 0;
    exp_54_ram[1936] = 0;
    exp_54_ram[1937] = 0;
    exp_54_ram[1938] = 0;
    exp_54_ram[1939] = 0;
    exp_54_ram[1940] = 231;
    exp_54_ram[1941] = 0;
    exp_54_ram[1942] = 250;
    exp_54_ram[1943] = 0;
    exp_54_ram[1944] = 246;
    exp_54_ram[1945] = 0;
    exp_54_ram[1946] = 0;
    exp_54_ram[1947] = 253;
    exp_54_ram[1948] = 253;
    exp_54_ram[1949] = 1;
    exp_54_ram[1950] = 0;
    exp_54_ram[1951] = 0;
    exp_54_ram[1952] = 1;
    exp_54_ram[1953] = 0;
    exp_54_ram[1954] = 0;
    exp_54_ram[1955] = 252;
    exp_54_ram[1956] = 252;
    exp_54_ram[1957] = 0;
    exp_54_ram[1958] = 139;
    exp_54_ram[1959] = 0;
    exp_54_ram[1960] = 0;
    exp_54_ram[1961] = 250;
    exp_54_ram[1962] = 250;
    exp_54_ram[1963] = 250;
    exp_54_ram[1964] = 0;
    exp_54_ram[1965] = 139;
    exp_54_ram[1966] = 0;
    exp_54_ram[1967] = 0;
    exp_54_ram[1968] = 203;
    exp_54_ram[1969] = 253;
    exp_54_ram[1970] = 0;
    exp_54_ram[1971] = 252;
    exp_54_ram[1972] = 253;
    exp_54_ram[1973] = 0;
    exp_54_ram[1974] = 242;
    exp_54_ram[1975] = 5;
    exp_54_ram[1976] = 5;
    exp_54_ram[1977] = 5;
    exp_54_ram[1978] = 5;
    exp_54_ram[1979] = 4;
    exp_54_ram[1980] = 4;
    exp_54_ram[1981] = 4;
    exp_54_ram[1982] = 4;
    exp_54_ram[1983] = 6;
    exp_54_ram[1984] = 0;
    exp_54_ram[1985] = 255;
    exp_54_ram[1986] = 0;
    exp_54_ram[1987] = 0;
    exp_54_ram[1988] = 1;
    exp_54_ram[1989] = 138;
    exp_54_ram[1990] = 134;
    exp_54_ram[1991] = 0;
    exp_54_ram[1992] = 0;
    exp_54_ram[1993] = 0;
    exp_54_ram[1994] = 1;
    exp_54_ram[1995] = 0;
    exp_54_ram[1996] = 0;
    exp_54_ram[1997] = 0;
    exp_54_ram[1998] = 2;
    exp_54_ram[1999] = 255;
    exp_54_ram[2000] = 2;
    exp_54_ram[2001] = 0;
    exp_54_ram[2002] = 0;
    exp_54_ram[2003] = 0;
    exp_54_ram[2004] = 64;
    exp_54_ram[2005] = 1;
    exp_54_ram[2006] = 0;
    exp_54_ram[2007] = 254;
    exp_54_ram[2008] = 255;
    exp_54_ram[2009] = 0;
    exp_54_ram[2010] = 254;
    exp_54_ram[2011] = 2;
    exp_54_ram[2012] = 128;
    exp_54_ram[2013] = 77;
    exp_54_ram[2014] = 117;
    exp_54_ram[2015] = 100;
    exp_54_ram[2016] = 70;
    exp_54_ram[2017] = 97;
    exp_54_ram[2018] = 0;
    exp_54_ram[2019] = 70;
    exp_54_ram[2020] = 97;
    exp_54_ram[2021] = 114;
    exp_54_ram[2022] = 74;
    exp_54_ram[2023] = 117;
    exp_54_ram[2024] = 103;
    exp_54_ram[2025] = 79;
    exp_54_ram[2026] = 111;
    exp_54_ram[2027] = 99;
    exp_54_ram[2028] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_52) begin
      exp_54_ram[exp_48] <= exp_50;
    end
  end
  assign exp_54 = exp_54_ram[exp_49];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_80) begin
        exp_54_ram[exp_76] <= exp_78;
    end
  end
  assign exp_82 = exp_54_ram[exp_77];
  assign exp_53 = exp_121;
  assign exp_121 = 1;
  assign exp_49 = exp_120;
  assign exp_120 = exp_10[31:2];
  assign exp_10 = exp_1;
  assign exp_52 = exp_116;
  assign exp_116 = exp_114 & exp_115;
  assign exp_114 = exp_14 & exp_15;
  assign exp_115 = exp_16[3:3];
  assign exp_16 = exp_7;
  assign exp_7 = exp_252;
  assign exp_252 = exp_533;

  reg [3:0] exp_533_reg;
  always@(*) begin
    case (exp_385)
      0:exp_533_reg <= exp_520;
      1:exp_533_reg <= exp_525;
      2:exp_533_reg <= exp_526;
      3:exp_533_reg <= exp_527;
      4:exp_533_reg <= exp_528;
      5:exp_533_reg <= exp_529;
      6:exp_533_reg <= exp_530;
      7:exp_533_reg <= exp_531;
      default:exp_533_reg <= exp_532;
    endcase
  end
  assign exp_533 = exp_533_reg;
  assign exp_532 = 0;
  assign exp_520 = exp_516 << exp_519;
  assign exp_516 = 1;
  assign exp_519 = exp_518 + exp_517;
  assign exp_518 = 0;
  assign exp_517 = exp_453[1:0];
  assign exp_525 = exp_521 << exp_524;
  assign exp_521 = 3;
  assign exp_524 = exp_523 + exp_522;
  assign exp_523 = 0;
  assign exp_522 = exp_453[1:1];
  assign exp_526 = 15;
  assign exp_527 = 0;
  assign exp_528 = 0;
  assign exp_529 = 0;
  assign exp_530 = 0;
  assign exp_531 = 0;
  assign exp_48 = exp_112;
  assign exp_112 = exp_10[31:2];
  assign exp_50 = exp_113;
  assign exp_113 = exp_11[31:24];
  assign exp_11 = exp_2;
  assign exp_2 = exp_247;
  assign exp_247 = exp_515;

  reg [31:0] exp_515_reg;
  always@(*) begin
    case (exp_385)
      0:exp_515_reg <= exp_502;
      1:exp_515_reg <= exp_506;
      2:exp_515_reg <= exp_508;
      3:exp_515_reg <= exp_509;
      4:exp_515_reg <= exp_510;
      5:exp_515_reg <= exp_511;
      6:exp_515_reg <= exp_512;
      7:exp_515_reg <= exp_513;
      default:exp_515_reg <= exp_514;
    endcase
  end
  assign exp_515 = exp_515_reg;
  assign exp_514 = 0;

  reg [31:0] exp_502_reg;
  always@(*) begin
    case (exp_456)
      0:exp_502_reg <= exp_488;
      1:exp_502_reg <= exp_496;
      2:exp_502_reg <= exp_498;
      3:exp_502_reg <= exp_500;
      default:exp_502_reg <= exp_501;
    endcase
  end
  assign exp_502 = exp_502_reg;
  assign exp_501 = 0;
  assign exp_488 = exp_487;
  assign exp_487 = exp_486 + exp_485;
  assign exp_486 = 0;
  assign exp_485 = exp_375[7:0];

      reg [31:0] exp_375_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_375_reg <= exp_318;
        end
      end
      assign exp_375 = exp_375_reg;
      assign exp_496 = exp_488 << exp_495;
  assign exp_495 = 8;
  assign exp_498 = exp_488 << exp_497;
  assign exp_497 = 16;
  assign exp_500 = exp_488 << exp_499;
  assign exp_499 = 24;

  reg [31:0] exp_506_reg;
  always@(*) begin
    case (exp_459)
      0:exp_506_reg <= exp_492;
      1:exp_506_reg <= exp_504;
      default:exp_506_reg <= exp_505;
    endcase
  end
  assign exp_506 = exp_506_reg;
  assign exp_459 = exp_458 + exp_457;
  assign exp_458 = 0;
  assign exp_457 = exp_453[1:1];
  assign exp_505 = 0;
  assign exp_492 = exp_491;
  assign exp_491 = exp_490 + exp_489;
  assign exp_490 = 0;
  assign exp_489 = exp_375[15:0];
  assign exp_504 = exp_492 << exp_503;
  assign exp_503 = 16;
  assign exp_508 = exp_507 + exp_494;
  assign exp_507 = 0;
  assign exp_494 = exp_493 + exp_375;
  assign exp_493 = 0;
  assign exp_509 = 0;
  assign exp_510 = 0;
  assign exp_511 = 0;
  assign exp_512 = 0;
  assign exp_513 = 0;

  //Create RAM
  reg [7:0] exp_47_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_47_ram[0] = 0;
    exp_47_ram[1] = 0;
    exp_47_ram[2] = 0;
    exp_47_ram[3] = 0;
    exp_47_ram[4] = 0;
    exp_47_ram[5] = 0;
    exp_47_ram[6] = 0;
    exp_47_ram[7] = 0;
    exp_47_ram[8] = 0;
    exp_47_ram[9] = 0;
    exp_47_ram[10] = 0;
    exp_47_ram[11] = 0;
    exp_47_ram[12] = 0;
    exp_47_ram[13] = 0;
    exp_47_ram[14] = 0;
    exp_47_ram[15] = 0;
    exp_47_ram[16] = 0;
    exp_47_ram[17] = 0;
    exp_47_ram[18] = 0;
    exp_47_ram[19] = 0;
    exp_47_ram[20] = 0;
    exp_47_ram[21] = 0;
    exp_47_ram[22] = 0;
    exp_47_ram[23] = 0;
    exp_47_ram[24] = 0;
    exp_47_ram[25] = 0;
    exp_47_ram[26] = 0;
    exp_47_ram[27] = 0;
    exp_47_ram[28] = 0;
    exp_47_ram[29] = 0;
    exp_47_ram[30] = 0;
    exp_47_ram[31] = 0;
    exp_47_ram[32] = 193;
    exp_47_ram[33] = 16;
    exp_47_ram[34] = 0;
    exp_47_ram[35] = 5;
    exp_47_ram[36] = 5;
    exp_47_ram[37] = 6;
    exp_47_ram[38] = 6;
    exp_47_ram[39] = 8;
    exp_47_ram[40] = 6;
    exp_47_ram[41] = 0;
    exp_47_ram[42] = 134;
    exp_47_ram[43] = 197;
    exp_47_ram[44] = 1;
    exp_47_ram[45] = 230;
    exp_47_ram[46] = 240;
    exp_47_ram[47] = 199;
    exp_47_ram[48] = 55;
    exp_47_ram[49] = 230;
    exp_47_ram[50] = 166;
    exp_47_ram[51] = 6;
    exp_47_ram[52] = 0;
    exp_47_ram[53] = 230;
    exp_47_ram[54] = 229;
    exp_47_ram[55] = 229;
    exp_47_ram[56] = 215;
    exp_47_ram[57] = 232;
    exp_47_ram[58] = 214;
    exp_47_ram[59] = 183;
    exp_47_ram[60] = 216;
    exp_47_ram[61] = 8;
    exp_47_ram[62] = 21;
    exp_47_ram[63] = 8;
    exp_47_ram[64] = 6;
    exp_47_ram[65] = 3;
    exp_47_ram[66] = 21;
    exp_47_ram[67] = 6;
    exp_47_ram[68] = 214;
    exp_47_ram[69] = 7;
    exp_47_ram[70] = 247;
    exp_47_ram[71] = 183;
    exp_47_ram[72] = 7;
    exp_47_ram[73] = 246;
    exp_47_ram[74] = 7;
    exp_47_ram[75] = 183;
    exp_47_ram[76] = 230;
    exp_47_ram[77] = 7;
    exp_47_ram[78] = 183;
    exp_47_ram[79] = 23;
    exp_47_ram[80] = 3;
    exp_47_ram[81] = 3;
    exp_47_ram[82] = 23;
    exp_47_ram[83] = 7;
    exp_47_ram[84] = 103;
    exp_47_ram[85] = 246;
    exp_47_ram[86] = 7;
    exp_47_ram[87] = 211;
    exp_47_ram[88] = 104;
    exp_47_ram[89] = 247;
    exp_47_ram[90] = 3;
    exp_47_ram[91] = 211;
    exp_47_ram[92] = 231;
    exp_47_ram[93] = 5;
    exp_47_ram[94] = 197;
    exp_47_ram[95] = 0;
    exp_47_ram[96] = 64;
    exp_47_ram[97] = 0;
    exp_47_ram[98] = 0;
    exp_47_ram[99] = 166;
    exp_47_ram[100] = 128;
    exp_47_ram[101] = 31;
    exp_47_ram[102] = 6;
    exp_47_ram[103] = 16;
    exp_47_ram[104] = 199;
    exp_47_ram[105] = 1;
    exp_47_ram[106] = 232;
    exp_47_ram[107] = 240;
    exp_47_ram[108] = 7;
    exp_47_ram[109] = 128;
    exp_47_ram[110] = 168;
    exp_47_ram[111] = 230;
    exp_47_ram[112] = 6;
    exp_47_ram[113] = 0;
    exp_47_ram[114] = 167;
    exp_47_ram[115] = 230;
    exp_47_ram[116] = 230;
    exp_47_ram[117] = 7;
    exp_47_ram[118] = 16;
    exp_47_ram[119] = 8;
    exp_47_ram[120] = 8;
    exp_47_ram[121] = 6;
    exp_47_ram[122] = 3;
    exp_47_ram[123] = 23;
    exp_47_ram[124] = 23;
    exp_47_ram[125] = 6;
    exp_47_ram[126] = 230;
    exp_47_ram[127] = 246;
    exp_47_ram[128] = 7;
    exp_47_ram[129] = 199;
    exp_47_ram[130] = 7;
    exp_47_ram[131] = 247;
    exp_47_ram[132] = 7;
    exp_47_ram[133] = 199;
    exp_47_ram[134] = 231;
    exp_47_ram[135] = 7;
    exp_47_ram[136] = 199;
    exp_47_ram[137] = 23;
    exp_47_ram[138] = 3;
    exp_47_ram[139] = 3;
    exp_47_ram[140] = 23;
    exp_47_ram[141] = 7;
    exp_47_ram[142] = 103;
    exp_47_ram[143] = 230;
    exp_47_ram[144] = 7;
    exp_47_ram[145] = 211;
    exp_47_ram[146] = 104;
    exp_47_ram[147] = 247;
    exp_47_ram[148] = 3;
    exp_47_ram[149] = 211;
    exp_47_ram[150] = 231;
    exp_47_ram[151] = 5;
    exp_47_ram[152] = 197;
    exp_47_ram[153] = 0;
    exp_47_ram[154] = 0;
    exp_47_ram[155] = 0;
    exp_47_ram[156] = 232;
    exp_47_ram[157] = 128;
    exp_47_ram[158] = 31;
    exp_47_ram[159] = 216;
    exp_47_ram[160] = 231;
    exp_47_ram[161] = 216;
    exp_47_ram[162] = 215;
    exp_47_ram[163] = 232;
    exp_47_ram[164] = 8;
    exp_47_ram[165] = 247;
    exp_47_ram[166] = 21;
    exp_47_ram[167] = 8;
    exp_47_ram[168] = 7;
    exp_47_ram[169] = 6;
    exp_47_ram[170] = 21;
    exp_47_ram[171] = 7;
    exp_47_ram[172] = 183;
    exp_47_ram[173] = 167;
    exp_47_ram[174] = 5;
    exp_47_ram[175] = 215;
    exp_47_ram[176] = 7;
    exp_47_ram[177] = 245;
    exp_47_ram[178] = 7;
    exp_47_ram[179] = 215;
    exp_47_ram[180] = 229;
    exp_47_ram[181] = 7;
    exp_47_ram[182] = 215;
    exp_47_ram[183] = 22;
    exp_47_ram[184] = 6;
    exp_47_ram[185] = 6;
    exp_47_ram[186] = 22;
    exp_47_ram[187] = 7;
    exp_47_ram[188] = 215;
    exp_47_ram[189] = 199;
    exp_47_ram[190] = 6;
    exp_47_ram[191] = 167;
    exp_47_ram[192] = 7;
    exp_47_ram[193] = 246;
    exp_47_ram[194] = 7;
    exp_47_ram[195] = 167;
    exp_47_ram[196] = 230;
    exp_47_ram[197] = 7;
    exp_47_ram[198] = 5;
    exp_47_ram[199] = 167;
    exp_47_ram[200] = 229;
    exp_47_ram[201] = 159;
    exp_47_ram[202] = 213;
    exp_47_ram[203] = 1;
    exp_47_ram[204] = 230;
    exp_47_ram[205] = 240;
    exp_47_ram[206] = 215;
    exp_47_ram[207] = 53;
    exp_47_ram[208] = 0;
    exp_47_ram[209] = 182;
    exp_47_ram[210] = 135;
    exp_47_ram[211] = 167;
    exp_47_ram[212] = 7;
    exp_47_ram[213] = 0;
    exp_47_ram[214] = 183;
    exp_47_ram[215] = 229;
    exp_47_ram[216] = 229;
    exp_47_ram[217] = 16;
    exp_47_ram[218] = 246;
    exp_47_ram[219] = 200;
    exp_47_ram[220] = 21;
    exp_47_ram[221] = 31;
    exp_47_ram[222] = 0;
    exp_47_ram[223] = 0;
    exp_47_ram[224] = 230;
    exp_47_ram[225] = 128;
    exp_47_ram[226] = 159;
    exp_47_ram[227] = 230;
    exp_47_ram[228] = 182;
    exp_47_ram[229] = 216;
    exp_47_ram[230] = 231;
    exp_47_ram[231] = 8;
    exp_47_ram[232] = 222;
    exp_47_ram[233] = 183;
    exp_47_ram[234] = 232;
    exp_47_ram[235] = 182;
    exp_47_ram[236] = 247;
    exp_47_ram[237] = 8;
    exp_47_ram[238] = 7;
    exp_47_ram[239] = 6;
    exp_47_ram[240] = 222;
    exp_47_ram[241] = 6;
    exp_47_ram[242] = 230;
    exp_47_ram[243] = 199;
    exp_47_ram[244] = 14;
    exp_47_ram[245] = 231;
    exp_47_ram[246] = 7;
    exp_47_ram[247] = 254;
    exp_47_ram[248] = 7;
    exp_47_ram[249] = 231;
    exp_47_ram[250] = 238;
    exp_47_ram[251] = 7;
    exp_47_ram[252] = 231;
    exp_47_ram[253] = 215;
    exp_47_ram[254] = 215;
    exp_47_ram[255] = 6;
    exp_47_ram[256] = 231;
    exp_47_ram[257] = 6;
    exp_47_ram[258] = 7;
    exp_47_ram[259] = 246;
    exp_47_ram[260] = 7;
    exp_47_ram[261] = 199;
    exp_47_ram[262] = 7;
    exp_47_ram[263] = 247;
    exp_47_ram[264] = 7;
    exp_47_ram[265] = 199;
    exp_47_ram[266] = 231;
    exp_47_ram[267] = 7;
    exp_47_ram[268] = 5;
    exp_47_ram[269] = 1;
    exp_47_ram[270] = 197;
    exp_47_ram[271] = 254;
    exp_47_ram[272] = 213;
    exp_47_ram[273] = 5;
    exp_47_ram[274] = 211;
    exp_47_ram[275] = 3;
    exp_47_ram[276] = 199;
    exp_47_ram[277] = 216;
    exp_47_ram[278] = 214;
    exp_47_ram[279] = 14;
    exp_47_ram[280] = 104;
    exp_47_ram[281] = 216;
    exp_47_ram[282] = 7;
    exp_47_ram[283] = 102;
    exp_47_ram[284] = 215;
    exp_47_ram[285] = 214;
    exp_47_ram[286] = 7;
    exp_47_ram[287] = 198;
    exp_47_ram[288] = 199;
    exp_47_ram[289] = 199;
    exp_47_ram[290] = 1;
    exp_47_ram[291] = 247;
    exp_47_ram[292] = 247;
    exp_47_ram[293] = 7;
    exp_47_ram[294] = 254;
    exp_47_ram[295] = 184;
    exp_47_ram[296] = 199;
    exp_47_ram[297] = 0;
    exp_47_ram[298] = 232;
    exp_47_ram[299] = 245;
    exp_47_ram[300] = 223;
    exp_47_ram[301] = 0;
    exp_47_ram[302] = 0;
    exp_47_ram[303] = 159;
    exp_47_ram[304] = 16;
    exp_47_ram[305] = 247;
    exp_47_ram[306] = 69;
    exp_47_ram[307] = 183;
    exp_47_ram[308] = 5;
    exp_47_ram[309] = 5;
    exp_47_ram[310] = 248;
    exp_47_ram[311] = 245;
    exp_47_ram[312] = 240;
    exp_47_ram[313] = 70;
    exp_47_ram[314] = 215;
    exp_47_ram[315] = 6;
    exp_47_ram[316] = 245;
    exp_47_ram[317] = 246;
    exp_47_ram[318] = 216;
    exp_47_ram[319] = 248;
    exp_47_ram[320] = 14;
    exp_47_ram[321] = 32;
    exp_47_ram[322] = 0;
    exp_47_ram[323] = 213;
    exp_47_ram[324] = 199;
    exp_47_ram[325] = 14;
    exp_47_ram[326] = 8;
    exp_47_ram[327] = 248;
    exp_47_ram[328] = 23;
    exp_47_ram[329] = 5;
    exp_47_ram[330] = 199;
    exp_47_ram[331] = 6;
    exp_47_ram[332] = 7;
    exp_47_ram[333] = 213;
    exp_47_ram[334] = 5;
    exp_47_ram[335] = 5;
    exp_47_ram[336] = 240;
    exp_47_ram[337] = 0;
    exp_47_ram[338] = 240;
    exp_47_ram[339] = 6;
    exp_47_ram[340] = 6;
    exp_47_ram[341] = 0;
    exp_47_ram[342] = 184;
    exp_47_ram[343] = 5;
    exp_47_ram[344] = 0;
    exp_47_ram[345] = 23;
    exp_47_ram[346] = 232;
    exp_47_ram[347] = 110;
    exp_47_ram[348] = 195;
    exp_47_ram[349] = 0;
    exp_47_ram[350] = 0;
    exp_47_ram[351] = 16;
    exp_47_ram[352] = 0;
    exp_47_ram[353] = 7;
    exp_47_ram[354] = 95;
    exp_47_ram[355] = 232;
    exp_47_ram[356] = 95;
    exp_47_ram[357] = 5;
    exp_47_ram[358] = 5;
    exp_47_ram[359] = 0;
    exp_47_ram[360] = 159;
    exp_47_ram[361] = 1;
    exp_47_ram[362] = 129;
    exp_47_ram[363] = 17;
    exp_47_ram[364] = 5;
    exp_47_ram[365] = 5;
    exp_47_ram[366] = 192;
    exp_47_ram[367] = 224;
    exp_47_ram[368] = 160;
    exp_47_ram[369] = 167;
    exp_47_ram[370] = 167;
    exp_47_ram[371] = 176;
    exp_47_ram[372] = 167;
    exp_47_ram[373] = 85;
    exp_47_ram[374] = 244;
    exp_47_ram[375] = 164;
    exp_47_ram[376] = 193;
    exp_47_ram[377] = 4;
    exp_47_ram[378] = 199;
    exp_47_ram[379] = 129;
    exp_47_ram[380] = 71;
    exp_47_ram[381] = 199;
    exp_47_ram[382] = 247;
    exp_47_ram[383] = 6;
    exp_47_ram[384] = 1;
    exp_47_ram[385] = 0;
    exp_47_ram[386] = 85;
    exp_47_ram[387] = 244;
    exp_47_ram[388] = 0;
    exp_47_ram[389] = 223;
    exp_47_ram[390] = 0;
    exp_47_ram[391] = 0;
    exp_47_ram[392] = 31;
    exp_47_ram[393] = 1;
    exp_47_ram[394] = 17;
    exp_47_ram[395] = 129;
    exp_47_ram[396] = 145;
    exp_47_ram[397] = 33;
    exp_47_ram[398] = 49;
    exp_47_ram[399] = 65;
    exp_47_ram[400] = 181;
    exp_47_ram[401] = 7;
    exp_47_ram[402] = 5;
    exp_47_ram[403] = 5;
    exp_47_ram[404] = 5;
    exp_47_ram[405] = 5;
    exp_47_ram[406] = 5;
    exp_47_ram[407] = 128;
    exp_47_ram[408] = 5;
    exp_47_ram[409] = 224;
    exp_47_ram[410] = 58;
    exp_47_ram[411] = 48;
    exp_47_ram[412] = 71;
    exp_47_ram[413] = 176;
    exp_47_ram[414] = 4;
    exp_47_ram[415] = 55;
    exp_47_ram[416] = 160;
    exp_47_ram[417] = 55;
    exp_47_ram[418] = 176;
    exp_47_ram[419] = 89;
    exp_47_ram[420] = 52;
    exp_47_ram[421] = 148;
    exp_47_ram[422] = 233;
    exp_47_ram[423] = 180;
    exp_47_ram[424] = 228;
    exp_47_ram[425] = 193;
    exp_47_ram[426] = 129;
    exp_47_ram[427] = 196;
    exp_47_ram[428] = 74;
    exp_47_ram[429] = 197;
    exp_47_ram[430] = 186;
    exp_47_ram[431] = 65;
    exp_47_ram[432] = 1;
    exp_47_ram[433] = 193;
    exp_47_ram[434] = 129;
    exp_47_ram[435] = 7;
    exp_47_ram[436] = 7;
    exp_47_ram[437] = 1;
    exp_47_ram[438] = 0;
    exp_47_ram[439] = 128;
    exp_47_ram[440] = 5;
    exp_47_ram[441] = 31;
    exp_47_ram[442] = 89;
    exp_47_ram[443] = 180;
    exp_47_ram[444] = 0;
    exp_47_ram[445] = 31;
    exp_47_ram[446] = 96;
    exp_47_ram[447] = 71;
    exp_47_ram[448] = 137;
    exp_47_ram[449] = 4;
    exp_47_ram[450] = 9;
    exp_47_ram[451] = 0;
    exp_47_ram[452] = 181;
    exp_47_ram[453] = 128;
    exp_47_ram[454] = 160;
    exp_47_ram[455] = 9;
    exp_47_ram[456] = 4;
    exp_47_ram[457] = 54;
    exp_47_ram[458] = 192;
    exp_47_ram[459] = 164;
    exp_47_ram[460] = 5;
    exp_47_ram[461] = 128;
    exp_47_ram[462] = 4;
    exp_47_ram[463] = 9;
    exp_47_ram[464] = 55;
    exp_47_ram[465] = 112;
    exp_47_ram[466] = 55;
    exp_47_ram[467] = 137;
    exp_47_ram[468] = 233;
    exp_47_ram[469] = 128;
    exp_47_ram[470] = 57;
    exp_47_ram[471] = 36;
    exp_47_ram[472] = 185;
    exp_47_ram[473] = 228;
    exp_47_ram[474] = 128;
    exp_47_ram[475] = 247;
    exp_47_ram[476] = 229;
    exp_47_ram[477] = 119;
    exp_47_ram[478] = 7;
    exp_47_ram[479] = 247;
    exp_47_ram[480] = 64;
    exp_47_ram[481] = 215;
    exp_47_ram[482] = 71;
    exp_47_ram[483] = 247;
    exp_47_ram[484] = 245;
    exp_47_ram[485] = 7;
    exp_47_ram[486] = 128;
    exp_47_ram[487] = 229;
    exp_47_ram[488] = 7;
    exp_47_ram[489] = 128;
    exp_47_ram[490] = 247;
    exp_47_ram[491] = 240;
    exp_47_ram[492] = 229;
    exp_47_ram[493] = 58;
    exp_47_ram[494] = 55;
    exp_47_ram[495] = 213;
    exp_47_ram[496] = 245;
    exp_47_ram[497] = 53;
    exp_47_ram[498] = 223;
    exp_47_ram[499] = 137;
    exp_47_ram[500] = 180;
    exp_47_ram[501] = 0;
    exp_47_ram[502] = 31;
    exp_47_ram[503] = 0;
    exp_47_ram[504] = 0;
    exp_47_ram[505] = 0;
    exp_47_ram[506] = 223;
    exp_47_ram[507] = 5;
    exp_47_ram[508] = 0;
    exp_47_ram[509] = 21;
    exp_47_ram[510] = 6;
    exp_47_ram[511] = 197;
    exp_47_ram[512] = 21;
    exp_47_ram[513] = 22;
    exp_47_ram[514] = 5;
    exp_47_ram[515] = 0;
    exp_47_ram[516] = 5;
    exp_47_ram[517] = 5;
    exp_47_ram[518] = 5;
    exp_47_ram[519] = 5;
    exp_47_ram[520] = 240;
    exp_47_ram[521] = 6;
    exp_47_ram[522] = 16;
    exp_47_ram[523] = 182;
    exp_47_ram[524] = 192;
    exp_47_ram[525] = 22;
    exp_47_ram[526] = 22;
    exp_47_ram[527] = 182;
    exp_47_ram[528] = 0;
    exp_47_ram[529] = 197;
    exp_47_ram[530] = 197;
    exp_47_ram[531] = 213;
    exp_47_ram[532] = 22;
    exp_47_ram[533] = 22;
    exp_47_ram[534] = 6;
    exp_47_ram[535] = 0;
    exp_47_ram[536] = 0;
    exp_47_ram[537] = 95;
    exp_47_ram[538] = 5;
    exp_47_ram[539] = 2;
    exp_47_ram[540] = 160;
    exp_47_ram[541] = 176;
    exp_47_ram[542] = 176;
    exp_47_ram[543] = 223;
    exp_47_ram[544] = 176;
    exp_47_ram[545] = 0;
    exp_47_ram[546] = 31;
    exp_47_ram[547] = 160;
    exp_47_ram[548] = 2;
    exp_47_ram[549] = 0;
    exp_47_ram[550] = 5;
    exp_47_ram[551] = 5;
    exp_47_ram[552] = 159;
    exp_47_ram[553] = 5;
    exp_47_ram[554] = 2;
    exp_47_ram[555] = 176;
    exp_47_ram[556] = 5;
    exp_47_ram[557] = 160;
    exp_47_ram[558] = 31;
    exp_47_ram[559] = 176;
    exp_47_ram[560] = 2;
    exp_47_ram[561] = 6;
    exp_47_ram[562] = 0;
    exp_47_ram[563] = 199;
    exp_47_ram[564] = 240;
    exp_47_ram[565] = 6;
    exp_47_ram[566] = 0;
    exp_47_ram[567] = 165;
    exp_47_ram[568] = 7;
    exp_47_ram[569] = 0;
    exp_47_ram[570] = 197;
    exp_47_ram[571] = 197;
    exp_47_ram[572] = 245;
    exp_47_ram[573] = 181;
    exp_47_ram[574] = 159;
    exp_47_ram[575] = 6;
    exp_47_ram[576] = 0;
    exp_47_ram[577] = 199;
    exp_47_ram[578] = 240;
    exp_47_ram[579] = 6;
    exp_47_ram[580] = 0;
    exp_47_ram[581] = 181;
    exp_47_ram[582] = 7;
    exp_47_ram[583] = 0;
    exp_47_ram[584] = 197;
    exp_47_ram[585] = 197;
    exp_47_ram[586] = 245;
    exp_47_ram[587] = 165;
    exp_47_ram[588] = 159;
    exp_47_ram[589] = 1;
    exp_47_ram[590] = 245;
    exp_47_ram[591] = 240;
    exp_47_ram[592] = 167;
    exp_47_ram[593] = 55;
    exp_47_ram[594] = 0;
    exp_47_ram[595] = 0;
    exp_47_ram[596] = 246;
    exp_47_ram[597] = 245;
    exp_47_ram[598] = 135;
    exp_47_ram[599] = 167;
    exp_47_ram[600] = 5;
    exp_47_ram[601] = 166;
    exp_47_ram[602] = 0;
    exp_47_ram[603] = 0;
    exp_47_ram[604] = 0;
    exp_47_ram[605] = 229;
    exp_47_ram[606] = 128;
    exp_47_ram[607] = 223;
    exp_47_ram[608] = 114;
    exp_47_ram[609] = 46;
    exp_47_ram[610] = 0;
    exp_47_ram[611] = 115;
    exp_47_ram[612] = 0;
    exp_47_ram[613] = 109;
    exp_47_ram[614] = 46;
    exp_47_ram[615] = 117;
    exp_47_ram[616] = 112;
    exp_47_ram[617] = 32;
    exp_47_ram[618] = 50;
    exp_47_ram[619] = 48;
    exp_47_ram[620] = 50;
    exp_47_ram[621] = 0;
    exp_47_ram[622] = 102;
    exp_47_ram[623] = 0;
    exp_47_ram[624] = 117;
    exp_47_ram[625] = 112;
    exp_47_ram[626] = 32;
    exp_47_ram[627] = 50;
    exp_47_ram[628] = 48;
    exp_47_ram[629] = 50;
    exp_47_ram[630] = 0;
    exp_47_ram[631] = 102;
    exp_47_ram[632] = 0;
    exp_47_ram[633] = 102;
    exp_47_ram[634] = 0;
    exp_47_ram[635] = 102;
    exp_47_ram[636] = 0;
    exp_47_ram[637] = 102;
    exp_47_ram[638] = 0;
    exp_47_ram[639] = 102;
    exp_47_ram[640] = 0;
    exp_47_ram[641] = 102;
    exp_47_ram[642] = 0;
    exp_47_ram[643] = 102;
    exp_47_ram[644] = 0;
    exp_47_ram[645] = 102;
    exp_47_ram[646] = 0;
    exp_47_ram[647] = 117;
    exp_47_ram[648] = 112;
    exp_47_ram[649] = 32;
    exp_47_ram[650] = 50;
    exp_47_ram[651] = 48;
    exp_47_ram[652] = 50;
    exp_47_ram[653] = 0;
    exp_47_ram[654] = 32;
    exp_47_ram[655] = 108;
    exp_47_ram[656] = 32;
    exp_47_ram[657] = 108;
    exp_47_ram[658] = 32;
    exp_47_ram[659] = 108;
    exp_47_ram[660] = 115;
    exp_47_ram[661] = 0;
    exp_47_ram[662] = 2;
    exp_47_ram[663] = 3;
    exp_47_ram[664] = 4;
    exp_47_ram[665] = 4;
    exp_47_ram[666] = 5;
    exp_47_ram[667] = 5;
    exp_47_ram[668] = 5;
    exp_47_ram[669] = 5;
    exp_47_ram[670] = 6;
    exp_47_ram[671] = 6;
    exp_47_ram[672] = 6;
    exp_47_ram[673] = 6;
    exp_47_ram[674] = 6;
    exp_47_ram[675] = 6;
    exp_47_ram[676] = 6;
    exp_47_ram[677] = 6;
    exp_47_ram[678] = 7;
    exp_47_ram[679] = 7;
    exp_47_ram[680] = 7;
    exp_47_ram[681] = 7;
    exp_47_ram[682] = 7;
    exp_47_ram[683] = 7;
    exp_47_ram[684] = 7;
    exp_47_ram[685] = 7;
    exp_47_ram[686] = 7;
    exp_47_ram[687] = 7;
    exp_47_ram[688] = 7;
    exp_47_ram[689] = 7;
    exp_47_ram[690] = 7;
    exp_47_ram[691] = 7;
    exp_47_ram[692] = 7;
    exp_47_ram[693] = 7;
    exp_47_ram[694] = 8;
    exp_47_ram[695] = 8;
    exp_47_ram[696] = 8;
    exp_47_ram[697] = 8;
    exp_47_ram[698] = 8;
    exp_47_ram[699] = 8;
    exp_47_ram[700] = 8;
    exp_47_ram[701] = 8;
    exp_47_ram[702] = 8;
    exp_47_ram[703] = 8;
    exp_47_ram[704] = 8;
    exp_47_ram[705] = 8;
    exp_47_ram[706] = 8;
    exp_47_ram[707] = 8;
    exp_47_ram[708] = 8;
    exp_47_ram[709] = 8;
    exp_47_ram[710] = 8;
    exp_47_ram[711] = 8;
    exp_47_ram[712] = 8;
    exp_47_ram[713] = 8;
    exp_47_ram[714] = 8;
    exp_47_ram[715] = 8;
    exp_47_ram[716] = 8;
    exp_47_ram[717] = 8;
    exp_47_ram[718] = 8;
    exp_47_ram[719] = 8;
    exp_47_ram[720] = 8;
    exp_47_ram[721] = 8;
    exp_47_ram[722] = 8;
    exp_47_ram[723] = 8;
    exp_47_ram[724] = 8;
    exp_47_ram[725] = 8;
    exp_47_ram[726] = 5;
    exp_47_ram[727] = 0;
    exp_47_ram[728] = 167;
    exp_47_ram[729] = 7;
    exp_47_ram[730] = 7;
    exp_47_ram[731] = 0;
    exp_47_ram[732] = 21;
    exp_47_ram[733] = 229;
    exp_47_ram[734] = 159;
    exp_47_ram[735] = 1;
    exp_47_ram[736] = 0;
    exp_47_ram[737] = 129;
    exp_47_ram[738] = 7;
    exp_47_ram[739] = 17;
    exp_47_ram[740] = 4;
    exp_47_ram[741] = 95;
    exp_47_ram[742] = 160;
    exp_47_ram[743] = 193;
    exp_47_ram[744] = 244;
    exp_47_ram[745] = 129;
    exp_47_ram[746] = 0;
    exp_47_ram[747] = 1;
    exp_47_ram[748] = 0;
    exp_47_ram[749] = 181;
    exp_47_ram[750] = 55;
    exp_47_ram[751] = 5;
    exp_47_ram[752] = 7;
    exp_47_ram[753] = 5;
    exp_47_ram[754] = 197;
    exp_47_ram[755] = 240;
    exp_47_ram[756] = 192;
    exp_47_ram[757] = 7;
    exp_47_ram[758] = 7;
    exp_47_ram[759] = 6;
    exp_47_ram[760] = 22;
    exp_47_ram[761] = 71;
    exp_47_ram[762] = 22;
    exp_47_ram[763] = 135;
    exp_47_ram[764] = 22;
    exp_47_ram[765] = 199;
    exp_47_ram[766] = 22;
    exp_47_ram[767] = 227;
    exp_47_ram[768] = 24;
    exp_47_ram[769] = 246;
    exp_47_ram[770] = 6;
    exp_47_ram[771] = 197;
    exp_47_ram[772] = 197;
    exp_47_ram[773] = 48;
    exp_47_ram[774] = 247;
    exp_47_ram[775] = 6;
    exp_47_ram[776] = 55;
    exp_47_ram[777] = 199;
    exp_47_ram[778] = 230;
    exp_47_ram[779] = 229;
    exp_47_ram[780] = 0;
    exp_47_ram[781] = 246;
    exp_47_ram[782] = 0;
    exp_47_ram[783] = 245;
    exp_47_ram[784] = 8;
    exp_47_ram[785] = 246;
    exp_47_ram[786] = 71;
    exp_47_ram[787] = 24;
    exp_47_ram[788] = 159;
    exp_47_ram[789] = 245;
    exp_47_ram[790] = 7;
    exp_47_ram[791] = 246;
    exp_47_ram[792] = 23;
    exp_47_ram[793] = 7;
    exp_47_ram[794] = 223;
    exp_47_ram[795] = 181;
    exp_47_ram[796] = 55;
    exp_47_ram[797] = 7;
    exp_47_ram[798] = 255;
    exp_47_ram[799] = 128;
    exp_47_ram[800] = 246;
    exp_47_ram[801] = 6;
    exp_47_ram[802] = 5;
    exp_47_ram[803] = 5;
    exp_47_ram[804] = 231;
    exp_47_ram[805] = 5;
    exp_47_ram[806] = 5;
    exp_47_ram[807] = 7;
    exp_47_ram[808] = 231;
    exp_47_ram[809] = 231;
    exp_47_ram[810] = 0;
    exp_47_ram[811] = 215;
    exp_47_ram[812] = 247;
    exp_47_ram[813] = 247;
    exp_47_ram[814] = 199;
    exp_47_ram[815] = 7;
    exp_47_ram[816] = 69;
    exp_47_ram[817] = 69;
    exp_47_ram[818] = 31;
    exp_47_ram[819] = 21;
    exp_47_ram[820] = 21;
    exp_47_ram[821] = 31;
    exp_47_ram[822] = 0;
    exp_47_ram[823] = 0;
    exp_47_ram[824] = 53;
    exp_47_ram[825] = 7;
    exp_47_ram[826] = 1;
    exp_47_ram[827] = 64;
    exp_47_ram[828] = 129;
    exp_47_ram[829] = 17;
    exp_47_ram[830] = 5;
    exp_47_ram[831] = 95;
    exp_47_ram[832] = 16;
    exp_47_ram[833] = 5;
    exp_47_ram[834] = 0;
    exp_47_ram[835] = 4;
    exp_47_ram[836] = 31;
    exp_47_ram[837] = 21;
    exp_47_ram[838] = 193;
    exp_47_ram[839] = 129;
    exp_47_ram[840] = 7;
    exp_47_ram[841] = 1;
    exp_47_ram[842] = 0;
    exp_47_ram[843] = 0;
    exp_47_ram[844] = 7;
    exp_47_ram[845] = 0;
    exp_47_ram[846] = 213;
    exp_47_ram[847] = 215;
    exp_47_ram[848] = 7;
    exp_47_ram[849] = 213;
    exp_47_ram[850] = 128;
    exp_47_ram[851] = 224;
    exp_47_ram[852] = 215;
    exp_47_ram[853] = 16;
    exp_47_ram[854] = 240;
    exp_47_ram[855] = 229;
    exp_47_ram[856] = 1;
    exp_47_ram[857] = 17;
    exp_47_ram[858] = 159;
    exp_47_ram[859] = 193;
    exp_47_ram[860] = 160;
    exp_47_ram[861] = 199;
    exp_47_ram[862] = 7;
    exp_47_ram[863] = 1;
    exp_47_ram[864] = 0;
    exp_47_ram[865] = 224;
    exp_47_ram[866] = 7;
    exp_47_ram[867] = 0;
    exp_47_ram[868] = 0;
    exp_47_ram[869] = 7;
    exp_47_ram[870] = 71;
    exp_47_ram[871] = 71;
    exp_47_ram[872] = 6;
    exp_47_ram[873] = 135;
    exp_47_ram[874] = 213;
    exp_47_ram[875] = 0;
    exp_47_ram[876] = 5;
    exp_47_ram[877] = 197;
    exp_47_ram[878] = 167;
    exp_47_ram[879] = 213;
    exp_47_ram[880] = 1;
    exp_47_ram[881] = 245;
    exp_47_ram[882] = 17;
    exp_47_ram[883] = 159;
    exp_47_ram[884] = 193;
    exp_47_ram[885] = 1;
    exp_47_ram[886] = 0;
    exp_47_ram[887] = 1;
    exp_47_ram[888] = 81;
    exp_47_ram[889] = 69;
    exp_47_ram[890] = 145;
    exp_47_ram[891] = 1;
    exp_47_ram[892] = 129;
    exp_47_ram[893] = 33;
    exp_47_ram[894] = 49;
    exp_47_ram[895] = 65;
    exp_47_ram[896] = 17;
    exp_47_ram[897] = 97;
    exp_47_ram[898] = 5;
    exp_47_ram[899] = 32;
    exp_47_ram[900] = 0;
    exp_47_ram[901] = 0;
    exp_47_ram[902] = 202;
    exp_47_ram[903] = 4;
    exp_47_ram[904] = 138;
    exp_47_ram[905] = 10;
    exp_47_ram[906] = 1;
    exp_47_ram[907] = 0;
    exp_47_ram[908] = 10;
    exp_47_ram[909] = 155;
    exp_47_ram[910] = 4;
    exp_47_ram[911] = 4;
    exp_47_ram[912] = 159;
    exp_47_ram[913] = 10;
    exp_47_ram[914] = 95;
    exp_47_ram[915] = 169;
    exp_47_ram[916] = 37;
    exp_47_ram[917] = 55;
    exp_47_ram[918] = 5;
    exp_47_ram[919] = 20;
    exp_47_ram[920] = 95;
    exp_47_ram[921] = 4;
    exp_47_ram[922] = 159;
    exp_47_ram[923] = 160;
    exp_47_ram[924] = 4;
    exp_47_ram[925] = 213;
    exp_47_ram[926] = 95;
    exp_47_ram[927] = 169;
    exp_47_ram[928] = 37;
    exp_47_ram[929] = 55;
    exp_47_ram[930] = 5;
    exp_47_ram[931] = 20;
    exp_47_ram[932] = 31;
    exp_47_ram[933] = 138;
    exp_47_ram[934] = 74;
    exp_47_ram[935] = 10;
    exp_47_ram[936] = 55;
    exp_47_ram[937] = 231;
    exp_47_ram[938] = 87;
    exp_47_ram[939] = 231;
    exp_47_ram[940] = 70;
    exp_47_ram[941] = 199;
    exp_47_ram[942] = 71;
    exp_47_ram[943] = 39;
    exp_47_ram[944] = 202;
    exp_47_ram[945] = 247;
    exp_47_ram[946] = 247;
    exp_47_ram[947] = 231;
    exp_47_ram[948] = 198;
    exp_47_ram[949] = 247;
    exp_47_ram[950] = 215;
    exp_47_ram[951] = 1;
    exp_47_ram[952] = 244;
    exp_47_ram[953] = 151;
    exp_47_ram[954] = 228;
    exp_47_ram[955] = 215;
    exp_47_ram[956] = 5;
    exp_47_ram[957] = 245;
    exp_47_ram[958] = 247;
    exp_47_ram[959] = 31;
    exp_47_ram[960] = 164;
    exp_47_ram[961] = 245;
    exp_47_ram[962] = 149;
    exp_47_ram[963] = 244;
    exp_47_ram[964] = 37;
    exp_47_ram[965] = 244;
    exp_47_ram[966] = 52;
    exp_47_ram[967] = 181;
    exp_47_ram[968] = 193;
    exp_47_ram[969] = 133;
    exp_47_ram[970] = 129;
    exp_47_ram[971] = 65;
    exp_47_ram[972] = 1;
    exp_47_ram[973] = 193;
    exp_47_ram[974] = 129;
    exp_47_ram[975] = 65;
    exp_47_ram[976] = 1;
    exp_47_ram[977] = 1;
    exp_47_ram[978] = 0;
    exp_47_ram[979] = 1;
    exp_47_ram[980] = 17;
    exp_47_ram[981] = 129;
    exp_47_ram[982] = 5;
    exp_47_ram[983] = 95;
    exp_47_ram[984] = 0;
    exp_47_ram[985] = 199;
    exp_47_ram[986] = 0;
    exp_47_ram[987] = 15;
    exp_47_ram[988] = 0;
    exp_47_ram[989] = 135;
    exp_47_ram[990] = 245;
    exp_47_ram[991] = 4;
    exp_47_ram[992] = 164;
    exp_47_ram[993] = 4;
    exp_47_ram[994] = 193;
    exp_47_ram[995] = 129;
    exp_47_ram[996] = 0;
    exp_47_ram[997] = 1;
    exp_47_ram[998] = 0;
    exp_47_ram[999] = 1;
    exp_47_ram[1000] = 17;
    exp_47_ram[1001] = 129;
    exp_47_ram[1002] = 145;
    exp_47_ram[1003] = 33;
    exp_47_ram[1004] = 5;
    exp_47_ram[1005] = 5;
    exp_47_ram[1006] = 159;
    exp_47_ram[1007] = 0;
    exp_47_ram[1008] = 199;
    exp_47_ram[1009] = 0;
    exp_47_ram[1010] = 0;
    exp_47_ram[1011] = 15;
    exp_47_ram[1012] = 164;
    exp_47_ram[1013] = 164;
    exp_47_ram[1014] = 180;
    exp_47_ram[1015] = 137;
    exp_47_ram[1016] = 148;
    exp_47_ram[1017] = 137;
    exp_47_ram[1018] = 193;
    exp_47_ram[1019] = 129;
    exp_47_ram[1020] = 169;
    exp_47_ram[1021] = 65;
    exp_47_ram[1022] = 1;
    exp_47_ram[1023] = 1;
    exp_47_ram[1024] = 0;
    exp_47_ram[1025] = 1;
    exp_47_ram[1026] = 0;
    exp_47_ram[1027] = 145;
    exp_47_ram[1028] = 96;
    exp_47_ram[1029] = 5;
    exp_47_ram[1030] = 69;
    exp_47_ram[1031] = 1;
    exp_47_ram[1032] = 17;
    exp_47_ram[1033] = 129;
    exp_47_ram[1034] = 33;
    exp_47_ram[1035] = 49;
    exp_47_ram[1036] = 65;
    exp_47_ram[1037] = 31;
    exp_47_ram[1038] = 0;
    exp_47_ram[1039] = 80;
    exp_47_ram[1040] = 197;
    exp_47_ram[1041] = 129;
    exp_47_ram[1042] = 223;
    exp_47_ram[1043] = 132;
    exp_47_ram[1044] = 0;
    exp_47_ram[1045] = 73;
    exp_47_ram[1046] = 23;
    exp_47_ram[1047] = 245;
    exp_47_ram[1048] = 1;
    exp_47_ram[1049] = 0;
    exp_47_ram[1050] = 183;
    exp_47_ram[1051] = 48;
    exp_47_ram[1052] = 73;
    exp_47_ram[1053] = 31;
    exp_47_ram[1054] = 36;
    exp_47_ram[1055] = 4;
    exp_47_ram[1056] = 48;
    exp_47_ram[1057] = 68;
    exp_47_ram[1058] = 23;
    exp_47_ram[1059] = 245;
    exp_47_ram[1060] = 129;
    exp_47_ram[1061] = 183;
    exp_47_ram[1062] = 223;
    exp_47_ram[1063] = 36;
    exp_47_ram[1064] = 196;
    exp_47_ram[1065] = 160;
    exp_47_ram[1066] = 160;
    exp_47_ram[1067] = 80;
    exp_47_ram[1068] = 161;
    exp_47_ram[1069] = 129;
    exp_47_ram[1070] = 177;
    exp_47_ram[1071] = 36;
    exp_47_ram[1072] = 7;
    exp_47_ram[1073] = 244;
    exp_47_ram[1074] = 193;
    exp_47_ram[1075] = 160;
    exp_47_ram[1076] = 7;
    exp_47_ram[1077] = 244;
    exp_47_ram[1078] = 132;
    exp_47_ram[1079] = 80;
    exp_47_ram[1080] = 161;
    exp_47_ram[1081] = 129;
    exp_47_ram[1082] = 177;
    exp_47_ram[1083] = 68;
    exp_47_ram[1084] = 7;
    exp_47_ram[1085] = 244;
    exp_47_ram[1086] = 193;
    exp_47_ram[1087] = 160;
    exp_47_ram[1088] = 7;
    exp_47_ram[1089] = 244;
    exp_47_ram[1090] = 68;
    exp_47_ram[1091] = 80;
    exp_47_ram[1092] = 161;
    exp_47_ram[1093] = 129;
    exp_47_ram[1094] = 177;
    exp_47_ram[1095] = 68;
    exp_47_ram[1096] = 7;
    exp_47_ram[1097] = 244;
    exp_47_ram[1098] = 193;
    exp_47_ram[1099] = 160;
    exp_47_ram[1100] = 7;
    exp_47_ram[1101] = 244;
    exp_47_ram[1102] = 4;
    exp_47_ram[1103] = 80;
    exp_47_ram[1104] = 161;
    exp_47_ram[1105] = 129;
    exp_47_ram[1106] = 177;
    exp_47_ram[1107] = 36;
    exp_47_ram[1108] = 7;
    exp_47_ram[1109] = 244;
    exp_47_ram[1110] = 193;
    exp_47_ram[1111] = 128;
    exp_47_ram[1112] = 7;
    exp_47_ram[1113] = 244;
    exp_47_ram[1114] = 68;
    exp_47_ram[1115] = 197;
    exp_47_ram[1116] = 16;
    exp_47_ram[1117] = 161;
    exp_47_ram[1118] = 177;
    exp_47_ram[1119] = 129;
    exp_47_ram[1120] = 193;
    exp_47_ram[1121] = 64;
    exp_47_ram[1122] = 7;
    exp_47_ram[1123] = 244;
    exp_47_ram[1124] = 16;
    exp_47_ram[1125] = 161;
    exp_47_ram[1126] = 177;
    exp_47_ram[1127] = 129;
    exp_47_ram[1128] = 193;
    exp_47_ram[1129] = 160;
    exp_47_ram[1130] = 7;
    exp_47_ram[1131] = 244;
    exp_47_ram[1132] = 16;
    exp_47_ram[1133] = 161;
    exp_47_ram[1134] = 129;
    exp_47_ram[1135] = 177;
    exp_47_ram[1136] = 193;
    exp_47_ram[1137] = 7;
    exp_47_ram[1138] = 244;
    exp_47_ram[1139] = 193;
    exp_47_ram[1140] = 65;
    exp_47_ram[1141] = 1;
    exp_47_ram[1142] = 7;
    exp_47_ram[1143] = 244;
    exp_47_ram[1144] = 160;
    exp_47_ram[1145] = 244;
    exp_47_ram[1146] = 129;
    exp_47_ram[1147] = 129;
    exp_47_ram[1148] = 73;
    exp_47_ram[1149] = 193;
    exp_47_ram[1150] = 1;
    exp_47_ram[1151] = 0;
    exp_47_ram[1152] = 1;
    exp_47_ram[1153] = 97;
    exp_47_ram[1154] = 1;
    exp_47_ram[1155] = 129;
    exp_47_ram[1156] = 145;
    exp_47_ram[1157] = 33;
    exp_47_ram[1158] = 49;
    exp_47_ram[1159] = 81;
    exp_47_ram[1160] = 17;
    exp_47_ram[1161] = 65;
    exp_47_ram[1162] = 113;
    exp_47_ram[1163] = 129;
    exp_47_ram[1164] = 145;
    exp_47_ram[1165] = 5;
    exp_47_ram[1166] = 5;
    exp_47_ram[1167] = 6;
    exp_47_ram[1168] = 32;
    exp_47_ram[1169] = 64;
    exp_47_ram[1170] = 11;
    exp_47_ram[1171] = 9;
    exp_47_ram[1172] = 31;
    exp_47_ram[1173] = 160;
    exp_47_ram[1174] = 218;
    exp_47_ram[1175] = 11;
    exp_47_ram[1176] = 10;
    exp_47_ram[1177] = 143;
    exp_47_ram[1178] = 25;
    exp_47_ram[1179] = 9;
    exp_47_ram[1180] = 164;
    exp_47_ram[1181] = 164;
    exp_47_ram[1182] = 164;
    exp_47_ram[1183] = 74;
    exp_47_ram[1184] = 5;
    exp_47_ram[1185] = 233;
    exp_47_ram[1186] = 7;
    exp_47_ram[1187] = 31;
    exp_47_ram[1188] = 1;
    exp_47_ram[1189] = 0;
    exp_47_ram[1190] = 0;
    exp_47_ram[1191] = 12;
    exp_47_ram[1192] = 12;
    exp_47_ram[1193] = 9;
    exp_47_ram[1194] = 31;
    exp_47_ram[1195] = 12;
    exp_47_ram[1196] = 12;
    exp_47_ram[1197] = 5;
    exp_47_ram[1198] = 28;
    exp_47_ram[1199] = 15;
    exp_47_ram[1200] = 9;
    exp_47_ram[1201] = 164;
    exp_47_ram[1202] = 164;
    exp_47_ram[1203] = 164;
    exp_47_ram[1204] = 122;
    exp_47_ram[1205] = 122;
    exp_47_ram[1206] = 5;
    exp_47_ram[1207] = 249;
    exp_47_ram[1208] = 31;
    exp_47_ram[1209] = 1;
    exp_47_ram[1210] = 4;
    exp_47_ram[1211] = 5;
    exp_47_ram[1212] = 16;
    exp_47_ram[1213] = 177;
    exp_47_ram[1214] = 5;
    exp_47_ram[1215] = 161;
    exp_47_ram[1216] = 170;
    exp_47_ram[1217] = 193;
    exp_47_ram[1218] = 0;
    exp_47_ram[1219] = 5;
    exp_47_ram[1220] = 16;
    exp_47_ram[1221] = 177;
    exp_47_ram[1222] = 5;
    exp_47_ram[1223] = 161;
    exp_47_ram[1224] = 193;
    exp_47_ram[1225] = 192;
    exp_47_ram[1226] = 73;
    exp_47_ram[1227] = 80;
    exp_47_ram[1228] = 20;
    exp_47_ram[1229] = 161;
    exp_47_ram[1230] = 177;
    exp_47_ram[1231] = 180;
    exp_47_ram[1232] = 164;
    exp_47_ram[1233] = 36;
    exp_47_ram[1234] = 100;
    exp_47_ram[1235] = 52;
    exp_47_ram[1236] = 154;
    exp_47_ram[1237] = 244;
    exp_47_ram[1238] = 112;
    exp_47_ram[1239] = 143;
    exp_47_ram[1240] = 164;
    exp_47_ram[1241] = 68;
    exp_47_ram[1242] = 193;
    exp_47_ram[1243] = 4;
    exp_47_ram[1244] = 129;
    exp_47_ram[1245] = 65;
    exp_47_ram[1246] = 1;
    exp_47_ram[1247] = 193;
    exp_47_ram[1248] = 129;
    exp_47_ram[1249] = 65;
    exp_47_ram[1250] = 1;
    exp_47_ram[1251] = 193;
    exp_47_ram[1252] = 129;
    exp_47_ram[1253] = 65;
    exp_47_ram[1254] = 1;
    exp_47_ram[1255] = 0;
    exp_47_ram[1256] = 1;
    exp_47_ram[1257] = 81;
    exp_47_ram[1258] = 69;
    exp_47_ram[1259] = 144;
    exp_47_ram[1260] = 145;
    exp_47_ram[1261] = 33;
    exp_47_ram[1262] = 65;
    exp_47_ram[1263] = 240;
    exp_47_ram[1264] = 16;
    exp_47_ram[1265] = 64;
    exp_47_ram[1266] = 5;
    exp_47_ram[1267] = 129;
    exp_47_ram[1268] = 1;
    exp_47_ram[1269] = 17;
    exp_47_ram[1270] = 241;
    exp_47_ram[1271] = 129;
    exp_47_ram[1272] = 49;
    exp_47_ram[1273] = 65;
    exp_47_ram[1274] = 145;
    exp_47_ram[1275] = 81;
    exp_47_ram[1276] = 1;
    exp_47_ram[1277] = 1;
    exp_47_ram[1278] = 1;
    exp_47_ram[1279] = 143;
    exp_47_ram[1280] = 1;
    exp_47_ram[1281] = 159;
    exp_47_ram[1282] = 5;
    exp_47_ram[1283] = 5;
    exp_47_ram[1284] = 129;
    exp_47_ram[1285] = 223;
    exp_47_ram[1286] = 1;
    exp_47_ram[1287] = 65;
    exp_47_ram[1288] = 64;
    exp_47_ram[1289] = 129;
    exp_47_ram[1290] = 231;
    exp_47_ram[1291] = 1;
    exp_47_ram[1292] = 241;
    exp_47_ram[1293] = 15;
    exp_47_ram[1294] = 1;
    exp_47_ram[1295] = 31;
    exp_47_ram[1296] = 32;
    exp_47_ram[1297] = 64;
    exp_47_ram[1298] = 5;
    exp_47_ram[1299] = 5;
    exp_47_ram[1300] = 1;
    exp_47_ram[1301] = 193;
    exp_47_ram[1302] = 241;
    exp_47_ram[1303] = 65;
    exp_47_ram[1304] = 145;
    exp_47_ram[1305] = 81;
    exp_47_ram[1306] = 1;
    exp_47_ram[1307] = 1;
    exp_47_ram[1308] = 79;
    exp_47_ram[1309] = 1;
    exp_47_ram[1310] = 95;
    exp_47_ram[1311] = 5;
    exp_47_ram[1312] = 5;
    exp_47_ram[1313] = 193;
    exp_47_ram[1314] = 159;
    exp_47_ram[1315] = 65;
    exp_47_ram[1316] = 129;
    exp_47_ram[1317] = 64;
    exp_47_ram[1318] = 193;
    exp_47_ram[1319] = 231;
    exp_47_ram[1320] = 1;
    exp_47_ram[1321] = 241;
    exp_47_ram[1322] = 207;
    exp_47_ram[1323] = 1;
    exp_47_ram[1324] = 223;
    exp_47_ram[1325] = 5;
    exp_47_ram[1326] = 5;
    exp_47_ram[1327] = 64;
    exp_47_ram[1328] = 9;
    exp_47_ram[1329] = 1;
    exp_47_ram[1330] = 207;
    exp_47_ram[1331] = 1;
    exp_47_ram[1332] = 223;
    exp_47_ram[1333] = 149;
    exp_47_ram[1334] = 5;
    exp_47_ram[1335] = 5;
    exp_47_ram[1336] = 180;
    exp_47_ram[1337] = 69;
    exp_47_ram[1338] = 16;
    exp_47_ram[1339] = 244;
    exp_47_ram[1340] = 135;
    exp_47_ram[1341] = 233;
    exp_47_ram[1342] = 0;
    exp_47_ram[1343] = 193;
    exp_47_ram[1344] = 129;
    exp_47_ram[1345] = 65;
    exp_47_ram[1346] = 1;
    exp_47_ram[1347] = 193;
    exp_47_ram[1348] = 129;
    exp_47_ram[1349] = 65;
    exp_47_ram[1350] = 1;
    exp_47_ram[1351] = 0;
    exp_47_ram[1352] = 1;
    exp_47_ram[1353] = 5;
    exp_47_ram[1354] = 33;
    exp_47_ram[1355] = 64;
    exp_47_ram[1356] = 5;
    exp_47_ram[1357] = 193;
    exp_47_ram[1358] = 17;
    exp_47_ram[1359] = 129;
    exp_47_ram[1360] = 145;
    exp_47_ram[1361] = 49;
    exp_47_ram[1362] = 207;
    exp_47_ram[1363] = 64;
    exp_47_ram[1364] = 193;
    exp_47_ram[1365] = 1;
    exp_47_ram[1366] = 9;
    exp_47_ram[1367] = 143;
    exp_47_ram[1368] = 1;
    exp_47_ram[1369] = 159;
    exp_47_ram[1370] = 5;
    exp_47_ram[1371] = 5;
    exp_47_ram[1372] = 48;
    exp_47_ram[1373] = 255;
    exp_47_ram[1374] = 7;
    exp_47_ram[1375] = 245;
    exp_47_ram[1376] = 167;
    exp_47_ram[1377] = 245;
    exp_47_ram[1378] = 7;
    exp_47_ram[1379] = 135;
    exp_47_ram[1380] = 4;
    exp_47_ram[1381] = 4;
    exp_47_ram[1382] = 1;
    exp_47_ram[1383] = 95;
    exp_47_ram[1384] = 64;
    exp_47_ram[1385] = 1;
    exp_47_ram[1386] = 9;
    exp_47_ram[1387] = 143;
    exp_47_ram[1388] = 48;
    exp_47_ram[1389] = 16;
    exp_47_ram[1390] = 249;
    exp_47_ram[1391] = 193;
    exp_47_ram[1392] = 4;
    exp_47_ram[1393] = 129;
    exp_47_ram[1394] = 1;
    exp_47_ram[1395] = 193;
    exp_47_ram[1396] = 4;
    exp_47_ram[1397] = 65;
    exp_47_ram[1398] = 1;
    exp_47_ram[1399] = 0;
    exp_47_ram[1400] = 9;
    exp_47_ram[1401] = 64;
    exp_47_ram[1402] = 193;
    exp_47_ram[1403] = 1;
    exp_47_ram[1404] = 79;
    exp_47_ram[1405] = 1;
    exp_47_ram[1406] = 159;
    exp_47_ram[1407] = 0;
    exp_47_ram[1408] = 5;
    exp_47_ram[1409] = 0;
    exp_47_ram[1410] = 7;
    exp_47_ram[1411] = 244;
    exp_47_ram[1412] = 244;
    exp_47_ram[1413] = 228;
    exp_47_ram[1414] = 7;
    exp_47_ram[1415] = 95;
    exp_47_ram[1416] = 9;
    exp_47_ram[1417] = 64;
    exp_47_ram[1418] = 193;
    exp_47_ram[1419] = 1;
    exp_47_ram[1420] = 79;
    exp_47_ram[1421] = 1;
    exp_47_ram[1422] = 159;
    exp_47_ram[1423] = 169;
    exp_47_ram[1424] = 223;
    exp_47_ram[1425] = 9;
    exp_47_ram[1426] = 95;
    exp_47_ram[1427] = 1;
    exp_47_ram[1428] = 5;
    exp_47_ram[1429] = 5;
    exp_47_ram[1430] = 193;
    exp_47_ram[1431] = 17;
    exp_47_ram[1432] = 31;
    exp_47_ram[1433] = 193;
    exp_47_ram[1434] = 64;
    exp_47_ram[1435] = 1;
    exp_47_ram[1436] = 79;
    exp_47_ram[1437] = 1;
    exp_47_ram[1438] = 159;
    exp_47_ram[1439] = 193;
    exp_47_ram[1440] = 1;
    exp_47_ram[1441] = 0;
    exp_47_ram[1442] = 5;
    exp_47_ram[1443] = 69;
    exp_47_ram[1444] = 1;
    exp_47_ram[1445] = 1;
    exp_47_ram[1446] = 17;
    exp_47_ram[1447] = 129;
    exp_47_ram[1448] = 31;
    exp_47_ram[1449] = 0;
    exp_47_ram[1450] = 1;
    exp_47_ram[1451] = 4;
    exp_47_ram[1452] = 64;
    exp_47_ram[1453] = 15;
    exp_47_ram[1454] = 193;
    exp_47_ram[1455] = 4;
    exp_47_ram[1456] = 129;
    exp_47_ram[1457] = 1;
    exp_47_ram[1458] = 0;
    exp_47_ram[1459] = 1;
    exp_47_ram[1460] = 145;
    exp_47_ram[1461] = 33;
    exp_47_ram[1462] = 69;
    exp_47_ram[1463] = 5;
    exp_47_ram[1464] = 17;
    exp_47_ram[1465] = 4;
    exp_47_ram[1466] = 9;
    exp_47_ram[1467] = 129;
    exp_47_ram[1468] = 49;
    exp_47_ram[1469] = 159;
    exp_47_ram[1470] = 0;
    exp_47_ram[1471] = 5;
    exp_47_ram[1472] = 0;
    exp_47_ram[1473] = 6;
    exp_47_ram[1474] = 38;
    exp_47_ram[1475] = 197;
    exp_47_ram[1476] = 150;
    exp_47_ram[1477] = 1;
    exp_47_ram[1478] = 159;
    exp_47_ram[1479] = 0;
    exp_47_ram[1480] = 1;
    exp_47_ram[1481] = 64;
    exp_47_ram[1482] = 4;
    exp_47_ram[1483] = 143;
    exp_47_ram[1484] = 9;
    exp_47_ram[1485] = 4;
    exp_47_ram[1486] = 95;
    exp_47_ram[1487] = 4;
    exp_47_ram[1488] = 169;
    exp_47_ram[1489] = 193;
    exp_47_ram[1490] = 4;
    exp_47_ram[1491] = 129;
    exp_47_ram[1492] = 65;
    exp_47_ram[1493] = 1;
    exp_47_ram[1494] = 193;
    exp_47_ram[1495] = 1;
    exp_47_ram[1496] = 0;
    exp_47_ram[1497] = 1;
    exp_47_ram[1498] = 17;
    exp_47_ram[1499] = 31;
    exp_47_ram[1500] = 193;
    exp_47_ram[1501] = 1;
    exp_47_ram[1502] = 223;
    exp_47_ram[1503] = 1;
    exp_47_ram[1504] = 17;
    exp_47_ram[1505] = 129;
    exp_47_ram[1506] = 1;
    exp_47_ram[1507] = 0;
    exp_47_ram[1508] = 7;
    exp_47_ram[1509] = 143;
    exp_47_ram[1510] = 0;
    exp_47_ram[1511] = 199;
    exp_47_ram[1512] = 207;
    exp_47_ram[1513] = 193;
    exp_47_ram[1514] = 129;
    exp_47_ram[1515] = 1;
    exp_47_ram[1516] = 0;
    exp_47_ram[1517] = 1;
    exp_47_ram[1518] = 17;
    exp_47_ram[1519] = 129;
    exp_47_ram[1520] = 33;
    exp_47_ram[1521] = 49;
    exp_47_ram[1522] = 65;
    exp_47_ram[1523] = 81;
    exp_47_ram[1524] = 97;
    exp_47_ram[1525] = 113;
    exp_47_ram[1526] = 1;
    exp_47_ram[1527] = 0;
    exp_47_ram[1528] = 71;
    exp_47_ram[1529] = 143;
    exp_47_ram[1530] = 128;
    exp_47_ram[1531] = 244;
    exp_47_ram[1532] = 128;
    exp_47_ram[1533] = 244;
    exp_47_ram[1534] = 16;
    exp_47_ram[1535] = 244;
    exp_47_ram[1536] = 16;
    exp_47_ram[1537] = 244;
    exp_47_ram[1538] = 80;
    exp_47_ram[1539] = 244;
    exp_47_ram[1540] = 4;
    exp_47_ram[1541] = 240;
    exp_47_ram[1542] = 244;
    exp_47_ram[1543] = 196;
    exp_47_ram[1544] = 7;
    exp_47_ram[1545] = 223;
    exp_47_ram[1546] = 5;
    exp_47_ram[1547] = 5;
    exp_47_ram[1548] = 228;
    exp_47_ram[1549] = 244;
    exp_47_ram[1550] = 196;
    exp_47_ram[1551] = 7;
    exp_47_ram[1552] = 79;
    exp_47_ram[1553] = 5;
    exp_47_ram[1554] = 0;
    exp_47_ram[1555] = 199;
    exp_47_ram[1556] = 7;
    exp_47_ram[1557] = 143;
    exp_47_ram[1558] = 5;
    exp_47_ram[1559] = 7;
    exp_47_ram[1560] = 0;
    exp_47_ram[1561] = 135;
    exp_47_ram[1562] = 79;
    exp_47_ram[1563] = 0;
    exp_47_ram[1564] = 4;
    exp_47_ram[1565] = 7;
    exp_47_ram[1566] = 95;
    exp_47_ram[1567] = 5;
    exp_47_ram[1568] = 7;
    exp_47_ram[1569] = 15;
    exp_47_ram[1570] = 5;
    exp_47_ram[1571] = 0;
    exp_47_ram[1572] = 7;
    exp_47_ram[1573] = 7;
    exp_47_ram[1574] = 79;
    exp_47_ram[1575] = 5;
    exp_47_ram[1576] = 7;
    exp_47_ram[1577] = 0;
    exp_47_ram[1578] = 199;
    exp_47_ram[1579] = 15;
    exp_47_ram[1580] = 192;
    exp_47_ram[1581] = 4;
    exp_47_ram[1582] = 7;
    exp_47_ram[1583] = 223;
    exp_47_ram[1584] = 5;
    exp_47_ram[1585] = 7;
    exp_47_ram[1586] = 207;
    exp_47_ram[1587] = 5;
    exp_47_ram[1588] = 0;
    exp_47_ram[1589] = 199;
    exp_47_ram[1590] = 7;
    exp_47_ram[1591] = 15;
    exp_47_ram[1592] = 5;
    exp_47_ram[1593] = 7;
    exp_47_ram[1594] = 0;
    exp_47_ram[1595] = 71;
    exp_47_ram[1596] = 207;
    exp_47_ram[1597] = 128;
    exp_47_ram[1598] = 4;
    exp_47_ram[1599] = 7;
    exp_47_ram[1600] = 95;
    exp_47_ram[1601] = 5;
    exp_47_ram[1602] = 0;
    exp_47_ram[1603] = 7;
    exp_47_ram[1604] = 7;
    exp_47_ram[1605] = 143;
    exp_47_ram[1606] = 5;
    exp_47_ram[1607] = 7;
    exp_47_ram[1608] = 0;
    exp_47_ram[1609] = 199;
    exp_47_ram[1610] = 79;
    exp_47_ram[1611] = 0;
    exp_47_ram[1612] = 128;
    exp_47_ram[1613] = 244;
    exp_47_ram[1614] = 128;
    exp_47_ram[1615] = 244;
    exp_47_ram[1616] = 16;
    exp_47_ram[1617] = 244;
    exp_47_ram[1618] = 16;
    exp_47_ram[1619] = 244;
    exp_47_ram[1620] = 80;
    exp_47_ram[1621] = 244;
    exp_47_ram[1622] = 4;
    exp_47_ram[1623] = 16;
    exp_47_ram[1624] = 244;
    exp_47_ram[1625] = 196;
    exp_47_ram[1626] = 7;
    exp_47_ram[1627] = 95;
    exp_47_ram[1628] = 5;
    exp_47_ram[1629] = 5;
    exp_47_ram[1630] = 228;
    exp_47_ram[1631] = 244;
    exp_47_ram[1632] = 196;
    exp_47_ram[1633] = 7;
    exp_47_ram[1634] = 207;
    exp_47_ram[1635] = 5;
    exp_47_ram[1636] = 0;
    exp_47_ram[1637] = 199;
    exp_47_ram[1638] = 7;
    exp_47_ram[1639] = 15;
    exp_47_ram[1640] = 5;
    exp_47_ram[1641] = 7;
    exp_47_ram[1642] = 0;
    exp_47_ram[1643] = 71;
    exp_47_ram[1644] = 207;
    exp_47_ram[1645] = 128;
    exp_47_ram[1646] = 4;
    exp_47_ram[1647] = 7;
    exp_47_ram[1648] = 223;
    exp_47_ram[1649] = 5;
    exp_47_ram[1650] = 7;
    exp_47_ram[1651] = 143;
    exp_47_ram[1652] = 5;
    exp_47_ram[1653] = 0;
    exp_47_ram[1654] = 7;
    exp_47_ram[1655] = 7;
    exp_47_ram[1656] = 207;
    exp_47_ram[1657] = 5;
    exp_47_ram[1658] = 7;
    exp_47_ram[1659] = 0;
    exp_47_ram[1660] = 199;
    exp_47_ram[1661] = 143;
    exp_47_ram[1662] = 64;
    exp_47_ram[1663] = 4;
    exp_47_ram[1664] = 7;
    exp_47_ram[1665] = 95;
    exp_47_ram[1666] = 5;
    exp_47_ram[1667] = 7;
    exp_47_ram[1668] = 79;
    exp_47_ram[1669] = 5;
    exp_47_ram[1670] = 0;
    exp_47_ram[1671] = 199;
    exp_47_ram[1672] = 7;
    exp_47_ram[1673] = 143;
    exp_47_ram[1674] = 5;
    exp_47_ram[1675] = 7;
    exp_47_ram[1676] = 0;
    exp_47_ram[1677] = 71;
    exp_47_ram[1678] = 79;
    exp_47_ram[1679] = 0;
    exp_47_ram[1680] = 4;
    exp_47_ram[1681] = 7;
    exp_47_ram[1682] = 223;
    exp_47_ram[1683] = 5;
    exp_47_ram[1684] = 0;
    exp_47_ram[1685] = 7;
    exp_47_ram[1686] = 7;
    exp_47_ram[1687] = 15;
    exp_47_ram[1688] = 5;
    exp_47_ram[1689] = 7;
    exp_47_ram[1690] = 0;
    exp_47_ram[1691] = 199;
    exp_47_ram[1692] = 207;
    exp_47_ram[1693] = 128;
    exp_47_ram[1694] = 128;
    exp_47_ram[1695] = 244;
    exp_47_ram[1696] = 128;
    exp_47_ram[1697] = 244;
    exp_47_ram[1698] = 16;
    exp_47_ram[1699] = 244;
    exp_47_ram[1700] = 16;
    exp_47_ram[1701] = 244;
    exp_47_ram[1702] = 80;
    exp_47_ram[1703] = 244;
    exp_47_ram[1704] = 4;
    exp_47_ram[1705] = 4;
    exp_47_ram[1706] = 196;
    exp_47_ram[1707] = 7;
    exp_47_ram[1708] = 31;
    exp_47_ram[1709] = 5;
    exp_47_ram[1710] = 5;
    exp_47_ram[1711] = 228;
    exp_47_ram[1712] = 244;
    exp_47_ram[1713] = 196;
    exp_47_ram[1714] = 7;
    exp_47_ram[1715] = 143;
    exp_47_ram[1716] = 5;
    exp_47_ram[1717] = 0;
    exp_47_ram[1718] = 7;
    exp_47_ram[1719] = 7;
    exp_47_ram[1720] = 207;
    exp_47_ram[1721] = 5;
    exp_47_ram[1722] = 7;
    exp_47_ram[1723] = 0;
    exp_47_ram[1724] = 71;
    exp_47_ram[1725] = 143;
    exp_47_ram[1726] = 64;
    exp_47_ram[1727] = 4;
    exp_47_ram[1728] = 7;
    exp_47_ram[1729] = 159;
    exp_47_ram[1730] = 5;
    exp_47_ram[1731] = 7;
    exp_47_ram[1732] = 79;
    exp_47_ram[1733] = 5;
    exp_47_ram[1734] = 0;
    exp_47_ram[1735] = 199;
    exp_47_ram[1736] = 7;
    exp_47_ram[1737] = 143;
    exp_47_ram[1738] = 5;
    exp_47_ram[1739] = 7;
    exp_47_ram[1740] = 0;
    exp_47_ram[1741] = 135;
    exp_47_ram[1742] = 79;
    exp_47_ram[1743] = 0;
    exp_47_ram[1744] = 4;
    exp_47_ram[1745] = 7;
    exp_47_ram[1746] = 31;
    exp_47_ram[1747] = 5;
    exp_47_ram[1748] = 7;
    exp_47_ram[1749] = 15;
    exp_47_ram[1750] = 5;
    exp_47_ram[1751] = 0;
    exp_47_ram[1752] = 7;
    exp_47_ram[1753] = 7;
    exp_47_ram[1754] = 79;
    exp_47_ram[1755] = 5;
    exp_47_ram[1756] = 7;
    exp_47_ram[1757] = 0;
    exp_47_ram[1758] = 7;
    exp_47_ram[1759] = 15;
    exp_47_ram[1760] = 192;
    exp_47_ram[1761] = 4;
    exp_47_ram[1762] = 7;
    exp_47_ram[1763] = 159;
    exp_47_ram[1764] = 5;
    exp_47_ram[1765] = 0;
    exp_47_ram[1766] = 199;
    exp_47_ram[1767] = 7;
    exp_47_ram[1768] = 207;
    exp_47_ram[1769] = 5;
    exp_47_ram[1770] = 7;
    exp_47_ram[1771] = 0;
    exp_47_ram[1772] = 135;
    exp_47_ram[1773] = 159;
    exp_47_ram[1774] = 64;
    exp_47_ram[1775] = 0;
    exp_47_ram[1776] = 7;
    exp_47_ram[1777] = 159;
    exp_47_ram[1778] = 128;
    exp_47_ram[1779] = 244;
    exp_47_ram[1780] = 32;
    exp_47_ram[1781] = 244;
    exp_47_ram[1782] = 208;
    exp_47_ram[1783] = 244;
    exp_47_ram[1784] = 4;
    exp_47_ram[1785] = 176;
    exp_47_ram[1786] = 244;
    exp_47_ram[1787] = 112;
    exp_47_ram[1788] = 244;
    exp_47_ram[1789] = 240;
    exp_47_ram[1790] = 244;
    exp_47_ram[1791] = 196;
    exp_47_ram[1792] = 7;
    exp_47_ram[1793] = 223;
    exp_47_ram[1794] = 5;
    exp_47_ram[1795] = 5;
    exp_47_ram[1796] = 228;
    exp_47_ram[1797] = 244;
    exp_47_ram[1798] = 4;
    exp_47_ram[1799] = 68;
    exp_47_ram[1800] = 7;
    exp_47_ram[1801] = 7;
    exp_47_ram[1802] = 79;
    exp_47_ram[1803] = 79;
    exp_47_ram[1804] = 164;
    exp_47_ram[1805] = 180;
    exp_47_ram[1806] = 4;
    exp_47_ram[1807] = 128;
    exp_47_ram[1808] = 0;
    exp_47_ram[1809] = 207;
    exp_47_ram[1810] = 5;
    exp_47_ram[1811] = 5;
    exp_47_ram[1812] = 132;
    exp_47_ram[1813] = 196;
    exp_47_ram[1814] = 7;
    exp_47_ram[1815] = 7;
    exp_47_ram[1816] = 15;
    exp_47_ram[1817] = 5;
    exp_47_ram[1818] = 5;
    exp_47_ram[1819] = 0;
    exp_47_ram[1820] = 199;
    exp_47_ram[1821] = 7;
    exp_47_ram[1822] = 223;
    exp_47_ram[1823] = 5;
    exp_47_ram[1824] = 5;
    exp_47_ram[1825] = 7;
    exp_47_ram[1826] = 7;
    exp_47_ram[1827] = 11;
    exp_47_ram[1828] = 11;
    exp_47_ram[1829] = 223;
    exp_47_ram[1830] = 5;
    exp_47_ram[1831] = 7;
    exp_47_ram[1832] = 0;
    exp_47_ram[1833] = 199;
    exp_47_ram[1834] = 7;
    exp_47_ram[1835] = 0;
    exp_47_ram[1836] = 132;
    exp_47_ram[1837] = 196;
    exp_47_ram[1838] = 70;
    exp_47_ram[1839] = 7;
    exp_47_ram[1840] = 197;
    exp_47_ram[1841] = 86;
    exp_47_ram[1842] = 245;
    exp_47_ram[1843] = 6;
    exp_47_ram[1844] = 228;
    exp_47_ram[1845] = 244;
    exp_47_ram[1846] = 0;
    exp_47_ram[1847] = 15;
    exp_47_ram[1848] = 5;
    exp_47_ram[1849] = 5;
    exp_47_ram[1850] = 228;
    exp_47_ram[1851] = 244;
    exp_47_ram[1852] = 4;
    exp_47_ram[1853] = 7;
    exp_47_ram[1854] = 223;
    exp_47_ram[1855] = 5;
    exp_47_ram[1856] = 7;
    exp_47_ram[1857] = 159;
    exp_47_ram[1858] = 68;
    exp_47_ram[1859] = 23;
    exp_47_ram[1860] = 244;
    exp_47_ram[1861] = 68;
    exp_47_ram[1862] = 144;
    exp_47_ram[1863] = 231;
    exp_47_ram[1864] = 128;
    exp_47_ram[1865] = 244;
    exp_47_ram[1866] = 144;
    exp_47_ram[1867] = 244;
    exp_47_ram[1868] = 144;
    exp_47_ram[1869] = 244;
    exp_47_ram[1870] = 16;
    exp_47_ram[1871] = 244;
    exp_47_ram[1872] = 176;
    exp_47_ram[1873] = 244;
    exp_47_ram[1874] = 112;
    exp_47_ram[1875] = 244;
    exp_47_ram[1876] = 16;
    exp_47_ram[1877] = 244;
    exp_47_ram[1878] = 196;
    exp_47_ram[1879] = 7;
    exp_47_ram[1880] = 15;
    exp_47_ram[1881] = 5;
    exp_47_ram[1882] = 5;
    exp_47_ram[1883] = 228;
    exp_47_ram[1884] = 244;
    exp_47_ram[1885] = 196;
    exp_47_ram[1886] = 7;
    exp_47_ram[1887] = 143;
    exp_47_ram[1888] = 5;
    exp_47_ram[1889] = 7;
    exp_47_ram[1890] = 95;
    exp_47_ram[1891] = 4;
    exp_47_ram[1892] = 7;
    exp_47_ram[1893] = 31;
    exp_47_ram[1894] = 5;
    exp_47_ram[1895] = 7;
    exp_47_ram[1896] = 223;
    exp_47_ram[1897] = 4;
    exp_47_ram[1898] = 68;
    exp_47_ram[1899] = 7;
    exp_47_ram[1900] = 7;
    exp_47_ram[1901] = 143;
    exp_47_ram[1902] = 0;
    exp_47_ram[1903] = 15;
    exp_47_ram[1904] = 5;
    exp_47_ram[1905] = 5;
    exp_47_ram[1906] = 228;
    exp_47_ram[1907] = 244;
    exp_47_ram[1908] = 4;
    exp_47_ram[1909] = 7;
    exp_47_ram[1910] = 223;
    exp_47_ram[1911] = 5;
    exp_47_ram[1912] = 7;
    exp_47_ram[1913] = 159;
    exp_47_ram[1914] = 159;
    exp_47_ram[1915] = 164;
    exp_47_ram[1916] = 180;
    exp_47_ram[1917] = 4;
    exp_47_ram[1918] = 128;
    exp_47_ram[1919] = 0;
    exp_47_ram[1920] = 31;
    exp_47_ram[1921] = 5;
    exp_47_ram[1922] = 5;
    exp_47_ram[1923] = 132;
    exp_47_ram[1924] = 196;
    exp_47_ram[1925] = 7;
    exp_47_ram[1926] = 7;
    exp_47_ram[1927] = 95;
    exp_47_ram[1928] = 5;
    exp_47_ram[1929] = 5;
    exp_47_ram[1930] = 0;
    exp_47_ram[1931] = 199;
    exp_47_ram[1932] = 7;
    exp_47_ram[1933] = 15;
    exp_47_ram[1934] = 5;
    exp_47_ram[1935] = 5;
    exp_47_ram[1936] = 7;
    exp_47_ram[1937] = 7;
    exp_47_ram[1938] = 10;
    exp_47_ram[1939] = 10;
    exp_47_ram[1940] = 15;
    exp_47_ram[1941] = 5;
    exp_47_ram[1942] = 7;
    exp_47_ram[1943] = 0;
    exp_47_ram[1944] = 199;
    exp_47_ram[1945] = 7;
    exp_47_ram[1946] = 0;
    exp_47_ram[1947] = 132;
    exp_47_ram[1948] = 196;
    exp_47_ram[1949] = 38;
    exp_47_ram[1950] = 7;
    exp_47_ram[1951] = 197;
    exp_47_ram[1952] = 54;
    exp_47_ram[1953] = 245;
    exp_47_ram[1954] = 6;
    exp_47_ram[1955] = 228;
    exp_47_ram[1956] = 244;
    exp_47_ram[1957] = 0;
    exp_47_ram[1958] = 79;
    exp_47_ram[1959] = 5;
    exp_47_ram[1960] = 5;
    exp_47_ram[1961] = 228;
    exp_47_ram[1962] = 244;
    exp_47_ram[1963] = 4;
    exp_47_ram[1964] = 7;
    exp_47_ram[1965] = 31;
    exp_47_ram[1966] = 5;
    exp_47_ram[1967] = 7;
    exp_47_ram[1968] = 223;
    exp_47_ram[1969] = 4;
    exp_47_ram[1970] = 23;
    exp_47_ram[1971] = 244;
    exp_47_ram[1972] = 4;
    exp_47_ram[1973] = 144;
    exp_47_ram[1974] = 231;
    exp_47_ram[1975] = 193;
    exp_47_ram[1976] = 129;
    exp_47_ram[1977] = 65;
    exp_47_ram[1978] = 1;
    exp_47_ram[1979] = 193;
    exp_47_ram[1980] = 129;
    exp_47_ram[1981] = 65;
    exp_47_ram[1982] = 1;
    exp_47_ram[1983] = 1;
    exp_47_ram[1984] = 0;
    exp_47_ram[1985] = 1;
    exp_47_ram[1986] = 17;
    exp_47_ram[1987] = 129;
    exp_47_ram[1988] = 1;
    exp_47_ram[1989] = 31;
    exp_47_ram[1990] = 95;
    exp_47_ram[1991] = 0;
    exp_47_ram[1992] = 193;
    exp_47_ram[1993] = 129;
    exp_47_ram[1994] = 1;
    exp_47_ram[1995] = 0;
    exp_47_ram[1996] = 5;
    exp_47_ram[1997] = 5;
    exp_47_ram[1998] = 181;
    exp_47_ram[1999] = 1;
    exp_47_ram[2000] = 183;
    exp_47_ram[2001] = 7;
    exp_47_ram[2002] = 5;
    exp_47_ram[2003] = 21;
    exp_47_ram[2004] = 245;
    exp_47_ram[2005] = 1;
    exp_47_ram[2006] = 0;
    exp_47_ram[2007] = 176;
    exp_47_ram[2008] = 245;
    exp_47_ram[2009] = 245;
    exp_47_ram[2010] = 223;
    exp_47_ram[2011] = 250;
    exp_47_ram[2012] = 0;
    exp_47_ram[2013] = 110;
    exp_47_ram[2014] = 84;
    exp_47_ram[2015] = 101;
    exp_47_ram[2016] = 117;
    exp_47_ram[2017] = 83;
    exp_47_ram[2018] = 0;
    exp_47_ram[2019] = 110;
    exp_47_ram[2020] = 77;
    exp_47_ram[2021] = 112;
    exp_47_ram[2022] = 121;
    exp_47_ram[2023] = 74;
    exp_47_ram[2024] = 117;
    exp_47_ram[2025] = 112;
    exp_47_ram[2026] = 78;
    exp_47_ram[2027] = 101;
    exp_47_ram[2028] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_45) begin
      exp_47_ram[exp_41] <= exp_43;
    end
  end
  assign exp_47 = exp_47_ram[exp_42];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_73) begin
        exp_47_ram[exp_69] <= exp_71;
    end
  end
  assign exp_75 = exp_47_ram[exp_70];
  assign exp_74 = exp_88;
  assign exp_88 = 1;
  assign exp_70 = exp_87;
  assign exp_87 = exp_8[31:2];
  assign exp_73 = exp_84;
  assign exp_84 = 0;
  assign exp_69 = exp_83;
  assign exp_83 = 0;
  assign exp_71 = exp_83;
  assign exp_46 = exp_123;
  assign exp_123 = 1;
  assign exp_42 = exp_122;
  assign exp_122 = exp_10[31:2];
  assign exp_45 = exp_111;
  assign exp_111 = exp_109 & exp_110;
  assign exp_109 = exp_14 & exp_15;
  assign exp_110 = exp_16[2:2];
  assign exp_41 = exp_107;
  assign exp_107 = exp_10[31:2];
  assign exp_43 = exp_108;
  assign exp_108 = exp_11[23:16];

  //Create RAM
  reg [7:0] exp_40_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_40_ram[0] = 0;
    exp_40_ram[1] = 1;
    exp_40_ram[2] = 1;
    exp_40_ram[3] = 2;
    exp_40_ram[4] = 2;
    exp_40_ram[5] = 3;
    exp_40_ram[6] = 3;
    exp_40_ram[7] = 4;
    exp_40_ram[8] = 4;
    exp_40_ram[9] = 5;
    exp_40_ram[10] = 5;
    exp_40_ram[11] = 6;
    exp_40_ram[12] = 6;
    exp_40_ram[13] = 7;
    exp_40_ram[14] = 7;
    exp_40_ram[15] = 8;
    exp_40_ram[16] = 8;
    exp_40_ram[17] = 9;
    exp_40_ram[18] = 9;
    exp_40_ram[19] = 10;
    exp_40_ram[20] = 10;
    exp_40_ram[21] = 11;
    exp_40_ram[22] = 11;
    exp_40_ram[23] = 12;
    exp_40_ram[24] = 12;
    exp_40_ram[25] = 13;
    exp_40_ram[26] = 13;
    exp_40_ram[27] = 14;
    exp_40_ram[28] = 14;
    exp_40_ram[29] = 15;
    exp_40_ram[30] = 15;
    exp_40_ram[31] = 65;
    exp_40_ram[32] = 1;
    exp_40_ram[33] = 16;
    exp_40_ram[34] = 0;
    exp_40_ram[35] = 8;
    exp_40_ram[36] = 135;
    exp_40_ram[37] = 8;
    exp_40_ram[38] = 133;
    exp_40_ram[39] = 131;
    exp_40_ram[40] = 148;
    exp_40_ram[41] = 22;
    exp_40_ram[42] = 134;
    exp_40_ram[43] = 246;
    exp_40_ram[44] = 7;
    exp_40_ram[45] = 120;
    exp_40_ram[46] = 7;
    exp_40_ram[47] = 55;
    exp_40_ram[48] = 23;
    exp_40_ram[49] = 85;
    exp_40_ram[50] = 134;
    exp_40_ram[51] = 198;
    exp_40_ram[52] = 5;
    exp_40_ram[53] = 135;
    exp_40_ram[54] = 6;
    exp_40_ram[55] = 12;
    exp_40_ram[56] = 149;
    exp_40_ram[57] = 215;
    exp_40_ram[58] = 24;
    exp_40_ram[59] = 101;
    exp_40_ram[60] = 147;
    exp_40_ram[61] = 88;
    exp_40_ram[62] = 214;
    exp_40_ram[63] = 22;
    exp_40_ram[64] = 86;
    exp_40_ram[65] = 87;
    exp_40_ram[66] = 247;
    exp_40_ram[67] = 133;
    exp_40_ram[68] = 5;
    exp_40_ram[69] = 23;
    exp_40_ram[70] = 103;
    exp_40_ram[71] = 254;
    exp_40_ram[72] = 135;
    exp_40_ram[73] = 133;
    exp_40_ram[74] = 232;
    exp_40_ram[75] = 246;
    exp_40_ram[76] = 133;
    exp_40_ram[77] = 135;
    exp_40_ram[78] = 135;
    exp_40_ram[79] = 247;
    exp_40_ram[80] = 19;
    exp_40_ram[81] = 83;
    exp_40_ram[82] = 215;
    exp_40_ram[83] = 23;
    exp_40_ram[84] = 99;
    exp_40_ram[85] = 6;
    exp_40_ram[86] = 134;
    exp_40_ram[87] = 124;
    exp_40_ram[88] = 3;
    exp_40_ram[89] = 134;
    exp_40_ram[90] = 102;
    exp_40_ram[91] = 116;
    exp_40_ram[92] = 134;
    exp_40_ram[93] = 21;
    exp_40_ram[94] = 101;
    exp_40_ram[95] = 5;
    exp_40_ram[96] = 0;
    exp_40_ram[97] = 5;
    exp_40_ram[98] = 7;
    exp_40_ram[99] = 108;
    exp_40_ram[100] = 7;
    exp_40_ram[101] = 240;
    exp_40_ram[102] = 22;
    exp_40_ram[103] = 7;
    exp_40_ram[104] = 88;
    exp_40_ram[105] = 7;
    exp_40_ram[106] = 112;
    exp_40_ram[107] = 7;
    exp_40_ram[108] = 116;
    exp_40_ram[109] = 5;
    exp_40_ram[110] = 87;
    exp_40_ram[111] = 134;
    exp_40_ram[112] = 199;
    exp_40_ram[113] = 6;
    exp_40_ram[114] = 7;
    exp_40_ram[115] = 6;
    exp_40_ram[116] = 22;
    exp_40_ram[117] = 135;
    exp_40_ram[118] = 5;
    exp_40_ram[119] = 88;
    exp_40_ram[120] = 22;
    exp_40_ram[121] = 86;
    exp_40_ram[122] = 87;
    exp_40_ram[123] = 246;
    exp_40_ram[124] = 215;
    exp_40_ram[125] = 150;
    exp_40_ram[126] = 231;
    exp_40_ram[127] = 14;
    exp_40_ram[128] = 133;
    exp_40_ram[129] = 126;
    exp_40_ram[130] = 7;
    exp_40_ram[131] = 133;
    exp_40_ram[132] = 104;
    exp_40_ram[133] = 118;
    exp_40_ram[134] = 133;
    exp_40_ram[135] = 7;
    exp_40_ram[136] = 7;
    exp_40_ram[137] = 119;
    exp_40_ram[138] = 19;
    exp_40_ram[139] = 83;
    exp_40_ram[140] = 87;
    exp_40_ram[141] = 151;
    exp_40_ram[142] = 227;
    exp_40_ram[143] = 6;
    exp_40_ram[144] = 6;
    exp_40_ram[145] = 124;
    exp_40_ram[146] = 3;
    exp_40_ram[147] = 6;
    exp_40_ram[148] = 102;
    exp_40_ram[149] = 116;
    exp_40_ram[150] = 6;
    exp_40_ram[151] = 21;
    exp_40_ram[152] = 101;
    exp_40_ram[153] = 128;
    exp_40_ram[154] = 7;
    exp_40_ram[155] = 5;
    exp_40_ram[156] = 100;
    exp_40_ram[157] = 5;
    exp_40_ram[158] = 240;
    exp_40_ram[159] = 24;
    exp_40_ram[160] = 213;
    exp_40_ram[161] = 147;
    exp_40_ram[162] = 151;
    exp_40_ram[163] = 215;
    exp_40_ram[164] = 88;
    exp_40_ram[165] = 102;
    exp_40_ram[166] = 119;
    exp_40_ram[167] = 23;
    exp_40_ram[168] = 215;
    exp_40_ram[169] = 85;
    exp_40_ram[170] = 85;
    exp_40_ram[171] = 23;
    exp_40_ram[172] = 103;
    exp_40_ram[173] = 134;
    exp_40_ram[174] = 5;
    exp_40_ram[175] = 126;
    exp_40_ram[176] = 7;
    exp_40_ram[177] = 5;
    exp_40_ram[178] = 104;
    exp_40_ram[179] = 118;
    exp_40_ram[180] = 5;
    exp_40_ram[181] = 7;
    exp_40_ram[182] = 6;
    exp_40_ram[183] = 247;
    exp_40_ram[184] = 22;
    exp_40_ram[185] = 86;
    exp_40_ram[186] = 214;
    exp_40_ram[187] = 23;
    exp_40_ram[188] = 133;
    exp_40_ram[189] = 103;
    exp_40_ram[190] = 135;
    exp_40_ram[191] = 254;
    exp_40_ram[192] = 135;
    exp_40_ram[193] = 135;
    exp_40_ram[194] = 232;
    exp_40_ram[195] = 246;
    exp_40_ram[196] = 135;
    exp_40_ram[197] = 135;
    exp_40_ram[198] = 149;
    exp_40_ram[199] = 135;
    exp_40_ram[200] = 229;
    exp_40_ram[201] = 240;
    exp_40_ram[202] = 230;
    exp_40_ram[203] = 7;
    exp_40_ram[204] = 244;
    exp_40_ram[205] = 7;
    exp_40_ram[206] = 53;
    exp_40_ram[207] = 149;
    exp_40_ram[208] = 23;
    exp_40_ram[209] = 213;
    exp_40_ram[210] = 7;
    exp_40_ram[211] = 7;
    exp_40_ram[212] = 71;
    exp_40_ram[213] = 5;
    exp_40_ram[214] = 7;
    exp_40_ram[215] = 5;
    exp_40_ram[216] = 22;
    exp_40_ram[217] = 5;
    exp_40_ram[218] = 238;
    exp_40_ram[219] = 181;
    exp_40_ram[220] = 69;
    exp_40_ram[221] = 240;
    exp_40_ram[222] = 7;
    exp_40_ram[223] = 5;
    exp_40_ram[224] = 224;
    exp_40_ram[225] = 5;
    exp_40_ram[226] = 240;
    exp_40_ram[227] = 88;
    exp_40_ram[228] = 150;
    exp_40_ram[229] = 104;
    exp_40_ram[230] = 222;
    exp_40_ram[231] = 94;
    exp_40_ram[232] = 118;
    exp_40_ram[233] = 151;
    exp_40_ram[234] = 215;
    exp_40_ram[235] = 19;
    exp_40_ram[236] = 102;
    exp_40_ram[237] = 23;
    exp_40_ram[238] = 215;
    exp_40_ram[239] = 87;
    exp_40_ram[240] = 94;
    exp_40_ram[241] = 150;
    exp_40_ram[242] = 231;
    exp_40_ram[243] = 143;
    exp_40_ram[244] = 5;
    exp_40_ram[245] = 126;
    exp_40_ram[246] = 7;
    exp_40_ram[247] = 5;
    exp_40_ram[248] = 104;
    exp_40_ram[249] = 118;
    exp_40_ram[250] = 5;
    exp_40_ram[251] = 7;
    exp_40_ram[252] = 7;
    exp_40_ram[253] = 118;
    exp_40_ram[254] = 87;
    exp_40_ram[255] = 150;
    exp_40_ram[256] = 142;
    exp_40_ram[257] = 23;
    exp_40_ram[258] = 215;
    exp_40_ram[259] = 231;
    exp_40_ram[260] = 6;
    exp_40_ram[261] = 254;
    exp_40_ram[262] = 135;
    exp_40_ram[263] = 6;
    exp_40_ram[264] = 232;
    exp_40_ram[265] = 246;
    exp_40_ram[266] = 6;
    exp_40_ram[267] = 135;
    exp_40_ram[268] = 21;
    exp_40_ram[269] = 14;
    exp_40_ram[270] = 101;
    exp_40_ram[271] = 134;
    exp_40_ram[272] = 120;
    exp_40_ram[273] = 86;
    exp_40_ram[274] = 118;
    exp_40_ram[275] = 83;
    exp_40_ram[276] = 135;
    exp_40_ram[277] = 14;
    exp_40_ram[278] = 6;
    exp_40_ram[279] = 87;
    exp_40_ram[280] = 8;
    exp_40_ram[281] = 8;
    exp_40_ram[282] = 7;
    exp_40_ram[283] = 6;
    exp_40_ram[284] = 116;
    exp_40_ram[285] = 6;
    exp_40_ram[286] = 86;
    exp_40_ram[287] = 134;
    exp_40_ram[288] = 230;
    exp_40_ram[289] = 156;
    exp_40_ram[290] = 7;
    exp_40_ram[291] = 135;
    exp_40_ram[292] = 119;
    exp_40_ram[293] = 23;
    exp_40_ram[294] = 126;
    exp_40_ram[295] = 152;
    exp_40_ram[296] = 7;
    exp_40_ram[297] = 5;
    exp_40_ram[298] = 254;
    exp_40_ram[299] = 5;
    exp_40_ram[300] = 240;
    exp_40_ram[301] = 5;
    exp_40_ram[302] = 5;
    exp_40_ram[303] = 240;
    exp_40_ram[304] = 7;
    exp_40_ram[305] = 7;
    exp_40_ram[306] = 216;
    exp_40_ram[307] = 120;
    exp_40_ram[308] = 7;
    exp_40_ram[309] = 3;
    exp_40_ram[310] = 120;
    exp_40_ram[311] = 213;
    exp_40_ram[312] = 14;
    exp_40_ram[313] = 213;
    exp_40_ram[314] = 119;
    exp_40_ram[315] = 14;
    exp_40_ram[316] = 245;
    exp_40_ram[317] = 214;
    exp_40_ram[318] = 26;
    exp_40_ram[319] = 238;
    exp_40_ram[320] = 138;
    exp_40_ram[321] = 5;
    exp_40_ram[322] = 128;
    exp_40_ram[323] = 150;
    exp_40_ram[324] = 110;
    exp_40_ram[325] = 152;
    exp_40_ram[326] = 16;
    exp_40_ram[327] = 231;
    exp_40_ram[328] = 183;
    exp_40_ram[329] = 150;
    exp_40_ram[330] = 102;
    exp_40_ram[331] = 12;
    exp_40_ram[332] = 156;
    exp_40_ram[333] = 20;
    exp_40_ram[334] = 208;
    exp_40_ram[335] = 0;
    exp_40_ram[336] = 5;
    exp_40_ram[337] = 128;
    exp_40_ram[338] = 5;
    exp_40_ram[339] = 138;
    exp_40_ram[340] = 133;
    exp_40_ram[341] = 128;
    exp_40_ram[342] = 86;
    exp_40_ram[343] = 2;
    exp_40_ram[344] = 128;
    exp_40_ram[345] = 108;
    exp_40_ram[346] = 146;
    exp_40_ram[347] = 104;
    exp_40_ram[348] = 102;
    exp_40_ram[349] = 5;
    exp_40_ram[350] = 128;
    exp_40_ram[351] = 5;
    exp_40_ram[352] = 128;
    exp_40_ram[353] = 152;
    exp_40_ram[354] = 240;
    exp_40_ram[355] = 232;
    exp_40_ram[356] = 240;
    exp_40_ram[357] = 142;
    exp_40_ram[358] = 158;
    exp_40_ram[359] = 7;
    exp_40_ram[360] = 240;
    exp_40_ram[361] = 1;
    exp_40_ram[362] = 36;
    exp_40_ram[363] = 38;
    exp_40_ram[364] = 4;
    exp_40_ram[365] = 2;
    exp_40_ram[366] = 0;
    exp_40_ram[367] = 7;
    exp_40_ram[368] = 7;
    exp_40_ram[369] = 7;
    exp_40_ram[370] = 192;
    exp_40_ram[371] = 7;
    exp_40_ram[372] = 135;
    exp_40_ram[373] = 5;
    exp_40_ram[374] = 87;
    exp_40_ram[375] = 20;
    exp_40_ram[376] = 32;
    exp_40_ram[377] = 5;
    exp_40_ram[378] = 151;
    exp_40_ram[379] = 36;
    exp_40_ram[380] = 23;
    exp_40_ram[381] = 215;
    exp_40_ram[382] = 102;
    exp_40_ram[383] = 133;
    exp_40_ram[384] = 1;
    exp_40_ram[385] = 128;
    exp_40_ram[386] = 7;
    exp_40_ram[387] = 23;
    exp_40_ram[388] = 4;
    exp_40_ram[389] = 240;
    exp_40_ram[390] = 7;
    exp_40_ram[391] = 7;
    exp_40_ram[392] = 240;
    exp_40_ram[393] = 1;
    exp_40_ram[394] = 46;
    exp_40_ram[395] = 44;
    exp_40_ram[396] = 42;
    exp_40_ram[397] = 40;
    exp_40_ram[398] = 38;
    exp_40_ram[399] = 36;
    exp_40_ram[400] = 103;
    exp_40_ram[401] = 140;
    exp_40_ram[402] = 4;
    exp_40_ram[403] = 137;
    exp_40_ram[404] = 132;
    exp_40_ram[405] = 132;
    exp_40_ram[406] = 133;
    exp_40_ram[407] = 0;
    exp_40_ram[408] = 9;
    exp_40_ram[409] = 10;
    exp_40_ram[410] = 10;
    exp_40_ram[411] = 7;
    exp_40_ram[412] = 196;
    exp_40_ram[413] = 7;
    exp_40_ram[414] = 7;
    exp_40_ram[415] = 84;
    exp_40_ram[416] = 7;
    exp_40_ram[417] = 66;
    exp_40_ram[418] = 4;
    exp_40_ram[419] = 135;
    exp_40_ram[420] = 132;
    exp_40_ram[421] = 84;
    exp_40_ram[422] = 21;
    exp_40_ram[423] = 228;
    exp_40_ram[424] = 23;
    exp_40_ram[425] = 32;
    exp_40_ram[426] = 36;
    exp_40_ram[427] = 149;
    exp_40_ram[428] = 26;
    exp_40_ram[429] = 213;
    exp_40_ram[430] = 103;
    exp_40_ram[431] = 36;
    exp_40_ram[432] = 41;
    exp_40_ram[433] = 41;
    exp_40_ram[434] = 42;
    exp_40_ram[435] = 133;
    exp_40_ram[436] = 5;
    exp_40_ram[437] = 1;
    exp_40_ram[438] = 128;
    exp_40_ram[439] = 0;
    exp_40_ram[440] = 9;
    exp_40_ram[441] = 240;
    exp_40_ram[442] = 133;
    exp_40_ram[443] = 20;
    exp_40_ram[444] = 7;
    exp_40_ram[445] = 240;
    exp_40_ram[446] = 7;
    exp_40_ram[447] = 220;
    exp_40_ram[448] = 134;
    exp_40_ram[449] = 5;
    exp_40_ram[450] = 5;
    exp_40_ram[451] = 0;
    exp_40_ram[452] = 101;
    exp_40_ram[453] = 6;
    exp_40_ram[454] = 52;
    exp_40_ram[455] = 5;
    exp_40_ram[456] = 5;
    exp_40_ram[457] = 6;
    exp_40_ram[458] = 0;
    exp_40_ram[459] = 228;
    exp_40_ram[460] = 137;
    exp_40_ram[461] = 7;
    exp_40_ram[462] = 7;
    exp_40_ram[463] = 5;
    exp_40_ram[464] = 84;
    exp_40_ram[465] = 7;
    exp_40_ram[466] = 66;
    exp_40_ram[467] = 135;
    exp_40_ram[468] = 21;
    exp_40_ram[469] = 9;
    exp_40_ram[470] = 9;
    exp_40_ram[471] = 89;
    exp_40_ram[472] = 101;
    exp_40_ram[473] = 23;
    exp_40_ram[474] = 7;
    exp_40_ram[475] = 7;
    exp_40_ram[476] = 245;
    exp_40_ram[477] = 247;
    exp_40_ram[478] = 0;
    exp_40_ram[479] = 247;
    exp_40_ram[480] = 6;
    exp_40_ram[481] = 10;
    exp_40_ram[482] = 135;
    exp_40_ram[483] = 55;
    exp_40_ram[484] = 133;
    exp_40_ram[485] = 7;
    exp_40_ram[486] = 7;
    exp_40_ram[487] = 247;
    exp_40_ram[488] = 12;
    exp_40_ram[489] = 7;
    exp_40_ram[490] = 7;
    exp_40_ram[491] = 10;
    exp_40_ram[492] = 245;
    exp_40_ram[493] = 10;
    exp_40_ram[494] = 215;
    exp_40_ram[495] = 149;
    exp_40_ram[496] = 103;
    exp_40_ram[497] = 212;
    exp_40_ram[498] = 240;
    exp_40_ram[499] = 133;
    exp_40_ram[500] = 21;
    exp_40_ram[501] = 7;
    exp_40_ram[502] = 240;
    exp_40_ram[503] = 4;
    exp_40_ram[504] = 7;
    exp_40_ram[505] = 10;
    exp_40_ram[506] = 240;
    exp_40_ram[507] = 6;
    exp_40_ram[508] = 5;
    exp_40_ram[509] = 246;
    exp_40_ram[510] = 132;
    exp_40_ram[511] = 5;
    exp_40_ram[512] = 213;
    exp_40_ram[513] = 22;
    exp_40_ram[514] = 150;
    exp_40_ram[515] = 128;
    exp_40_ram[516] = 64;
    exp_40_ram[517] = 198;
    exp_40_ram[518] = 134;
    exp_40_ram[519] = 5;
    exp_40_ram[520] = 5;
    exp_40_ram[521] = 12;
    exp_40_ram[522] = 6;
    exp_40_ram[523] = 122;
    exp_40_ram[524] = 88;
    exp_40_ram[525] = 22;
    exp_40_ram[526] = 150;
    exp_40_ram[527] = 106;
    exp_40_ram[528] = 5;
    exp_40_ram[529] = 230;
    exp_40_ram[530] = 133;
    exp_40_ram[531] = 101;
    exp_40_ram[532] = 214;
    exp_40_ram[533] = 86;
    exp_40_ram[534] = 150;
    exp_40_ram[535] = 128;
    exp_40_ram[536] = 130;
    exp_40_ram[537] = 240;
    exp_40_ram[538] = 133;
    exp_40_ram[539] = 128;
    exp_40_ram[540] = 5;
    exp_40_ram[541] = 72;
    exp_40_ram[542] = 5;
    exp_40_ram[543] = 240;
    exp_40_ram[544] = 5;
    exp_40_ram[545] = 130;
    exp_40_ram[546] = 240;
    exp_40_ram[547] = 5;
    exp_40_ram[548] = 128;
    exp_40_ram[549] = 130;
    exp_40_ram[550] = 202;
    exp_40_ram[551] = 76;
    exp_40_ram[552] = 240;
    exp_40_ram[553] = 133;
    exp_40_ram[554] = 128;
    exp_40_ram[555] = 5;
    exp_40_ram[556] = 88;
    exp_40_ram[557] = 5;
    exp_40_ram[558] = 240;
    exp_40_ram[559] = 5;
    exp_40_ram[560] = 128;
    exp_40_ram[561] = 0;
    exp_40_ram[562] = 7;
    exp_40_ram[563] = 135;
    exp_40_ram[564] = 76;
    exp_40_ram[565] = 5;
    exp_40_ram[566] = 7;
    exp_40_ram[567] = 213;
    exp_40_ram[568] = 5;
    exp_40_ram[569] = 128;
    exp_40_ram[570] = 215;
    exp_40_ram[571] = 85;
    exp_40_ram[572] = 149;
    exp_40_ram[573] = 101;
    exp_40_ram[574] = 240;
    exp_40_ram[575] = 0;
    exp_40_ram[576] = 7;
    exp_40_ram[577] = 135;
    exp_40_ram[578] = 76;
    exp_40_ram[579] = 5;
    exp_40_ram[580] = 7;
    exp_40_ram[581] = 21;
    exp_40_ram[582] = 5;
    exp_40_ram[583] = 128;
    exp_40_ram[584] = 23;
    exp_40_ram[585] = 149;
    exp_40_ram[586] = 85;
    exp_40_ram[587] = 229;
    exp_40_ram[588] = 240;
    exp_40_ram[589] = 7;
    exp_40_ram[590] = 122;
    exp_40_ram[591] = 7;
    exp_40_ram[592] = 183;
    exp_40_ram[593] = 151;
    exp_40_ram[594] = 23;
    exp_40_ram[595] = 6;
    exp_40_ram[596] = 134;
    exp_40_ram[597] = 85;
    exp_40_ram[598] = 7;
    exp_40_ram[599] = 133;
    exp_40_ram[600] = 69;
    exp_40_ram[601] = 133;
    exp_40_ram[602] = 128;
    exp_40_ram[603] = 7;
    exp_40_ram[604] = 7;
    exp_40_ram[605] = 106;
    exp_40_ram[606] = 7;
    exp_40_ram[607] = 240;
    exp_40_ram[608] = 116;
    exp_40_ram[609] = 112;
    exp_40_ram[610] = 0;
    exp_40_ram[611] = 97;
    exp_40_ram[612] = 0;
    exp_40_ram[613] = 105;
    exp_40_ram[614] = 46;
    exp_40_ram[615] = 104;
    exp_40_ram[616] = 101;
    exp_40_ram[617] = 55;
    exp_40_ram[618] = 58;
    exp_40_ram[619] = 48;
    exp_40_ram[620] = 48;
    exp_40_ram[621] = 0;
    exp_40_ram[622] = 32;
    exp_40_ram[623] = 108;
    exp_40_ram[624] = 104;
    exp_40_ram[625] = 101;
    exp_40_ram[626] = 55;
    exp_40_ram[627] = 58;
    exp_40_ram[628] = 48;
    exp_40_ram[629] = 48;
    exp_40_ram[630] = 0;
    exp_40_ram[631] = 32;
    exp_40_ram[632] = 108;
    exp_40_ram[633] = 32;
    exp_40_ram[634] = 108;
    exp_40_ram[635] = 32;
    exp_40_ram[636] = 108;
    exp_40_ram[637] = 32;
    exp_40_ram[638] = 108;
    exp_40_ram[639] = 32;
    exp_40_ram[640] = 108;
    exp_40_ram[641] = 32;
    exp_40_ram[642] = 108;
    exp_40_ram[643] = 32;
    exp_40_ram[644] = 108;
    exp_40_ram[645] = 32;
    exp_40_ram[646] = 108;
    exp_40_ram[647] = 104;
    exp_40_ram[648] = 101;
    exp_40_ram[649] = 55;
    exp_40_ram[650] = 58;
    exp_40_ram[651] = 48;
    exp_40_ram[652] = 48;
    exp_40_ram[653] = 0;
    exp_40_ram[654] = 48;
    exp_40_ram[655] = 105;
    exp_40_ram[656] = 49;
    exp_40_ram[657] = 105;
    exp_40_ram[658] = 50;
    exp_40_ram[659] = 105;
    exp_40_ram[660] = 97;
    exp_40_ram[661] = 0;
    exp_40_ram[662] = 1;
    exp_40_ram[663] = 3;
    exp_40_ram[664] = 4;
    exp_40_ram[665] = 4;
    exp_40_ram[666] = 5;
    exp_40_ram[667] = 5;
    exp_40_ram[668] = 5;
    exp_40_ram[669] = 5;
    exp_40_ram[670] = 6;
    exp_40_ram[671] = 6;
    exp_40_ram[672] = 6;
    exp_40_ram[673] = 6;
    exp_40_ram[674] = 6;
    exp_40_ram[675] = 6;
    exp_40_ram[676] = 6;
    exp_40_ram[677] = 6;
    exp_40_ram[678] = 7;
    exp_40_ram[679] = 7;
    exp_40_ram[680] = 7;
    exp_40_ram[681] = 7;
    exp_40_ram[682] = 7;
    exp_40_ram[683] = 7;
    exp_40_ram[684] = 7;
    exp_40_ram[685] = 7;
    exp_40_ram[686] = 7;
    exp_40_ram[687] = 7;
    exp_40_ram[688] = 7;
    exp_40_ram[689] = 7;
    exp_40_ram[690] = 7;
    exp_40_ram[691] = 7;
    exp_40_ram[692] = 7;
    exp_40_ram[693] = 7;
    exp_40_ram[694] = 8;
    exp_40_ram[695] = 8;
    exp_40_ram[696] = 8;
    exp_40_ram[697] = 8;
    exp_40_ram[698] = 8;
    exp_40_ram[699] = 8;
    exp_40_ram[700] = 8;
    exp_40_ram[701] = 8;
    exp_40_ram[702] = 8;
    exp_40_ram[703] = 8;
    exp_40_ram[704] = 8;
    exp_40_ram[705] = 8;
    exp_40_ram[706] = 8;
    exp_40_ram[707] = 8;
    exp_40_ram[708] = 8;
    exp_40_ram[709] = 8;
    exp_40_ram[710] = 8;
    exp_40_ram[711] = 8;
    exp_40_ram[712] = 8;
    exp_40_ram[713] = 8;
    exp_40_ram[714] = 8;
    exp_40_ram[715] = 8;
    exp_40_ram[716] = 8;
    exp_40_ram[717] = 8;
    exp_40_ram[718] = 8;
    exp_40_ram[719] = 8;
    exp_40_ram[720] = 8;
    exp_40_ram[721] = 8;
    exp_40_ram[722] = 8;
    exp_40_ram[723] = 8;
    exp_40_ram[724] = 8;
    exp_40_ram[725] = 8;
    exp_40_ram[726] = 7;
    exp_40_ram[727] = 5;
    exp_40_ram[728] = 135;
    exp_40_ram[729] = 71;
    exp_40_ram[730] = 20;
    exp_40_ram[731] = 128;
    exp_40_ram[732] = 5;
    exp_40_ram[733] = 160;
    exp_40_ram[734] = 240;
    exp_40_ram[735] = 1;
    exp_40_ram[736] = 39;
    exp_40_ram[737] = 36;
    exp_40_ram[738] = 164;
    exp_40_ram[739] = 38;
    exp_40_ram[740] = 5;
    exp_40_ram[741] = 240;
    exp_40_ram[742] = 7;
    exp_40_ram[743] = 32;
    exp_40_ram[744] = 32;
    exp_40_ram[745] = 36;
    exp_40_ram[746] = 5;
    exp_40_ram[747] = 1;
    exp_40_ram[748] = 128;
    exp_40_ram[749] = 103;
    exp_40_ram[750] = 247;
    exp_40_ram[751] = 6;
    exp_40_ram[752] = 152;
    exp_40_ram[753] = 135;
    exp_40_ram[754] = 131;
    exp_40_ram[755] = 8;
    exp_40_ram[756] = 0;
    exp_40_ram[757] = 40;
    exp_40_ram[758] = 7;
    exp_40_ram[759] = 134;
    exp_40_ram[760] = 168;
    exp_40_ram[761] = 40;
    exp_40_ram[762] = 170;
    exp_40_ram[763] = 40;
    exp_40_ram[764] = 172;
    exp_40_ram[765] = 40;
    exp_40_ram[766] = 174;
    exp_40_ram[767] = 8;
    exp_40_ram[768] = 106;
    exp_40_ram[769] = 119;
    exp_40_ram[770] = 118;
    exp_40_ram[771] = 6;
    exp_40_ram[772] = 133;
    exp_40_ram[773] = 6;
    exp_40_ram[774] = 8;
    exp_40_ram[775] = 96;
    exp_40_ram[776] = 118;
    exp_40_ram[777] = 119;
    exp_40_ram[778] = 134;
    exp_40_ram[779] = 133;
    exp_40_ram[780] = 7;
    exp_40_ram[781] = 16;
    exp_40_ram[782] = 128;
    exp_40_ram[783] = 136;
    exp_40_ram[784] = 40;
    exp_40_ram[785] = 136;
    exp_40_ram[786] = 135;
    exp_40_ram[787] = 32;
    exp_40_ram[788] = 240;
    exp_40_ram[789] = 135;
    exp_40_ram[790] = 72;
    exp_40_ram[791] = 135;
    exp_40_ram[792] = 135;
    exp_40_ram[793] = 0;
    exp_40_ram[794] = 240;
    exp_40_ram[795] = 103;
    exp_40_ram[796] = 247;
    exp_40_ram[797] = 144;
    exp_40_ram[798] = 6;
    exp_40_ram[799] = 134;
    exp_40_ram[800] = 134;
    exp_40_ram[801] = 6;
    exp_40_ram[802] = 167;
    exp_40_ram[803] = 39;
    exp_40_ram[804] = 142;
    exp_40_ram[805] = 71;
    exp_40_ram[806] = 199;
    exp_40_ram[807] = 132;
    exp_40_ram[808] = 134;
    exp_40_ram[809] = 133;
    exp_40_ram[810] = 128;
    exp_40_ram[811] = 135;
    exp_40_ram[812] = 199;
    exp_40_ram[813] = 119;
    exp_40_ram[814] = 247;
    exp_40_ram[815] = 142;
    exp_40_ram[816] = 5;
    exp_40_ram[817] = 133;
    exp_40_ram[818] = 240;
    exp_40_ram[819] = 5;
    exp_40_ram[820] = 133;
    exp_40_ram[821] = 240;
    exp_40_ram[822] = 5;
    exp_40_ram[823] = 128;
    exp_40_ram[824] = 119;
    exp_40_ram[825] = 148;
    exp_40_ram[826] = 1;
    exp_40_ram[827] = 5;
    exp_40_ram[828] = 36;
    exp_40_ram[829] = 38;
    exp_40_ram[830] = 4;
    exp_40_ram[831] = 240;
    exp_40_ram[832] = 7;
    exp_40_ram[833] = 26;
    exp_40_ram[834] = 5;
    exp_40_ram[835] = 5;
    exp_40_ram[836] = 240;
    exp_40_ram[837] = 55;
    exp_40_ram[838] = 32;
    exp_40_ram[839] = 36;
    exp_40_ram[840] = 133;
    exp_40_ram[841] = 1;
    exp_40_ram[842] = 128;
    exp_40_ram[843] = 7;
    exp_40_ram[844] = 133;
    exp_40_ram[845] = 128;
    exp_40_ram[846] = 135;
    exp_40_ram[847] = 247;
    exp_40_ram[848] = 130;
    exp_40_ram[849] = 247;
    exp_40_ram[850] = 6;
    exp_40_ram[851] = 7;
    exp_40_ram[852] = 12;
    exp_40_ram[853] = 7;
    exp_40_ram[854] = 7;
    exp_40_ram[855] = 150;
    exp_40_ram[856] = 1;
    exp_40_ram[857] = 38;
    exp_40_ram[858] = 240;
    exp_40_ram[859] = 32;
    exp_40_ram[860] = 55;
    exp_40_ram[861] = 135;
    exp_40_ram[862] = 133;
    exp_40_ram[863] = 1;
    exp_40_ram[864] = 128;
    exp_40_ram[865] = 7;
    exp_40_ram[866] = 133;
    exp_40_ram[867] = 128;
    exp_40_ram[868] = 7;
    exp_40_ram[869] = 166;
    exp_40_ram[870] = 166;
    exp_40_ram[871] = 165;
    exp_40_ram[872] = 5;
    exp_40_ram[873] = 167;
    exp_40_ram[874] = 229;
    exp_40_ram[875] = 128;
    exp_40_ram[876] = 7;
    exp_40_ram[877] = 5;
    exp_40_ram[878] = 183;
    exp_40_ram[879] = 133;
    exp_40_ram[880] = 1;
    exp_40_ram[881] = 133;
    exp_40_ram[882] = 38;
    exp_40_ram[883] = 240;
    exp_40_ram[884] = 32;
    exp_40_ram[885] = 1;
    exp_40_ram[886] = 128;
    exp_40_ram[887] = 1;
    exp_40_ram[888] = 34;
    exp_40_ram[889] = 42;
    exp_40_ram[890] = 42;
    exp_40_ram[891] = 84;
    exp_40_ram[892] = 44;
    exp_40_ram[893] = 40;
    exp_40_ram[894] = 38;
    exp_40_ram[895] = 36;
    exp_40_ram[896] = 46;
    exp_40_ram[897] = 32;
    exp_40_ram[898] = 10;
    exp_40_ram[899] = 4;
    exp_40_ram[900] = 9;
    exp_40_ram[901] = 9;
    exp_40_ram[902] = 138;
    exp_40_ram[903] = 132;
    exp_40_ram[904] = 146;
    exp_40_ram[905] = 43;
    exp_40_ram[906] = 90;
    exp_40_ram[907] = 4;
    exp_40_ram[908] = 138;
    exp_40_ram[909] = 0;
    exp_40_ram[910] = 133;
    exp_40_ram[911] = 5;
    exp_40_ram[912] = 240;
    exp_40_ram[913] = 133;
    exp_40_ram[914] = 240;
    exp_40_ram[915] = 5;
    exp_40_ram[916] = 55;
    exp_40_ram[917] = 137;
    exp_40_ram[918] = 9;
    exp_40_ram[919] = 132;
    exp_40_ram[920] = 240;
    exp_40_ram[921] = 5;
    exp_40_ram[922] = 240;
    exp_40_ram[923] = 53;
    exp_40_ram[924] = 133;
    exp_40_ram[925] = 5;
    exp_40_ram[926] = 240;
    exp_40_ram[927] = 5;
    exp_40_ram[928] = 55;
    exp_40_ram[929] = 137;
    exp_40_ram[930] = 9;
    exp_40_ram[931] = 4;
    exp_40_ram[932] = 240;
    exp_40_ram[933] = 39;
    exp_40_ram[934] = 38;
    exp_40_ram[935] = 36;
    exp_40_ram[936] = 23;
    exp_40_ram[937] = 135;
    exp_40_ram[938] = 151;
    exp_40_ram[939] = 135;
    exp_40_ram[940] = 23;
    exp_40_ram[941] = 7;
    exp_40_ram[942] = 151;
    exp_40_ram[943] = 23;
    exp_40_ram[944] = 37;
    exp_40_ram[945] = 86;
    exp_40_ram[946] = 214;
    exp_40_ram[947] = 135;
    exp_40_ram[948] = 134;
    exp_40_ram[949] = 55;
    exp_40_ram[950] = 135;
    exp_40_ram[951] = 85;
    exp_40_ram[952] = 214;
    exp_40_ram[953] = 4;
    exp_40_ram[954] = 183;
    exp_40_ram[955] = 135;
    exp_40_ram[956] = 133;
    exp_40_ram[957] = 5;
    exp_40_ram[958] = 4;
    exp_40_ram[959] = 240;
    exp_40_ram[960] = 133;
    exp_40_ram[961] = 87;
    exp_40_ram[962] = 180;
    exp_40_ram[963] = 7;
    exp_40_ram[964] = 133;
    exp_40_ram[965] = 132;
    exp_40_ram[966] = 4;
    exp_40_ram[967] = 53;
    exp_40_ram[968] = 32;
    exp_40_ram[969] = 133;
    exp_40_ram[970] = 36;
    exp_40_ram[971] = 36;
    exp_40_ram[972] = 41;
    exp_40_ram[973] = 41;
    exp_40_ram[974] = 42;
    exp_40_ram[975] = 42;
    exp_40_ram[976] = 43;
    exp_40_ram[977] = 1;
    exp_40_ram[978] = 128;
    exp_40_ram[979] = 1;
    exp_40_ram[980] = 38;
    exp_40_ram[981] = 36;
    exp_40_ram[982] = 4;
    exp_40_ram[983] = 240;
    exp_40_ram[984] = 39;
    exp_40_ram[985] = 166;
    exp_40_ram[986] = 6;
    exp_40_ram[987] = 240;
    exp_40_ram[988] = 39;
    exp_40_ram[989] = 167;
    exp_40_ram[990] = 5;
    exp_40_ram[991] = 6;
    exp_40_ram[992] = 32;
    exp_40_ram[993] = 34;
    exp_40_ram[994] = 32;
    exp_40_ram[995] = 36;
    exp_40_ram[996] = 5;
    exp_40_ram[997] = 1;
    exp_40_ram[998] = 128;
    exp_40_ram[999] = 1;
    exp_40_ram[1000] = 38;
    exp_40_ram[1001] = 36;
    exp_40_ram[1002] = 34;
    exp_40_ram[1003] = 32;
    exp_40_ram[1004] = 4;
    exp_40_ram[1005] = 132;
    exp_40_ram[1006] = 240;
    exp_40_ram[1007] = 39;
    exp_40_ram[1008] = 166;
    exp_40_ram[1009] = 6;
    exp_40_ram[1010] = 41;
    exp_40_ram[1011] = 240;
    exp_40_ram[1012] = 133;
    exp_40_ram[1013] = 180;
    exp_40_ram[1014] = 4;
    exp_40_ram[1015] = 9;
    exp_40_ram[1016] = 4;
    exp_40_ram[1017] = 34;
    exp_40_ram[1018] = 32;
    exp_40_ram[1019] = 36;
    exp_40_ram[1020] = 32;
    exp_40_ram[1021] = 36;
    exp_40_ram[1022] = 41;
    exp_40_ram[1023] = 1;
    exp_40_ram[1024] = 128;
    exp_40_ram[1025] = 1;
    exp_40_ram[1026] = 37;
    exp_40_ram[1027] = 34;
    exp_40_ram[1028] = 6;
    exp_40_ram[1029] = 4;
    exp_40_ram[1030] = 133;
    exp_40_ram[1031] = 5;
    exp_40_ram[1032] = 38;
    exp_40_ram[1033] = 36;
    exp_40_ram[1034] = 32;
    exp_40_ram[1035] = 46;
    exp_40_ram[1036] = 44;
    exp_40_ram[1037] = 240;
    exp_40_ram[1038] = 37;
    exp_40_ram[1039] = 6;
    exp_40_ram[1040] = 133;
    exp_40_ram[1041] = 5;
    exp_40_ram[1042] = 240;
    exp_40_ram[1043] = 167;
    exp_40_ram[1044] = 41;
    exp_40_ram[1045] = 132;
    exp_40_ram[1046] = 149;
    exp_40_ram[1047] = 133;
    exp_40_ram[1048] = 7;
    exp_40_ram[1049] = 9;
    exp_40_ram[1050] = 133;
    exp_40_ram[1051] = 6;
    exp_40_ram[1052] = 133;
    exp_40_ram[1053] = 240;
    exp_40_ram[1054] = 1;
    exp_40_ram[1055] = 167;
    exp_40_ram[1056] = 6;
    exp_40_ram[1057] = 5;
    exp_40_ram[1058] = 149;
    exp_40_ram[1059] = 133;
    exp_40_ram[1060] = 7;
    exp_40_ram[1061] = 133;
    exp_40_ram[1062] = 240;
    exp_40_ram[1063] = 3;
    exp_40_ram[1064] = 165;
    exp_40_ram[1065] = 5;
    exp_40_ram[1066] = 10;
    exp_40_ram[1067] = 0;
    exp_40_ram[1068] = 36;
    exp_40_ram[1069] = 39;
    exp_40_ram[1070] = 38;
    exp_40_ram[1071] = 5;
    exp_40_ram[1072] = 135;
    exp_40_ram[1073] = 4;
    exp_40_ram[1074] = 39;
    exp_40_ram[1075] = 5;
    exp_40_ram[1076] = 135;
    exp_40_ram[1077] = 4;
    exp_40_ram[1078] = 165;
    exp_40_ram[1079] = 0;
    exp_40_ram[1080] = 36;
    exp_40_ram[1081] = 39;
    exp_40_ram[1082] = 38;
    exp_40_ram[1083] = 6;
    exp_40_ram[1084] = 135;
    exp_40_ram[1085] = 5;
    exp_40_ram[1086] = 39;
    exp_40_ram[1087] = 5;
    exp_40_ram[1088] = 135;
    exp_40_ram[1089] = 6;
    exp_40_ram[1090] = 165;
    exp_40_ram[1091] = 0;
    exp_40_ram[1092] = 36;
    exp_40_ram[1093] = 39;
    exp_40_ram[1094] = 38;
    exp_40_ram[1095] = 8;
    exp_40_ram[1096] = 135;
    exp_40_ram[1097] = 7;
    exp_40_ram[1098] = 39;
    exp_40_ram[1099] = 5;
    exp_40_ram[1100] = 135;
    exp_40_ram[1101] = 7;
    exp_40_ram[1102] = 165;
    exp_40_ram[1103] = 0;
    exp_40_ram[1104] = 36;
    exp_40_ram[1105] = 39;
    exp_40_ram[1106] = 38;
    exp_40_ram[1107] = 9;
    exp_40_ram[1108] = 135;
    exp_40_ram[1109] = 8;
    exp_40_ram[1110] = 39;
    exp_40_ram[1111] = 5;
    exp_40_ram[1112] = 135;
    exp_40_ram[1113] = 9;
    exp_40_ram[1114] = 165;
    exp_40_ram[1115] = 5;
    exp_40_ram[1116] = 0;
    exp_40_ram[1117] = 36;
    exp_40_ram[1118] = 38;
    exp_40_ram[1119] = 39;
    exp_40_ram[1120] = 37;
    exp_40_ram[1121] = 5;
    exp_40_ram[1122] = 135;
    exp_40_ram[1123] = 10;
    exp_40_ram[1124] = 0;
    exp_40_ram[1125] = 36;
    exp_40_ram[1126] = 38;
    exp_40_ram[1127] = 39;
    exp_40_ram[1128] = 37;
    exp_40_ram[1129] = 5;
    exp_40_ram[1130] = 135;
    exp_40_ram[1131] = 10;
    exp_40_ram[1132] = 0;
    exp_40_ram[1133] = 36;
    exp_40_ram[1134] = 39;
    exp_40_ram[1135] = 38;
    exp_40_ram[1136] = 32;
    exp_40_ram[1137] = 135;
    exp_40_ram[1138] = 11;
    exp_40_ram[1139] = 39;
    exp_40_ram[1140] = 36;
    exp_40_ram[1141] = 41;
    exp_40_ram[1142] = 135;
    exp_40_ram[1143] = 11;
    exp_40_ram[1144] = 7;
    exp_40_ram[1145] = 28;
    exp_40_ram[1146] = 36;
    exp_40_ram[1147] = 42;
    exp_40_ram[1148] = 133;
    exp_40_ram[1149] = 41;
    exp_40_ram[1150] = 1;
    exp_40_ram[1151] = 128;
    exp_40_ram[1152] = 1;
    exp_40_ram[1153] = 32;
    exp_40_ram[1154] = 91;
    exp_40_ram[1155] = 44;
    exp_40_ram[1156] = 42;
    exp_40_ram[1157] = 40;
    exp_40_ram[1158] = 38;
    exp_40_ram[1159] = 34;
    exp_40_ram[1160] = 46;
    exp_40_ram[1161] = 36;
    exp_40_ram[1162] = 46;
    exp_40_ram[1163] = 44;
    exp_40_ram[1164] = 42;
    exp_40_ram[1165] = 4;
    exp_40_ram[1166] = 132;
    exp_40_ram[1167] = 9;
    exp_40_ram[1168] = 9;
    exp_40_ram[1169] = 10;
    exp_40_ram[1170] = 11;
    exp_40_ram[1171] = 133;
    exp_40_ram[1172] = 240;
    exp_40_ram[1173] = 58;
    exp_40_ram[1174] = 10;
    exp_40_ram[1175] = 5;
    exp_40_ram[1176] = 5;
    exp_40_ram[1177] = 240;
    exp_40_ram[1178] = 135;
    exp_40_ram[1179] = 20;
    exp_40_ram[1180] = 224;
    exp_40_ram[1181] = 133;
    exp_40_ram[1182] = 183;
    exp_40_ram[1183] = 138;
    exp_40_ram[1184] = 4;
    exp_40_ram[1185] = 9;
    exp_40_ram[1186] = 137;
    exp_40_ram[1187] = 240;
    exp_40_ram[1188] = 92;
    exp_40_ram[1189] = 12;
    exp_40_ram[1190] = 10;
    exp_40_ram[1191] = 12;
    exp_40_ram[1192] = 133;
    exp_40_ram[1193] = 133;
    exp_40_ram[1194] = 240;
    exp_40_ram[1195] = 5;
    exp_40_ram[1196] = 139;
    exp_40_ram[1197] = 11;
    exp_40_ram[1198] = 140;
    exp_40_ram[1199] = 240;
    exp_40_ram[1200] = 20;
    exp_40_ram[1201] = 224;
    exp_40_ram[1202] = 133;
    exp_40_ram[1203] = 183;
    exp_40_ram[1204] = 138;
    exp_40_ram[1205] = 10;
    exp_40_ram[1206] = 4;
    exp_40_ram[1207] = 9;
    exp_40_ram[1208] = 240;
    exp_40_ram[1209] = 85;
    exp_40_ram[1210] = 133;
    exp_40_ram[1211] = 133;
    exp_40_ram[1212] = 0;
    exp_40_ram[1213] = 38;
    exp_40_ram[1214] = 4;
    exp_40_ram[1215] = 36;
    exp_40_ram[1216] = 10;
    exp_40_ram[1217] = 37;
    exp_40_ram[1218] = 21;
    exp_40_ram[1219] = 133;
    exp_40_ram[1220] = 0;
    exp_40_ram[1221] = 38;
    exp_40_ram[1222] = 9;
    exp_40_ram[1223] = 36;
    exp_40_ram[1224] = 37;
    exp_40_ram[1225] = 5;
    exp_40_ram[1226] = 137;
    exp_40_ram[1227] = 0;
    exp_40_ram[1228] = 135;
    exp_40_ram[1229] = 36;
    exp_40_ram[1230] = 38;
    exp_40_ram[1231] = 32;
    exp_40_ram[1232] = 34;
    exp_40_ram[1233] = 36;
    exp_40_ram[1234] = 40;
    exp_40_ram[1235] = 42;
    exp_40_ram[1236] = 133;
    exp_40_ram[1237] = 38;
    exp_40_ram[1238] = 5;
    exp_40_ram[1239] = 240;
    exp_40_ram[1240] = 44;
    exp_40_ram[1241] = 46;
    exp_40_ram[1242] = 32;
    exp_40_ram[1243] = 5;
    exp_40_ram[1244] = 36;
    exp_40_ram[1245] = 36;
    exp_40_ram[1246] = 41;
    exp_40_ram[1247] = 41;
    exp_40_ram[1248] = 42;
    exp_40_ram[1249] = 42;
    exp_40_ram[1250] = 43;
    exp_40_ram[1251] = 43;
    exp_40_ram[1252] = 44;
    exp_40_ram[1253] = 44;
    exp_40_ram[1254] = 1;
    exp_40_ram[1255] = 128;
    exp_40_ram[1256] = 1;
    exp_40_ram[1257] = 34;
    exp_40_ram[1258] = 42;
    exp_40_ram[1259] = 7;
    exp_40_ram[1260] = 42;
    exp_40_ram[1261] = 40;
    exp_40_ram[1262] = 36;
    exp_40_ram[1263] = 4;
    exp_40_ram[1264] = 10;
    exp_40_ram[1265] = 6;
    exp_40_ram[1266] = 9;
    exp_40_ram[1267] = 5;
    exp_40_ram[1268] = 5;
    exp_40_ram[1269] = 46;
    exp_40_ram[1270] = 36;
    exp_40_ram[1271] = 44;
    exp_40_ram[1272] = 38;
    exp_40_ram[1273] = 32;
    exp_40_ram[1274] = 34;
    exp_40_ram[1275] = 38;
    exp_40_ram[1276] = 46;
    exp_40_ram[1277] = 44;
    exp_40_ram[1278] = 44;
    exp_40_ram[1279] = 240;
    exp_40_ram[1280] = 5;
    exp_40_ram[1281] = 240;
    exp_40_ram[1282] = 134;
    exp_40_ram[1283] = 5;
    exp_40_ram[1284] = 5;
    exp_40_ram[1285] = 240;
    exp_40_ram[1286] = 39;
    exp_40_ram[1287] = 39;
    exp_40_ram[1288] = 6;
    exp_40_ram[1289] = 5;
    exp_40_ram[1290] = 135;
    exp_40_ram[1291] = 5;
    exp_40_ram[1292] = 34;
    exp_40_ram[1293] = 240;
    exp_40_ram[1294] = 5;
    exp_40_ram[1295] = 240;
    exp_40_ram[1296] = 7;
    exp_40_ram[1297] = 6;
    exp_40_ram[1298] = 9;
    exp_40_ram[1299] = 132;
    exp_40_ram[1300] = 5;
    exp_40_ram[1301] = 5;
    exp_40_ram[1302] = 38;
    exp_40_ram[1303] = 34;
    exp_40_ram[1304] = 36;
    exp_40_ram[1305] = 40;
    exp_40_ram[1306] = 32;
    exp_40_ram[1307] = 46;
    exp_40_ram[1308] = 240;
    exp_40_ram[1309] = 5;
    exp_40_ram[1310] = 240;
    exp_40_ram[1311] = 134;
    exp_40_ram[1312] = 5;
    exp_40_ram[1313] = 5;
    exp_40_ram[1314] = 240;
    exp_40_ram[1315] = 39;
    exp_40_ram[1316] = 39;
    exp_40_ram[1317] = 6;
    exp_40_ram[1318] = 5;
    exp_40_ram[1319] = 135;
    exp_40_ram[1320] = 5;
    exp_40_ram[1321] = 36;
    exp_40_ram[1322] = 240;
    exp_40_ram[1323] = 5;
    exp_40_ram[1324] = 240;
    exp_40_ram[1325] = 132;
    exp_40_ram[1326] = 10;
    exp_40_ram[1327] = 6;
    exp_40_ram[1328] = 5;
    exp_40_ram[1329] = 5;
    exp_40_ram[1330] = 240;
    exp_40_ram[1331] = 5;
    exp_40_ram[1332] = 240;
    exp_40_ram[1333] = 226;
    exp_40_ram[1334] = 7;
    exp_40_ram[1335] = 135;
    exp_40_ram[1336] = 148;
    exp_40_ram[1337] = 106;
    exp_40_ram[1338] = 5;
    exp_40_ram[1339] = 102;
    exp_40_ram[1340] = 150;
    exp_40_ram[1341] = 244;
    exp_40_ram[1342] = 5;
    exp_40_ram[1343] = 32;
    exp_40_ram[1344] = 36;
    exp_40_ram[1345] = 36;
    exp_40_ram[1346] = 41;
    exp_40_ram[1347] = 41;
    exp_40_ram[1348] = 42;
    exp_40_ram[1349] = 42;
    exp_40_ram[1350] = 1;
    exp_40_ram[1351] = 128;
    exp_40_ram[1352] = 1;
    exp_40_ram[1353] = 5;
    exp_40_ram[1354] = 40;
    exp_40_ram[1355] = 6;
    exp_40_ram[1356] = 9;
    exp_40_ram[1357] = 5;
    exp_40_ram[1358] = 46;
    exp_40_ram[1359] = 44;
    exp_40_ram[1360] = 42;
    exp_40_ram[1361] = 38;
    exp_40_ram[1362] = 240;
    exp_40_ram[1363] = 6;
    exp_40_ram[1364] = 5;
    exp_40_ram[1365] = 5;
    exp_40_ram[1366] = 41;
    exp_40_ram[1367] = 240;
    exp_40_ram[1368] = 5;
    exp_40_ram[1369] = 240;
    exp_40_ram[1370] = 4;
    exp_40_ram[1371] = 132;
    exp_40_ram[1372] = 88;
    exp_40_ram[1373] = 247;
    exp_40_ram[1374] = 135;
    exp_40_ram[1375] = 7;
    exp_40_ram[1376] = 183;
    exp_40_ram[1377] = 132;
    exp_40_ram[1378] = 132;
    exp_40_ram[1379] = 4;
    exp_40_ram[1380] = 133;
    exp_40_ram[1381] = 6;
    exp_40_ram[1382] = 5;
    exp_40_ram[1383] = 240;
    exp_40_ram[1384] = 6;
    exp_40_ram[1385] = 5;
    exp_40_ram[1386] = 5;
    exp_40_ram[1387] = 240;
    exp_40_ram[1388] = 88;
    exp_40_ram[1389] = 7;
    exp_40_ram[1390] = 32;
    exp_40_ram[1391] = 32;
    exp_40_ram[1392] = 5;
    exp_40_ram[1393] = 36;
    exp_40_ram[1394] = 41;
    exp_40_ram[1395] = 41;
    exp_40_ram[1396] = 133;
    exp_40_ram[1397] = 36;
    exp_40_ram[1398] = 1;
    exp_40_ram[1399] = 128;
    exp_40_ram[1400] = 136;
    exp_40_ram[1401] = 6;
    exp_40_ram[1402] = 5;
    exp_40_ram[1403] = 5;
    exp_40_ram[1404] = 240;
    exp_40_ram[1405] = 5;
    exp_40_ram[1406] = 240;
    exp_40_ram[1407] = 7;
    exp_40_ram[1408] = 6;
    exp_40_ram[1409] = 23;
    exp_40_ram[1410] = 135;
    exp_40_ram[1411] = 135;
    exp_40_ram[1412] = 183;
    exp_40_ram[1413] = 4;
    exp_40_ram[1414] = 132;
    exp_40_ram[1415] = 240;
    exp_40_ram[1416] = 130;
    exp_40_ram[1417] = 6;
    exp_40_ram[1418] = 5;
    exp_40_ram[1419] = 5;
    exp_40_ram[1420] = 240;
    exp_40_ram[1421] = 5;
    exp_40_ram[1422] = 240;
    exp_40_ram[1423] = 32;
    exp_40_ram[1424] = 240;
    exp_40_ram[1425] = 32;
    exp_40_ram[1426] = 240;
    exp_40_ram[1427] = 1;
    exp_40_ram[1428] = 134;
    exp_40_ram[1429] = 5;
    exp_40_ram[1430] = 5;
    exp_40_ram[1431] = 38;
    exp_40_ram[1432] = 240;
    exp_40_ram[1433] = 5;
    exp_40_ram[1434] = 6;
    exp_40_ram[1435] = 5;
    exp_40_ram[1436] = 240;
    exp_40_ram[1437] = 5;
    exp_40_ram[1438] = 240;
    exp_40_ram[1439] = 32;
    exp_40_ram[1440] = 1;
    exp_40_ram[1441] = 128;
    exp_40_ram[1442] = 37;
    exp_40_ram[1443] = 38;
    exp_40_ram[1444] = 1;
    exp_40_ram[1445] = 5;
    exp_40_ram[1446] = 46;
    exp_40_ram[1447] = 44;
    exp_40_ram[1448] = 240;
    exp_40_ram[1449] = 36;
    exp_40_ram[1450] = 5;
    exp_40_ram[1451] = 5;
    exp_40_ram[1452] = 6;
    exp_40_ram[1453] = 240;
    exp_40_ram[1454] = 32;
    exp_40_ram[1455] = 5;
    exp_40_ram[1456] = 36;
    exp_40_ram[1457] = 1;
    exp_40_ram[1458] = 128;
    exp_40_ram[1459] = 1;
    exp_40_ram[1460] = 34;
    exp_40_ram[1461] = 32;
    exp_40_ram[1462] = 36;
    exp_40_ram[1463] = 41;
    exp_40_ram[1464] = 38;
    exp_40_ram[1465] = 133;
    exp_40_ram[1466] = 5;
    exp_40_ram[1467] = 36;
    exp_40_ram[1468] = 46;
    exp_40_ram[1469] = 240;
    exp_40_ram[1470] = 6;
    exp_40_ram[1471] = 6;
    exp_40_ram[1472] = 22;
    exp_40_ram[1473] = 6;
    exp_40_ram[1474] = 5;
    exp_40_ram[1475] = 182;
    exp_40_ram[1476] = 6;
    exp_40_ram[1477] = 5;
    exp_40_ram[1478] = 240;
    exp_40_ram[1479] = 36;
    exp_40_ram[1480] = 5;
    exp_40_ram[1481] = 6;
    exp_40_ram[1482] = 5;
    exp_40_ram[1483] = 240;
    exp_40_ram[1484] = 5;
    exp_40_ram[1485] = 133;
    exp_40_ram[1486] = 240;
    exp_40_ram[1487] = 9;
    exp_40_ram[1488] = 160;
    exp_40_ram[1489] = 32;
    exp_40_ram[1490] = 5;
    exp_40_ram[1491] = 36;
    exp_40_ram[1492] = 36;
    exp_40_ram[1493] = 41;
    exp_40_ram[1494] = 41;
    exp_40_ram[1495] = 1;
    exp_40_ram[1496] = 128;
    exp_40_ram[1497] = 1;
    exp_40_ram[1498] = 38;
    exp_40_ram[1499] = 240;
    exp_40_ram[1500] = 32;
    exp_40_ram[1501] = 1;
    exp_40_ram[1502] = 240;
    exp_40_ram[1503] = 1;
    exp_40_ram[1504] = 38;
    exp_40_ram[1505] = 36;
    exp_40_ram[1506] = 4;
    exp_40_ram[1507] = 23;
    exp_40_ram[1508] = 133;
    exp_40_ram[1509] = 240;
    exp_40_ram[1510] = 23;
    exp_40_ram[1511] = 133;
    exp_40_ram[1512] = 240;
    exp_40_ram[1513] = 32;
    exp_40_ram[1514] = 36;
    exp_40_ram[1515] = 1;
    exp_40_ram[1516] = 128;
    exp_40_ram[1517] = 1;
    exp_40_ram[1518] = 46;
    exp_40_ram[1519] = 44;
    exp_40_ram[1520] = 42;
    exp_40_ram[1521] = 40;
    exp_40_ram[1522] = 38;
    exp_40_ram[1523] = 36;
    exp_40_ram[1524] = 34;
    exp_40_ram[1525] = 32;
    exp_40_ram[1526] = 4;
    exp_40_ram[1527] = 23;
    exp_40_ram[1528] = 133;
    exp_40_ram[1529] = 240;
    exp_40_ram[1530] = 7;
    exp_40_ram[1531] = 32;
    exp_40_ram[1532] = 7;
    exp_40_ram[1533] = 46;
    exp_40_ram[1534] = 7;
    exp_40_ram[1535] = 44;
    exp_40_ram[1536] = 7;
    exp_40_ram[1537] = 42;
    exp_40_ram[1538] = 7;
    exp_40_ram[1539] = 40;
    exp_40_ram[1540] = 38;
    exp_40_ram[1541] = 7;
    exp_40_ram[1542] = 38;
    exp_40_ram[1543] = 7;
    exp_40_ram[1544] = 133;
    exp_40_ram[1545] = 240;
    exp_40_ram[1546] = 7;
    exp_40_ram[1547] = 135;
    exp_40_ram[1548] = 32;
    exp_40_ram[1549] = 34;
    exp_40_ram[1550] = 7;
    exp_40_ram[1551] = 133;
    exp_40_ram[1552] = 240;
    exp_40_ram[1553] = 7;
    exp_40_ram[1554] = 23;
    exp_40_ram[1555] = 133;
    exp_40_ram[1556] = 5;
    exp_40_ram[1557] = 240;
    exp_40_ram[1558] = 7;
    exp_40_ram[1559] = 138;
    exp_40_ram[1560] = 23;
    exp_40_ram[1561] = 133;
    exp_40_ram[1562] = 240;
    exp_40_ram[1563] = 0;
    exp_40_ram[1564] = 7;
    exp_40_ram[1565] = 133;
    exp_40_ram[1566] = 240;
    exp_40_ram[1567] = 7;
    exp_40_ram[1568] = 133;
    exp_40_ram[1569] = 240;
    exp_40_ram[1570] = 7;
    exp_40_ram[1571] = 23;
    exp_40_ram[1572] = 133;
    exp_40_ram[1573] = 5;
    exp_40_ram[1574] = 240;
    exp_40_ram[1575] = 7;
    exp_40_ram[1576] = 138;
    exp_40_ram[1577] = 23;
    exp_40_ram[1578] = 133;
    exp_40_ram[1579] = 240;
    exp_40_ram[1580] = 0;
    exp_40_ram[1581] = 7;
    exp_40_ram[1582] = 133;
    exp_40_ram[1583] = 240;
    exp_40_ram[1584] = 7;
    exp_40_ram[1585] = 133;
    exp_40_ram[1586] = 240;
    exp_40_ram[1587] = 7;
    exp_40_ram[1588] = 23;
    exp_40_ram[1589] = 133;
    exp_40_ram[1590] = 5;
    exp_40_ram[1591] = 240;
    exp_40_ram[1592] = 7;
    exp_40_ram[1593] = 138;
    exp_40_ram[1594] = 23;
    exp_40_ram[1595] = 133;
    exp_40_ram[1596] = 240;
    exp_40_ram[1597] = 0;
    exp_40_ram[1598] = 7;
    exp_40_ram[1599] = 133;
    exp_40_ram[1600] = 240;
    exp_40_ram[1601] = 7;
    exp_40_ram[1602] = 23;
    exp_40_ram[1603] = 133;
    exp_40_ram[1604] = 5;
    exp_40_ram[1605] = 240;
    exp_40_ram[1606] = 7;
    exp_40_ram[1607] = 138;
    exp_40_ram[1608] = 23;
    exp_40_ram[1609] = 133;
    exp_40_ram[1610] = 240;
    exp_40_ram[1611] = 0;
    exp_40_ram[1612] = 7;
    exp_40_ram[1613] = 32;
    exp_40_ram[1614] = 7;
    exp_40_ram[1615] = 46;
    exp_40_ram[1616] = 7;
    exp_40_ram[1617] = 44;
    exp_40_ram[1618] = 7;
    exp_40_ram[1619] = 42;
    exp_40_ram[1620] = 7;
    exp_40_ram[1621] = 40;
    exp_40_ram[1622] = 38;
    exp_40_ram[1623] = 7;
    exp_40_ram[1624] = 38;
    exp_40_ram[1625] = 7;
    exp_40_ram[1626] = 133;
    exp_40_ram[1627] = 240;
    exp_40_ram[1628] = 7;
    exp_40_ram[1629] = 135;
    exp_40_ram[1630] = 32;
    exp_40_ram[1631] = 34;
    exp_40_ram[1632] = 7;
    exp_40_ram[1633] = 133;
    exp_40_ram[1634] = 240;
    exp_40_ram[1635] = 7;
    exp_40_ram[1636] = 23;
    exp_40_ram[1637] = 133;
    exp_40_ram[1638] = 5;
    exp_40_ram[1639] = 240;
    exp_40_ram[1640] = 7;
    exp_40_ram[1641] = 138;
    exp_40_ram[1642] = 23;
    exp_40_ram[1643] = 133;
    exp_40_ram[1644] = 240;
    exp_40_ram[1645] = 0;
    exp_40_ram[1646] = 7;
    exp_40_ram[1647] = 133;
    exp_40_ram[1648] = 240;
    exp_40_ram[1649] = 7;
    exp_40_ram[1650] = 133;
    exp_40_ram[1651] = 240;
    exp_40_ram[1652] = 7;
    exp_40_ram[1653] = 23;
    exp_40_ram[1654] = 133;
    exp_40_ram[1655] = 5;
    exp_40_ram[1656] = 240;
    exp_40_ram[1657] = 7;
    exp_40_ram[1658] = 138;
    exp_40_ram[1659] = 23;
    exp_40_ram[1660] = 133;
    exp_40_ram[1661] = 240;
    exp_40_ram[1662] = 0;
    exp_40_ram[1663] = 7;
    exp_40_ram[1664] = 133;
    exp_40_ram[1665] = 240;
    exp_40_ram[1666] = 7;
    exp_40_ram[1667] = 133;
    exp_40_ram[1668] = 240;
    exp_40_ram[1669] = 7;
    exp_40_ram[1670] = 23;
    exp_40_ram[1671] = 133;
    exp_40_ram[1672] = 5;
    exp_40_ram[1673] = 240;
    exp_40_ram[1674] = 7;
    exp_40_ram[1675] = 138;
    exp_40_ram[1676] = 23;
    exp_40_ram[1677] = 133;
    exp_40_ram[1678] = 240;
    exp_40_ram[1679] = 0;
    exp_40_ram[1680] = 7;
    exp_40_ram[1681] = 133;
    exp_40_ram[1682] = 240;
    exp_40_ram[1683] = 7;
    exp_40_ram[1684] = 23;
    exp_40_ram[1685] = 133;
    exp_40_ram[1686] = 5;
    exp_40_ram[1687] = 240;
    exp_40_ram[1688] = 7;
    exp_40_ram[1689] = 138;
    exp_40_ram[1690] = 23;
    exp_40_ram[1691] = 133;
    exp_40_ram[1692] = 240;
    exp_40_ram[1693] = 0;
    exp_40_ram[1694] = 7;
    exp_40_ram[1695] = 32;
    exp_40_ram[1696] = 7;
    exp_40_ram[1697] = 46;
    exp_40_ram[1698] = 7;
    exp_40_ram[1699] = 44;
    exp_40_ram[1700] = 7;
    exp_40_ram[1701] = 42;
    exp_40_ram[1702] = 7;
    exp_40_ram[1703] = 40;
    exp_40_ram[1704] = 38;
    exp_40_ram[1705] = 38;
    exp_40_ram[1706] = 7;
    exp_40_ram[1707] = 133;
    exp_40_ram[1708] = 240;
    exp_40_ram[1709] = 7;
    exp_40_ram[1710] = 135;
    exp_40_ram[1711] = 32;
    exp_40_ram[1712] = 34;
    exp_40_ram[1713] = 7;
    exp_40_ram[1714] = 133;
    exp_40_ram[1715] = 240;
    exp_40_ram[1716] = 7;
    exp_40_ram[1717] = 23;
    exp_40_ram[1718] = 133;
    exp_40_ram[1719] = 5;
    exp_40_ram[1720] = 240;
    exp_40_ram[1721] = 7;
    exp_40_ram[1722] = 138;
    exp_40_ram[1723] = 23;
    exp_40_ram[1724] = 133;
    exp_40_ram[1725] = 240;
    exp_40_ram[1726] = 0;
    exp_40_ram[1727] = 7;
    exp_40_ram[1728] = 133;
    exp_40_ram[1729] = 240;
    exp_40_ram[1730] = 7;
    exp_40_ram[1731] = 133;
    exp_40_ram[1732] = 240;
    exp_40_ram[1733] = 7;
    exp_40_ram[1734] = 23;
    exp_40_ram[1735] = 133;
    exp_40_ram[1736] = 5;
    exp_40_ram[1737] = 240;
    exp_40_ram[1738] = 7;
    exp_40_ram[1739] = 138;
    exp_40_ram[1740] = 23;
    exp_40_ram[1741] = 133;
    exp_40_ram[1742] = 240;
    exp_40_ram[1743] = 0;
    exp_40_ram[1744] = 7;
    exp_40_ram[1745] = 133;
    exp_40_ram[1746] = 240;
    exp_40_ram[1747] = 7;
    exp_40_ram[1748] = 133;
    exp_40_ram[1749] = 240;
    exp_40_ram[1750] = 7;
    exp_40_ram[1751] = 23;
    exp_40_ram[1752] = 133;
    exp_40_ram[1753] = 5;
    exp_40_ram[1754] = 240;
    exp_40_ram[1755] = 7;
    exp_40_ram[1756] = 138;
    exp_40_ram[1757] = 23;
    exp_40_ram[1758] = 133;
    exp_40_ram[1759] = 240;
    exp_40_ram[1760] = 0;
    exp_40_ram[1761] = 7;
    exp_40_ram[1762] = 133;
    exp_40_ram[1763] = 240;
    exp_40_ram[1764] = 7;
    exp_40_ram[1765] = 23;
    exp_40_ram[1766] = 133;
    exp_40_ram[1767] = 5;
    exp_40_ram[1768] = 240;
    exp_40_ram[1769] = 7;
    exp_40_ram[1770] = 138;
    exp_40_ram[1771] = 23;
    exp_40_ram[1772] = 133;
    exp_40_ram[1773] = 224;
    exp_40_ram[1774] = 0;
    exp_40_ram[1775] = 23;
    exp_40_ram[1776] = 133;
    exp_40_ram[1777] = 224;
    exp_40_ram[1778] = 7;
    exp_40_ram[1779] = 32;
    exp_40_ram[1780] = 7;
    exp_40_ram[1781] = 46;
    exp_40_ram[1782] = 7;
    exp_40_ram[1783] = 44;
    exp_40_ram[1784] = 42;
    exp_40_ram[1785] = 7;
    exp_40_ram[1786] = 40;
    exp_40_ram[1787] = 7;
    exp_40_ram[1788] = 38;
    exp_40_ram[1789] = 7;
    exp_40_ram[1790] = 38;
    exp_40_ram[1791] = 7;
    exp_40_ram[1792] = 133;
    exp_40_ram[1793] = 240;
    exp_40_ram[1794] = 7;
    exp_40_ram[1795] = 135;
    exp_40_ram[1796] = 32;
    exp_40_ram[1797] = 34;
    exp_40_ram[1798] = 39;
    exp_40_ram[1799] = 39;
    exp_40_ram[1800] = 5;
    exp_40_ram[1801] = 133;
    exp_40_ram[1802] = 240;
    exp_40_ram[1803] = 240;
    exp_40_ram[1804] = 44;
    exp_40_ram[1805] = 46;
    exp_40_ram[1806] = 42;
    exp_40_ram[1807] = 0;
    exp_40_ram[1808] = 0;
    exp_40_ram[1809] = 240;
    exp_40_ram[1810] = 7;
    exp_40_ram[1811] = 135;
    exp_40_ram[1812] = 38;
    exp_40_ram[1813] = 38;
    exp_40_ram[1814] = 5;
    exp_40_ram[1815] = 133;
    exp_40_ram[1816] = 240;
    exp_40_ram[1817] = 11;
    exp_40_ram[1818] = 139;
    exp_40_ram[1819] = 39;
    exp_40_ram[1820] = 167;
    exp_40_ram[1821] = 133;
    exp_40_ram[1822] = 224;
    exp_40_ram[1823] = 7;
    exp_40_ram[1824] = 135;
    exp_40_ram[1825] = 6;
    exp_40_ram[1826] = 134;
    exp_40_ram[1827] = 5;
    exp_40_ram[1828] = 133;
    exp_40_ram[1829] = 224;
    exp_40_ram[1830] = 7;
    exp_40_ram[1831] = 196;
    exp_40_ram[1832] = 39;
    exp_40_ram[1833] = 167;
    exp_40_ram[1834] = 138;
    exp_40_ram[1835] = 10;
    exp_40_ram[1836] = 38;
    exp_40_ram[1837] = 38;
    exp_40_ram[1838] = 7;
    exp_40_ram[1839] = 5;
    exp_40_ram[1840] = 181;
    exp_40_ram[1841] = 135;
    exp_40_ram[1842] = 134;
    exp_40_ram[1843] = 135;
    exp_40_ram[1844] = 44;
    exp_40_ram[1845] = 46;
    exp_40_ram[1846] = 5;
    exp_40_ram[1847] = 240;
    exp_40_ram[1848] = 7;
    exp_40_ram[1849] = 135;
    exp_40_ram[1850] = 32;
    exp_40_ram[1851] = 34;
    exp_40_ram[1852] = 7;
    exp_40_ram[1853] = 133;
    exp_40_ram[1854] = 240;
    exp_40_ram[1855] = 7;
    exp_40_ram[1856] = 133;
    exp_40_ram[1857] = 224;
    exp_40_ram[1858] = 39;
    exp_40_ram[1859] = 135;
    exp_40_ram[1860] = 42;
    exp_40_ram[1861] = 39;
    exp_40_ram[1862] = 7;
    exp_40_ram[1863] = 210;
    exp_40_ram[1864] = 7;
    exp_40_ram[1865] = 32;
    exp_40_ram[1866] = 7;
    exp_40_ram[1867] = 46;
    exp_40_ram[1868] = 7;
    exp_40_ram[1869] = 44;
    exp_40_ram[1870] = 7;
    exp_40_ram[1871] = 42;
    exp_40_ram[1872] = 7;
    exp_40_ram[1873] = 40;
    exp_40_ram[1874] = 7;
    exp_40_ram[1875] = 38;
    exp_40_ram[1876] = 7;
    exp_40_ram[1877] = 38;
    exp_40_ram[1878] = 7;
    exp_40_ram[1879] = 133;
    exp_40_ram[1880] = 240;
    exp_40_ram[1881] = 7;
    exp_40_ram[1882] = 135;
    exp_40_ram[1883] = 32;
    exp_40_ram[1884] = 34;
    exp_40_ram[1885] = 7;
    exp_40_ram[1886] = 133;
    exp_40_ram[1887] = 240;
    exp_40_ram[1888] = 7;
    exp_40_ram[1889] = 133;
    exp_40_ram[1890] = 224;
    exp_40_ram[1891] = 7;
    exp_40_ram[1892] = 133;
    exp_40_ram[1893] = 240;
    exp_40_ram[1894] = 7;
    exp_40_ram[1895] = 133;
    exp_40_ram[1896] = 224;
    exp_40_ram[1897] = 39;
    exp_40_ram[1898] = 39;
    exp_40_ram[1899] = 5;
    exp_40_ram[1900] = 133;
    exp_40_ram[1901] = 240;
    exp_40_ram[1902] = 5;
    exp_40_ram[1903] = 240;
    exp_40_ram[1904] = 7;
    exp_40_ram[1905] = 135;
    exp_40_ram[1906] = 32;
    exp_40_ram[1907] = 34;
    exp_40_ram[1908] = 7;
    exp_40_ram[1909] = 133;
    exp_40_ram[1910] = 240;
    exp_40_ram[1911] = 7;
    exp_40_ram[1912] = 133;
    exp_40_ram[1913] = 224;
    exp_40_ram[1914] = 224;
    exp_40_ram[1915] = 44;
    exp_40_ram[1916] = 46;
    exp_40_ram[1917] = 40;
    exp_40_ram[1918] = 0;
    exp_40_ram[1919] = 0;
    exp_40_ram[1920] = 224;
    exp_40_ram[1921] = 7;
    exp_40_ram[1922] = 135;
    exp_40_ram[1923] = 38;
    exp_40_ram[1924] = 38;
    exp_40_ram[1925] = 5;
    exp_40_ram[1926] = 133;
    exp_40_ram[1927] = 224;
    exp_40_ram[1928] = 10;
    exp_40_ram[1929] = 138;
    exp_40_ram[1930] = 39;
    exp_40_ram[1931] = 167;
    exp_40_ram[1932] = 133;
    exp_40_ram[1933] = 224;
    exp_40_ram[1934] = 7;
    exp_40_ram[1935] = 135;
    exp_40_ram[1936] = 6;
    exp_40_ram[1937] = 134;
    exp_40_ram[1938] = 5;
    exp_40_ram[1939] = 133;
    exp_40_ram[1940] = 224;
    exp_40_ram[1941] = 7;
    exp_40_ram[1942] = 196;
    exp_40_ram[1943] = 39;
    exp_40_ram[1944] = 167;
    exp_40_ram[1945] = 137;
    exp_40_ram[1946] = 9;
    exp_40_ram[1947] = 38;
    exp_40_ram[1948] = 38;
    exp_40_ram[1949] = 7;
    exp_40_ram[1950] = 5;
    exp_40_ram[1951] = 181;
    exp_40_ram[1952] = 135;
    exp_40_ram[1953] = 134;
    exp_40_ram[1954] = 135;
    exp_40_ram[1955] = 44;
    exp_40_ram[1956] = 46;
    exp_40_ram[1957] = 5;
    exp_40_ram[1958] = 240;
    exp_40_ram[1959] = 7;
    exp_40_ram[1960] = 135;
    exp_40_ram[1961] = 32;
    exp_40_ram[1962] = 34;
    exp_40_ram[1963] = 7;
    exp_40_ram[1964] = 133;
    exp_40_ram[1965] = 240;
    exp_40_ram[1966] = 7;
    exp_40_ram[1967] = 133;
    exp_40_ram[1968] = 224;
    exp_40_ram[1969] = 39;
    exp_40_ram[1970] = 135;
    exp_40_ram[1971] = 40;
    exp_40_ram[1972] = 39;
    exp_40_ram[1973] = 7;
    exp_40_ram[1974] = 210;
    exp_40_ram[1975] = 32;
    exp_40_ram[1976] = 36;
    exp_40_ram[1977] = 41;
    exp_40_ram[1978] = 41;
    exp_40_ram[1979] = 42;
    exp_40_ram[1980] = 42;
    exp_40_ram[1981] = 43;
    exp_40_ram[1982] = 43;
    exp_40_ram[1983] = 1;
    exp_40_ram[1984] = 128;
    exp_40_ram[1985] = 1;
    exp_40_ram[1986] = 38;
    exp_40_ram[1987] = 36;
    exp_40_ram[1988] = 4;
    exp_40_ram[1989] = 240;
    exp_40_ram[1990] = 240;
    exp_40_ram[1991] = 0;
    exp_40_ram[1992] = 32;
    exp_40_ram[1993] = 36;
    exp_40_ram[1994] = 1;
    exp_40_ram[1995] = 128;
    exp_40_ram[1996] = 7;
    exp_40_ram[1997] = 135;
    exp_40_ram[1998] = 69;
    exp_40_ram[1999] = 1;
    exp_40_ram[2000] = 101;
    exp_40_ram[2001] = 76;
    exp_40_ram[2002] = 214;
    exp_40_ram[2003] = 5;
    exp_40_ram[2004] = 133;
    exp_40_ram[2005] = 1;
    exp_40_ram[2006] = 128;
    exp_40_ram[2007] = 92;
    exp_40_ram[2008] = 5;
    exp_40_ram[2009] = 133;
    exp_40_ram[2010] = 240;
    exp_40_ram[2011] = 240;
    exp_40_ram[2012] = 0;
    exp_40_ram[2013] = 117;
    exp_40_ram[2014] = 110;
    exp_40_ram[2015] = 87;
    exp_40_ram[2016] = 104;
    exp_40_ram[2017] = 105;
    exp_40_ram[2018] = 0;
    exp_40_ram[2019] = 97;
    exp_40_ram[2020] = 98;
    exp_40_ram[2021] = 65;
    exp_40_ram[2022] = 97;
    exp_40_ram[2023] = 110;
    exp_40_ram[2024] = 65;
    exp_40_ram[2025] = 101;
    exp_40_ram[2026] = 116;
    exp_40_ram[2027] = 68;
    exp_40_ram[2028] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_38) begin
      exp_40_ram[exp_34] <= exp_36;
    end
  end
  assign exp_40 = exp_40_ram[exp_35];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_66) begin
        exp_40_ram[exp_62] <= exp_64;
    end
  end
  assign exp_68 = exp_40_ram[exp_63];
  assign exp_67 = exp_90;
  assign exp_90 = 1;
  assign exp_63 = exp_89;
  assign exp_89 = exp_8[31:2];
  assign exp_66 = exp_84;
  assign exp_62 = exp_83;
  assign exp_64 = exp_83;
  assign exp_39 = exp_125;
  assign exp_125 = 1;
  assign exp_35 = exp_124;
  assign exp_124 = exp_10[31:2];
  assign exp_38 = exp_106;
  assign exp_106 = exp_104 & exp_105;
  assign exp_104 = exp_14 & exp_15;
  assign exp_105 = exp_16[1:1];
  assign exp_34 = exp_102;
  assign exp_102 = exp_10[31:2];
  assign exp_36 = exp_103;
  assign exp_103 = exp_11[15:8];

  //Create RAM
  reg [7:0] exp_33_ram [4095:0];


  //Initialise RAM contents
  initial
  begin
    exp_33_ram[0] = 147;
    exp_33_ram[1] = 19;
    exp_33_ram[2] = 147;
    exp_33_ram[3] = 19;
    exp_33_ram[4] = 147;
    exp_33_ram[5] = 19;
    exp_33_ram[6] = 147;
    exp_33_ram[7] = 19;
    exp_33_ram[8] = 147;
    exp_33_ram[9] = 19;
    exp_33_ram[10] = 147;
    exp_33_ram[11] = 19;
    exp_33_ram[12] = 147;
    exp_33_ram[13] = 19;
    exp_33_ram[14] = 147;
    exp_33_ram[15] = 19;
    exp_33_ram[16] = 147;
    exp_33_ram[17] = 19;
    exp_33_ram[18] = 147;
    exp_33_ram[19] = 19;
    exp_33_ram[20] = 147;
    exp_33_ram[21] = 19;
    exp_33_ram[22] = 147;
    exp_33_ram[23] = 19;
    exp_33_ram[24] = 147;
    exp_33_ram[25] = 19;
    exp_33_ram[26] = 147;
    exp_33_ram[27] = 19;
    exp_33_ram[28] = 147;
    exp_33_ram[29] = 19;
    exp_33_ram[30] = 147;
    exp_33_ram[31] = 55;
    exp_33_ram[32] = 19;
    exp_33_ram[33] = 239;
    exp_33_ram[34] = 111;
    exp_33_ram[35] = 147;
    exp_33_ram[36] = 147;
    exp_33_ram[37] = 19;
    exp_33_ram[38] = 19;
    exp_33_ram[39] = 19;
    exp_33_ram[40] = 99;
    exp_33_ram[41] = 183;
    exp_33_ram[42] = 147;
    exp_33_ram[43] = 99;
    exp_33_ram[44] = 55;
    exp_33_ram[45] = 99;
    exp_33_ram[46] = 19;
    exp_33_ram[47] = 51;
    exp_33_ram[48] = 19;
    exp_33_ram[49] = 51;
    exp_33_ram[50] = 179;
    exp_33_ram[51] = 131;
    exp_33_ram[52] = 19;
    exp_33_ram[53] = 51;
    exp_33_ram[54] = 179;
    exp_33_ram[55] = 99;
    exp_33_ram[56] = 179;
    exp_33_ram[57] = 51;
    exp_33_ram[58] = 51;
    exp_33_ram[59] = 179;
    exp_33_ram[60] = 51;
    exp_33_ram[61] = 147;
    exp_33_ram[62] = 179;
    exp_33_ram[63] = 19;
    exp_33_ram[64] = 19;
    exp_33_ram[65] = 147;
    exp_33_ram[66] = 51;
    exp_33_ram[67] = 19;
    exp_33_ram[68] = 179;
    exp_33_ram[69] = 19;
    exp_33_ram[70] = 179;
    exp_33_ram[71] = 99;
    exp_33_ram[72] = 179;
    exp_33_ram[73] = 19;
    exp_33_ram[74] = 99;
    exp_33_ram[75] = 99;
    exp_33_ram[76] = 19;
    exp_33_ram[77] = 179;
    exp_33_ram[78] = 179;
    exp_33_ram[79] = 51;
    exp_33_ram[80] = 19;
    exp_33_ram[81] = 19;
    exp_33_ram[82] = 179;
    exp_33_ram[83] = 19;
    exp_33_ram[84] = 51;
    exp_33_ram[85] = 179;
    exp_33_ram[86] = 19;
    exp_33_ram[87] = 99;
    exp_33_ram[88] = 51;
    exp_33_ram[89] = 19;
    exp_33_ram[90] = 99;
    exp_33_ram[91] = 99;
    exp_33_ram[92] = 19;
    exp_33_ram[93] = 19;
    exp_33_ram[94] = 51;
    exp_33_ram[95] = 147;
    exp_33_ram[96] = 111;
    exp_33_ram[97] = 55;
    exp_33_ram[98] = 19;
    exp_33_ram[99] = 227;
    exp_33_ram[100] = 19;
    exp_33_ram[101] = 111;
    exp_33_ram[102] = 99;
    exp_33_ram[103] = 19;
    exp_33_ram[104] = 51;
    exp_33_ram[105] = 55;
    exp_33_ram[106] = 99;
    exp_33_ram[107] = 19;
    exp_33_ram[108] = 99;
    exp_33_ram[109] = 19;
    exp_33_ram[110] = 51;
    exp_33_ram[111] = 179;
    exp_33_ram[112] = 3;
    exp_33_ram[113] = 19;
    exp_33_ram[114] = 51;
    exp_33_ram[115] = 179;
    exp_33_ram[116] = 99;
    exp_33_ram[117] = 179;
    exp_33_ram[118] = 147;
    exp_33_ram[119] = 147;
    exp_33_ram[120] = 19;
    exp_33_ram[121] = 19;
    exp_33_ram[122] = 19;
    exp_33_ram[123] = 179;
    exp_33_ram[124] = 179;
    exp_33_ram[125] = 147;
    exp_33_ram[126] = 51;
    exp_33_ram[127] = 51;
    exp_33_ram[128] = 19;
    exp_33_ram[129] = 99;
    exp_33_ram[130] = 51;
    exp_33_ram[131] = 19;
    exp_33_ram[132] = 99;
    exp_33_ram[133] = 99;
    exp_33_ram[134] = 19;
    exp_33_ram[135] = 51;
    exp_33_ram[136] = 51;
    exp_33_ram[137] = 179;
    exp_33_ram[138] = 19;
    exp_33_ram[139] = 19;
    exp_33_ram[140] = 51;
    exp_33_ram[141] = 147;
    exp_33_ram[142] = 51;
    exp_33_ram[143] = 179;
    exp_33_ram[144] = 19;
    exp_33_ram[145] = 99;
    exp_33_ram[146] = 51;
    exp_33_ram[147] = 19;
    exp_33_ram[148] = 99;
    exp_33_ram[149] = 99;
    exp_33_ram[150] = 19;
    exp_33_ram[151] = 19;
    exp_33_ram[152] = 51;
    exp_33_ram[153] = 103;
    exp_33_ram[154] = 55;
    exp_33_ram[155] = 19;
    exp_33_ram[156] = 227;
    exp_33_ram[157] = 19;
    exp_33_ram[158] = 111;
    exp_33_ram[159] = 51;
    exp_33_ram[160] = 51;
    exp_33_ram[161] = 51;
    exp_33_ram[162] = 179;
    exp_33_ram[163] = 51;
    exp_33_ram[164] = 147;
    exp_33_ram[165] = 51;
    exp_33_ram[166] = 51;
    exp_33_ram[167] = 147;
    exp_33_ram[168] = 147;
    exp_33_ram[169] = 147;
    exp_33_ram[170] = 51;
    exp_33_ram[171] = 19;
    exp_33_ram[172] = 51;
    exp_33_ram[173] = 179;
    exp_33_ram[174] = 147;
    exp_33_ram[175] = 99;
    exp_33_ram[176] = 51;
    exp_33_ram[177] = 147;
    exp_33_ram[178] = 99;
    exp_33_ram[179] = 99;
    exp_33_ram[180] = 147;
    exp_33_ram[181] = 51;
    exp_33_ram[182] = 179;
    exp_33_ram[183] = 51;
    exp_33_ram[184] = 19;
    exp_33_ram[185] = 19;
    exp_33_ram[186] = 179;
    exp_33_ram[187] = 19;
    exp_33_ram[188] = 51;
    exp_33_ram[189] = 179;
    exp_33_ram[190] = 19;
    exp_33_ram[191] = 99;
    exp_33_ram[192] = 179;
    exp_33_ram[193] = 19;
    exp_33_ram[194] = 99;
    exp_33_ram[195] = 99;
    exp_33_ram[196] = 19;
    exp_33_ram[197] = 179;
    exp_33_ram[198] = 147;
    exp_33_ram[199] = 179;
    exp_33_ram[200] = 179;
    exp_33_ram[201] = 111;
    exp_33_ram[202] = 99;
    exp_33_ram[203] = 55;
    exp_33_ram[204] = 99;
    exp_33_ram[205] = 19;
    exp_33_ram[206] = 179;
    exp_33_ram[207] = 147;
    exp_33_ram[208] = 55;
    exp_33_ram[209] = 51;
    exp_33_ram[210] = 19;
    exp_33_ram[211] = 51;
    exp_33_ram[212] = 3;
    exp_33_ram[213] = 19;
    exp_33_ram[214] = 51;
    exp_33_ram[215] = 179;
    exp_33_ram[216] = 99;
    exp_33_ram[217] = 19;
    exp_33_ram[218] = 227;
    exp_33_ram[219] = 51;
    exp_33_ram[220] = 19;
    exp_33_ram[221] = 111;
    exp_33_ram[222] = 55;
    exp_33_ram[223] = 147;
    exp_33_ram[224] = 227;
    exp_33_ram[225] = 147;
    exp_33_ram[226] = 111;
    exp_33_ram[227] = 51;
    exp_33_ram[228] = 179;
    exp_33_ram[229] = 51;
    exp_33_ram[230] = 51;
    exp_33_ram[231] = 147;
    exp_33_ram[232] = 179;
    exp_33_ram[233] = 179;
    exp_33_ram[234] = 51;
    exp_33_ram[235] = 51;
    exp_33_ram[236] = 51;
    exp_33_ram[237] = 147;
    exp_33_ram[238] = 147;
    exp_33_ram[239] = 19;
    exp_33_ram[240] = 51;
    exp_33_ram[241] = 147;
    exp_33_ram[242] = 51;
    exp_33_ram[243] = 51;
    exp_33_ram[244] = 19;
    exp_33_ram[245] = 99;
    exp_33_ram[246] = 51;
    exp_33_ram[247] = 19;
    exp_33_ram[248] = 99;
    exp_33_ram[249] = 99;
    exp_33_ram[250] = 19;
    exp_33_ram[251] = 51;
    exp_33_ram[252] = 51;
    exp_33_ram[253] = 179;
    exp_33_ram[254] = 51;
    exp_33_ram[255] = 147;
    exp_33_ram[256] = 51;
    exp_33_ram[257] = 147;
    exp_33_ram[258] = 147;
    exp_33_ram[259] = 179;
    exp_33_ram[260] = 19;
    exp_33_ram[261] = 99;
    exp_33_ram[262] = 179;
    exp_33_ram[263] = 19;
    exp_33_ram[264] = 99;
    exp_33_ram[265] = 99;
    exp_33_ram[266] = 19;
    exp_33_ram[267] = 179;
    exp_33_ram[268] = 19;
    exp_33_ram[269] = 183;
    exp_33_ram[270] = 51;
    exp_33_ram[271] = 147;
    exp_33_ram[272] = 51;
    exp_33_ram[273] = 19;
    exp_33_ram[274] = 179;
    exp_33_ram[275] = 19;
    exp_33_ram[276] = 179;
    exp_33_ram[277] = 51;
    exp_33_ram[278] = 179;
    exp_33_ram[279] = 19;
    exp_33_ram[280] = 51;
    exp_33_ram[281] = 51;
    exp_33_ram[282] = 51;
    exp_33_ram[283] = 51;
    exp_33_ram[284] = 99;
    exp_33_ram[285] = 51;
    exp_33_ram[286] = 147;
    exp_33_ram[287] = 51;
    exp_33_ram[288] = 99;
    exp_33_ram[289] = 227;
    exp_33_ram[290] = 183;
    exp_33_ram[291] = 147;
    exp_33_ram[292] = 51;
    exp_33_ram[293] = 19;
    exp_33_ram[294] = 51;
    exp_33_ram[295] = 179;
    exp_33_ram[296] = 51;
    exp_33_ram[297] = 147;
    exp_33_ram[298] = 227;
    exp_33_ram[299] = 19;
    exp_33_ram[300] = 111;
    exp_33_ram[301] = 147;
    exp_33_ram[302] = 19;
    exp_33_ram[303] = 111;
    exp_33_ram[304] = 55;
    exp_33_ram[305] = 19;
    exp_33_ram[306] = 19;
    exp_33_ram[307] = 179;
    exp_33_ram[308] = 147;
    exp_33_ram[309] = 19;
    exp_33_ram[310] = 19;
    exp_33_ram[311] = 19;
    exp_33_ram[312] = 147;
    exp_33_ram[313] = 147;
    exp_33_ram[314] = 51;
    exp_33_ram[315] = 19;
    exp_33_ram[316] = 147;
    exp_33_ram[317] = 147;
    exp_33_ram[318] = 99;
    exp_33_ram[319] = 179;
    exp_33_ram[320] = 99;
    exp_33_ram[321] = 19;
    exp_33_ram[322] = 103;
    exp_33_ram[323] = 99;
    exp_33_ram[324] = 179;
    exp_33_ram[325] = 227;
    exp_33_ram[326] = 99;
    exp_33_ram[327] = 179;
    exp_33_ram[328] = 147;
    exp_33_ram[329] = 99;
    exp_33_ram[330] = 51;
    exp_33_ram[331] = 99;
    exp_33_ram[332] = 99;
    exp_33_ram[333] = 99;
    exp_33_ram[334] = 99;
    exp_33_ram[335] = 99;
    exp_33_ram[336] = 19;
    exp_33_ram[337] = 103;
    exp_33_ram[338] = 19;
    exp_33_ram[339] = 99;
    exp_33_ram[340] = 19;
    exp_33_ram[341] = 103;
    exp_33_ram[342] = 99;
    exp_33_ram[343] = 227;
    exp_33_ram[344] = 103;
    exp_33_ram[345] = 227;
    exp_33_ram[346] = 99;
    exp_33_ram[347] = 227;
    exp_33_ram[348] = 227;
    exp_33_ram[349] = 19;
    exp_33_ram[350] = 103;
    exp_33_ram[351] = 19;
    exp_33_ram[352] = 103;
    exp_33_ram[353] = 227;
    exp_33_ram[354] = 111;
    exp_33_ram[355] = 227;
    exp_33_ram[356] = 111;
    exp_33_ram[357] = 227;
    exp_33_ram[358] = 227;
    exp_33_ram[359] = 147;
    exp_33_ram[360] = 111;
    exp_33_ram[361] = 19;
    exp_33_ram[362] = 35;
    exp_33_ram[363] = 35;
    exp_33_ram[364] = 19;
    exp_33_ram[365] = 99;
    exp_33_ram[366] = 239;
    exp_33_ram[367] = 19;
    exp_33_ram[368] = 147;
    exp_33_ram[369] = 51;
    exp_33_ram[370] = 99;
    exp_33_ram[371] = 147;
    exp_33_ram[372] = 179;
    exp_33_ram[373] = 19;
    exp_33_ram[374] = 179;
    exp_33_ram[375] = 51;
    exp_33_ram[376] = 131;
    exp_33_ram[377] = 19;
    exp_33_ram[378] = 147;
    exp_33_ram[379] = 3;
    exp_33_ram[380] = 19;
    exp_33_ram[381] = 147;
    exp_33_ram[382] = 179;
    exp_33_ram[383] = 147;
    exp_33_ram[384] = 19;
    exp_33_ram[385] = 103;
    exp_33_ram[386] = 147;
    exp_33_ram[387] = 179;
    exp_33_ram[388] = 19;
    exp_33_ram[389] = 111;
    exp_33_ram[390] = 147;
    exp_33_ram[391] = 19;
    exp_33_ram[392] = 111;
    exp_33_ram[393] = 19;
    exp_33_ram[394] = 35;
    exp_33_ram[395] = 35;
    exp_33_ram[396] = 35;
    exp_33_ram[397] = 35;
    exp_33_ram[398] = 35;
    exp_33_ram[399] = 35;
    exp_33_ram[400] = 179;
    exp_33_ram[401] = 99;
    exp_33_ram[402] = 19;
    exp_33_ram[403] = 19;
    exp_33_ram[404] = 147;
    exp_33_ram[405] = 99;
    exp_33_ram[406] = 19;
    exp_33_ram[407] = 239;
    exp_33_ram[408] = 147;
    exp_33_ram[409] = 19;
    exp_33_ram[410] = 51;
    exp_33_ram[411] = 147;
    exp_33_ram[412] = 99;
    exp_33_ram[413] = 19;
    exp_33_ram[414] = 147;
    exp_33_ram[415] = 99;
    exp_33_ram[416] = 19;
    exp_33_ram[417] = 99;
    exp_33_ram[418] = 147;
    exp_33_ram[419] = 19;
    exp_33_ram[420] = 179;
    exp_33_ram[421] = 179;
    exp_33_ram[422] = 179;
    exp_33_ram[423] = 179;
    exp_33_ram[424] = 179;
    exp_33_ram[425] = 131;
    exp_33_ram[426] = 3;
    exp_33_ram[427] = 147;
    exp_33_ram[428] = 19;
    exp_33_ram[429] = 147;
    exp_33_ram[430] = 51;
    exp_33_ram[431] = 131;
    exp_33_ram[432] = 3;
    exp_33_ram[433] = 131;
    exp_33_ram[434] = 3;
    exp_33_ram[435] = 19;
    exp_33_ram[436] = 147;
    exp_33_ram[437] = 19;
    exp_33_ram[438] = 103;
    exp_33_ram[439] = 239;
    exp_33_ram[440] = 147;
    exp_33_ram[441] = 111;
    exp_33_ram[442] = 147;
    exp_33_ram[443] = 179;
    exp_33_ram[444] = 147;
    exp_33_ram[445] = 111;
    exp_33_ram[446] = 147;
    exp_33_ram[447] = 99;
    exp_33_ram[448] = 19;
    exp_33_ram[449] = 19;
    exp_33_ram[450] = 147;
    exp_33_ram[451] = 239;
    exp_33_ram[452] = 51;
    exp_33_ram[453] = 19;
    exp_33_ram[454] = 179;
    exp_33_ram[455] = 147;
    exp_33_ram[456] = 19;
    exp_33_ram[457] = 51;
    exp_33_ram[458] = 239;
    exp_33_ram[459] = 51;
    exp_33_ram[460] = 19;
    exp_33_ram[461] = 19;
    exp_33_ram[462] = 147;
    exp_33_ram[463] = 147;
    exp_33_ram[464] = 99;
    exp_33_ram[465] = 19;
    exp_33_ram[466] = 99;
    exp_33_ram[467] = 19;
    exp_33_ram[468] = 179;
    exp_33_ram[469] = 19;
    exp_33_ram[470] = 51;
    exp_33_ram[471] = 51;
    exp_33_ram[472] = 179;
    exp_33_ram[473] = 179;
    exp_33_ram[474] = 55;
    exp_33_ram[475] = 19;
    exp_33_ram[476] = 179;
    exp_33_ram[477] = 19;
    exp_33_ram[478] = 99;
    exp_33_ram[479] = 19;
    exp_33_ram[480] = 147;
    exp_33_ram[481] = 99;
    exp_33_ram[482] = 19;
    exp_33_ram[483] = 179;
    exp_33_ram[484] = 179;
    exp_33_ram[485] = 147;
    exp_33_ram[486] = 55;
    exp_33_ram[487] = 51;
    exp_33_ram[488] = 99;
    exp_33_ram[489] = 55;
    exp_33_ram[490] = 19;
    exp_33_ram[491] = 19;
    exp_33_ram[492] = 179;
    exp_33_ram[493] = 51;
    exp_33_ram[494] = 147;
    exp_33_ram[495] = 19;
    exp_33_ram[496] = 179;
    exp_33_ram[497] = 147;
    exp_33_ram[498] = 111;
    exp_33_ram[499] = 147;
    exp_33_ram[500] = 179;
    exp_33_ram[501] = 147;
    exp_33_ram[502] = 111;
    exp_33_ram[503] = 147;
    exp_33_ram[504] = 147;
    exp_33_ram[505] = 19;
    exp_33_ram[506] = 111;
    exp_33_ram[507] = 19;
    exp_33_ram[508] = 19;
    exp_33_ram[509] = 147;
    exp_33_ram[510] = 99;
    exp_33_ram[511] = 51;
    exp_33_ram[512] = 147;
    exp_33_ram[513] = 19;
    exp_33_ram[514] = 227;
    exp_33_ram[515] = 103;
    exp_33_ram[516] = 99;
    exp_33_ram[517] = 99;
    exp_33_ram[518] = 19;
    exp_33_ram[519] = 147;
    exp_33_ram[520] = 19;
    exp_33_ram[521] = 99;
    exp_33_ram[522] = 147;
    exp_33_ram[523] = 99;
    exp_33_ram[524] = 99;
    exp_33_ram[525] = 19;
    exp_33_ram[526] = 147;
    exp_33_ram[527] = 227;
    exp_33_ram[528] = 19;
    exp_33_ram[529] = 99;
    exp_33_ram[530] = 179;
    exp_33_ram[531] = 51;
    exp_33_ram[532] = 147;
    exp_33_ram[533] = 19;
    exp_33_ram[534] = 227;
    exp_33_ram[535] = 103;
    exp_33_ram[536] = 147;
    exp_33_ram[537] = 239;
    exp_33_ram[538] = 19;
    exp_33_ram[539] = 103;
    exp_33_ram[540] = 51;
    exp_33_ram[541] = 99;
    exp_33_ram[542] = 179;
    exp_33_ram[543] = 111;
    exp_33_ram[544] = 179;
    exp_33_ram[545] = 147;
    exp_33_ram[546] = 239;
    exp_33_ram[547] = 51;
    exp_33_ram[548] = 103;
    exp_33_ram[549] = 147;
    exp_33_ram[550] = 99;
    exp_33_ram[551] = 99;
    exp_33_ram[552] = 239;
    exp_33_ram[553] = 19;
    exp_33_ram[554] = 103;
    exp_33_ram[555] = 179;
    exp_33_ram[556] = 227;
    exp_33_ram[557] = 51;
    exp_33_ram[558] = 239;
    exp_33_ram[559] = 51;
    exp_33_ram[560] = 103;
    exp_33_ram[561] = 99;
    exp_33_ram[562] = 147;
    exp_33_ram[563] = 179;
    exp_33_ram[564] = 99;
    exp_33_ram[565] = 19;
    exp_33_ram[566] = 19;
    exp_33_ram[567] = 51;
    exp_33_ram[568] = 147;
    exp_33_ram[569] = 103;
    exp_33_ram[570] = 51;
    exp_33_ram[571] = 51;
    exp_33_ram[572] = 179;
    exp_33_ram[573] = 51;
    exp_33_ram[574] = 111;
    exp_33_ram[575] = 99;
    exp_33_ram[576] = 147;
    exp_33_ram[577] = 179;
    exp_33_ram[578] = 99;
    exp_33_ram[579] = 147;
    exp_33_ram[580] = 19;
    exp_33_ram[581] = 179;
    exp_33_ram[582] = 19;
    exp_33_ram[583] = 103;
    exp_33_ram[584] = 51;
    exp_33_ram[585] = 179;
    exp_33_ram[586] = 51;
    exp_33_ram[587] = 179;
    exp_33_ram[588] = 111;
    exp_33_ram[589] = 183;
    exp_33_ram[590] = 99;
    exp_33_ram[591] = 147;
    exp_33_ram[592] = 179;
    exp_33_ram[593] = 147;
    exp_33_ram[594] = 55;
    exp_33_ram[595] = 147;
    exp_33_ram[596] = 179;
    exp_33_ram[597] = 51;
    exp_33_ram[598] = 147;
    exp_33_ram[599] = 51;
    exp_33_ram[600] = 3;
    exp_33_ram[601] = 51;
    exp_33_ram[602] = 103;
    exp_33_ram[603] = 55;
    exp_33_ram[604] = 147;
    exp_33_ram[605] = 227;
    exp_33_ram[606] = 147;
    exp_33_ram[607] = 111;
    exp_33_ram[608] = 115;
    exp_33_ram[609] = 109;
    exp_33_ram[610] = 46;
    exp_33_ram[611] = 112;
    exp_33_ram[612] = 10;
    exp_33_ram[613] = 116;
    exp_33_ram[614] = 46;
    exp_33_ram[615] = 84;
    exp_33_ram[616] = 83;
    exp_33_ram[617] = 49;
    exp_33_ram[618] = 48;
    exp_33_ram[619] = 58;
    exp_33_ram[620] = 50;
    exp_33_ram[621] = 10;
    exp_33_ram[622] = 49;
    exp_33_ram[623] = 105;
    exp_33_ram[624] = 84;
    exp_33_ram[625] = 83;
    exp_33_ram[626] = 49;
    exp_33_ram[627] = 49;
    exp_33_ram[628] = 58;
    exp_33_ram[629] = 50;
    exp_33_ram[630] = 10;
    exp_33_ram[631] = 50;
    exp_33_ram[632] = 105;
    exp_33_ram[633] = 51;
    exp_33_ram[634] = 105;
    exp_33_ram[635] = 52;
    exp_33_ram[636] = 105;
    exp_33_ram[637] = 53;
    exp_33_ram[638] = 105;
    exp_33_ram[639] = 54;
    exp_33_ram[640] = 105;
    exp_33_ram[641] = 55;
    exp_33_ram[642] = 105;
    exp_33_ram[643] = 56;
    exp_33_ram[644] = 105;
    exp_33_ram[645] = 57;
    exp_33_ram[646] = 105;
    exp_33_ram[647] = 84;
    exp_33_ram[648] = 83;
    exp_33_ram[649] = 49;
    exp_33_ram[650] = 50;
    exp_33_ram[651] = 58;
    exp_33_ram[652] = 50;
    exp_33_ram[653] = 10;
    exp_33_ram[654] = 49;
    exp_33_ram[655] = 97;
    exp_33_ram[656] = 49;
    exp_33_ram[657] = 97;
    exp_33_ram[658] = 49;
    exp_33_ram[659] = 97;
    exp_33_ram[660] = 112;
    exp_33_ram[661] = 0;
    exp_33_ram[662] = 0;
    exp_33_ram[663] = 3;
    exp_33_ram[664] = 4;
    exp_33_ram[665] = 4;
    exp_33_ram[666] = 5;
    exp_33_ram[667] = 5;
    exp_33_ram[668] = 5;
    exp_33_ram[669] = 5;
    exp_33_ram[670] = 6;
    exp_33_ram[671] = 6;
    exp_33_ram[672] = 6;
    exp_33_ram[673] = 6;
    exp_33_ram[674] = 6;
    exp_33_ram[675] = 6;
    exp_33_ram[676] = 6;
    exp_33_ram[677] = 6;
    exp_33_ram[678] = 7;
    exp_33_ram[679] = 7;
    exp_33_ram[680] = 7;
    exp_33_ram[681] = 7;
    exp_33_ram[682] = 7;
    exp_33_ram[683] = 7;
    exp_33_ram[684] = 7;
    exp_33_ram[685] = 7;
    exp_33_ram[686] = 7;
    exp_33_ram[687] = 7;
    exp_33_ram[688] = 7;
    exp_33_ram[689] = 7;
    exp_33_ram[690] = 7;
    exp_33_ram[691] = 7;
    exp_33_ram[692] = 7;
    exp_33_ram[693] = 7;
    exp_33_ram[694] = 8;
    exp_33_ram[695] = 8;
    exp_33_ram[696] = 8;
    exp_33_ram[697] = 8;
    exp_33_ram[698] = 8;
    exp_33_ram[699] = 8;
    exp_33_ram[700] = 8;
    exp_33_ram[701] = 8;
    exp_33_ram[702] = 8;
    exp_33_ram[703] = 8;
    exp_33_ram[704] = 8;
    exp_33_ram[705] = 8;
    exp_33_ram[706] = 8;
    exp_33_ram[707] = 8;
    exp_33_ram[708] = 8;
    exp_33_ram[709] = 8;
    exp_33_ram[710] = 8;
    exp_33_ram[711] = 8;
    exp_33_ram[712] = 8;
    exp_33_ram[713] = 8;
    exp_33_ram[714] = 8;
    exp_33_ram[715] = 8;
    exp_33_ram[716] = 8;
    exp_33_ram[717] = 8;
    exp_33_ram[718] = 8;
    exp_33_ram[719] = 8;
    exp_33_ram[720] = 8;
    exp_33_ram[721] = 8;
    exp_33_ram[722] = 8;
    exp_33_ram[723] = 8;
    exp_33_ram[724] = 8;
    exp_33_ram[725] = 8;
    exp_33_ram[726] = 147;
    exp_33_ram[727] = 19;
    exp_33_ram[728] = 51;
    exp_33_ram[729] = 3;
    exp_33_ram[730] = 99;
    exp_33_ram[731] = 103;
    exp_33_ram[732] = 19;
    exp_33_ram[733] = 35;
    exp_33_ram[734] = 111;
    exp_33_ram[735] = 19;
    exp_33_ram[736] = 183;
    exp_33_ram[737] = 35;
    exp_33_ram[738] = 3;
    exp_33_ram[739] = 35;
    exp_33_ram[740] = 147;
    exp_33_ram[741] = 239;
    exp_33_ram[742] = 147;
    exp_33_ram[743] = 131;
    exp_33_ram[744] = 35;
    exp_33_ram[745] = 3;
    exp_33_ram[746] = 19;
    exp_33_ram[747] = 19;
    exp_33_ram[748] = 103;
    exp_33_ram[749] = 179;
    exp_33_ram[750] = 147;
    exp_33_ram[751] = 147;
    exp_33_ram[752] = 99;
    exp_33_ram[753] = 19;
    exp_33_ram[754] = 51;
    exp_33_ram[755] = 19;
    exp_33_ram[756] = 111;
    exp_33_ram[757] = 131;
    exp_33_ram[758] = 19;
    exp_33_ram[759] = 147;
    exp_33_ram[760] = 35;
    exp_33_ram[761] = 131;
    exp_33_ram[762] = 35;
    exp_33_ram[763] = 131;
    exp_33_ram[764] = 35;
    exp_33_ram[765] = 131;
    exp_33_ram[766] = 35;
    exp_33_ram[767] = 179;
    exp_33_ram[768] = 227;
    exp_33_ram[769] = 19;
    exp_33_ram[770] = 19;
    exp_33_ram[771] = 179;
    exp_33_ram[772] = 179;
    exp_33_ram[773] = 19;
    exp_33_ram[774] = 51;
    exp_33_ram[775] = 99;
    exp_33_ram[776] = 19;
    exp_33_ram[777] = 19;
    exp_33_ram[778] = 179;
    exp_33_ram[779] = 179;
    exp_33_ram[780] = 147;
    exp_33_ram[781] = 99;
    exp_33_ram[782] = 103;
    exp_33_ram[783] = 51;
    exp_33_ram[784] = 131;
    exp_33_ram[785] = 51;
    exp_33_ram[786] = 147;
    exp_33_ram[787] = 35;
    exp_33_ram[788] = 111;
    exp_33_ram[789] = 51;
    exp_33_ram[790] = 3;
    exp_33_ram[791] = 51;
    exp_33_ram[792] = 147;
    exp_33_ram[793] = 35;
    exp_33_ram[794] = 111;
    exp_33_ram[795] = 179;
    exp_33_ram[796] = 147;
    exp_33_ram[797] = 99;
    exp_33_ram[798] = 183;
    exp_33_ram[799] = 55;
    exp_33_ram[800] = 147;
    exp_33_ram[801] = 19;
    exp_33_ram[802] = 3;
    exp_33_ram[803] = 131;
    exp_33_ram[804] = 99;
    exp_33_ram[805] = 131;
    exp_33_ram[806] = 3;
    exp_33_ram[807] = 99;
    exp_33_ram[808] = 99;
    exp_33_ram[809] = 51;
    exp_33_ram[810] = 103;
    exp_33_ram[811] = 51;
    exp_33_ram[812] = 147;
    exp_33_ram[813] = 179;
    exp_33_ram[814] = 179;
    exp_33_ram[815] = 99;
    exp_33_ram[816] = 19;
    exp_33_ram[817] = 147;
    exp_33_ram[818] = 111;
    exp_33_ram[819] = 19;
    exp_33_ram[820] = 147;
    exp_33_ram[821] = 111;
    exp_33_ram[822] = 19;
    exp_33_ram[823] = 103;
    exp_33_ram[824] = 147;
    exp_33_ram[825] = 99;
    exp_33_ram[826] = 19;
    exp_33_ram[827] = 147;
    exp_33_ram[828] = 35;
    exp_33_ram[829] = 35;
    exp_33_ram[830] = 19;
    exp_33_ram[831] = 239;
    exp_33_ram[832] = 147;
    exp_33_ram[833] = 99;
    exp_33_ram[834] = 147;
    exp_33_ram[835] = 19;
    exp_33_ram[836] = 239;
    exp_33_ram[837] = 147;
    exp_33_ram[838] = 131;
    exp_33_ram[839] = 3;
    exp_33_ram[840] = 19;
    exp_33_ram[841] = 19;
    exp_33_ram[842] = 103;
    exp_33_ram[843] = 147;
    exp_33_ram[844] = 19;
    exp_33_ram[845] = 103;
    exp_33_ram[846] = 147;
    exp_33_ram[847] = 147;
    exp_33_ram[848] = 99;
    exp_33_ram[849] = 19;
    exp_33_ram[850] = 147;
    exp_33_ram[851] = 147;
    exp_33_ram[852] = 99;
    exp_33_ram[853] = 19;
    exp_33_ram[854] = 147;
    exp_33_ram[855] = 99;
    exp_33_ram[856] = 19;
    exp_33_ram[857] = 35;
    exp_33_ram[858] = 239;
    exp_33_ram[859] = 131;
    exp_33_ram[860] = 179;
    exp_33_ram[861] = 147;
    exp_33_ram[862] = 19;
    exp_33_ram[863] = 19;
    exp_33_ram[864] = 103;
    exp_33_ram[865] = 147;
    exp_33_ram[866] = 19;
    exp_33_ram[867] = 103;
    exp_33_ram[868] = 183;
    exp_33_ram[869] = 3;
    exp_33_ram[870] = 131;
    exp_33_ram[871] = 131;
    exp_33_ram[872] = 19;
    exp_33_ram[873] = 131;
    exp_33_ram[874] = 179;
    exp_33_ram[875] = 103;
    exp_33_ram[876] = 147;
    exp_33_ram[877] = 51;
    exp_33_ram[878] = 179;
    exp_33_ram[879] = 179;
    exp_33_ram[880] = 19;
    exp_33_ram[881] = 179;
    exp_33_ram[882] = 35;
    exp_33_ram[883] = 239;
    exp_33_ram[884] = 131;
    exp_33_ram[885] = 19;
    exp_33_ram[886] = 103;
    exp_33_ram[887] = 19;
    exp_33_ram[888] = 35;
    exp_33_ram[889] = 131;
    exp_33_ram[890] = 35;
    exp_33_ram[891] = 183;
    exp_33_ram[892] = 35;
    exp_33_ram[893] = 35;
    exp_33_ram[894] = 35;
    exp_33_ram[895] = 35;
    exp_33_ram[896] = 35;
    exp_33_ram[897] = 35;
    exp_33_ram[898] = 19;
    exp_33_ram[899] = 19;
    exp_33_ram[900] = 19;
    exp_33_ram[901] = 147;
    exp_33_ram[902] = 147;
    exp_33_ram[903] = 147;
    exp_33_ram[904] = 99;
    exp_33_ram[905] = 3;
    exp_33_ram[906] = 183;
    exp_33_ram[907] = 147;
    exp_33_ram[908] = 147;
    exp_33_ram[909] = 99;
    exp_33_ram[910] = 147;
    exp_33_ram[911] = 19;
    exp_33_ram[912] = 239;
    exp_33_ram[913] = 147;
    exp_33_ram[914] = 239;
    exp_33_ram[915] = 51;
    exp_33_ram[916] = 179;
    exp_33_ram[917] = 179;
    exp_33_ram[918] = 19;
    exp_33_ram[919] = 147;
    exp_33_ram[920] = 111;
    exp_33_ram[921] = 19;
    exp_33_ram[922] = 239;
    exp_33_ram[923] = 51;
    exp_33_ram[924] = 147;
    exp_33_ram[925] = 19;
    exp_33_ram[926] = 239;
    exp_33_ram[927] = 51;
    exp_33_ram[928] = 179;
    exp_33_ram[929] = 179;
    exp_33_ram[930] = 19;
    exp_33_ram[931] = 19;
    exp_33_ram[932] = 111;
    exp_33_ram[933] = 3;
    exp_33_ram[934] = 3;
    exp_33_ram[935] = 131;
    exp_33_ram[936] = 147;
    exp_33_ram[937] = 179;
    exp_33_ram[938] = 147;
    exp_33_ram[939] = 179;
    exp_33_ram[940] = 19;
    exp_33_ram[941] = 51;
    exp_33_ram[942] = 147;
    exp_33_ram[943] = 19;
    exp_33_ram[944] = 3;
    exp_33_ram[945] = 19;
    exp_33_ram[946] = 147;
    exp_33_ram[947] = 51;
    exp_33_ram[948] = 179;
    exp_33_ram[949] = 179;
    exp_33_ram[950] = 179;
    exp_33_ram[951] = 183;
    exp_33_ram[952] = 147;
    exp_33_ram[953] = 179;
    exp_33_ram[954] = 51;
    exp_33_ram[955] = 179;
    exp_33_ram[956] = 147;
    exp_33_ram[957] = 19;
    exp_33_ram[958] = 51;
    exp_33_ram[959] = 239;
    exp_33_ram[960] = 179;
    exp_33_ram[961] = 147;
    exp_33_ram[962] = 179;
    exp_33_ram[963] = 179;
    exp_33_ram[964] = 51;
    exp_33_ram[965] = 51;
    exp_33_ram[966] = 51;
    exp_33_ram[967] = 179;
    exp_33_ram[968] = 131;
    exp_33_ram[969] = 179;
    exp_33_ram[970] = 3;
    exp_33_ram[971] = 131;
    exp_33_ram[972] = 3;
    exp_33_ram[973] = 131;
    exp_33_ram[974] = 3;
    exp_33_ram[975] = 131;
    exp_33_ram[976] = 3;
    exp_33_ram[977] = 19;
    exp_33_ram[978] = 103;
    exp_33_ram[979] = 19;
    exp_33_ram[980] = 35;
    exp_33_ram[981] = 35;
    exp_33_ram[982] = 19;
    exp_33_ram[983] = 239;
    exp_33_ram[984] = 183;
    exp_33_ram[985] = 3;
    exp_33_ram[986] = 147;
    exp_33_ram[987] = 239;
    exp_33_ram[988] = 183;
    exp_33_ram[989] = 131;
    exp_33_ram[990] = 51;
    exp_33_ram[991] = 99;
    exp_33_ram[992] = 35;
    exp_33_ram[993] = 35;
    exp_33_ram[994] = 131;
    exp_33_ram[995] = 3;
    exp_33_ram[996] = 147;
    exp_33_ram[997] = 19;
    exp_33_ram[998] = 103;
    exp_33_ram[999] = 19;
    exp_33_ram[1000] = 35;
    exp_33_ram[1001] = 35;
    exp_33_ram[1002] = 35;
    exp_33_ram[1003] = 35;
    exp_33_ram[1004] = 147;
    exp_33_ram[1005] = 19;
    exp_33_ram[1006] = 239;
    exp_33_ram[1007] = 183;
    exp_33_ram[1008] = 3;
    exp_33_ram[1009] = 147;
    exp_33_ram[1010] = 55;
    exp_33_ram[1011] = 239;
    exp_33_ram[1012] = 51;
    exp_33_ram[1013] = 179;
    exp_33_ram[1014] = 51;
    exp_33_ram[1015] = 19;
    exp_33_ram[1016] = 51;
    exp_33_ram[1017] = 35;
    exp_33_ram[1018] = 131;
    exp_33_ram[1019] = 3;
    exp_33_ram[1020] = 35;
    exp_33_ram[1021] = 131;
    exp_33_ram[1022] = 3;
    exp_33_ram[1023] = 19;
    exp_33_ram[1024] = 103;
    exp_33_ram[1025] = 19;
    exp_33_ram[1026] = 183;
    exp_33_ram[1027] = 35;
    exp_33_ram[1028] = 19;
    exp_33_ram[1029] = 147;
    exp_33_ram[1030] = 147;
    exp_33_ram[1031] = 19;
    exp_33_ram[1032] = 35;
    exp_33_ram[1033] = 35;
    exp_33_ram[1034] = 35;
    exp_33_ram[1035] = 35;
    exp_33_ram[1036] = 35;
    exp_33_ram[1037] = 239;
    exp_33_ram[1038] = 183;
    exp_33_ram[1039] = 19;
    exp_33_ram[1040] = 147;
    exp_33_ram[1041] = 19;
    exp_33_ram[1042] = 239;
    exp_33_ram[1043] = 131;
    exp_33_ram[1044] = 183;
    exp_33_ram[1045] = 19;
    exp_33_ram[1046] = 147;
    exp_33_ram[1047] = 179;
    exp_33_ram[1048] = 147;
    exp_33_ram[1049] = 19;
    exp_33_ram[1050] = 179;
    exp_33_ram[1051] = 19;
    exp_33_ram[1052] = 19;
    exp_33_ram[1053] = 239;
    exp_33_ram[1054] = 163;
    exp_33_ram[1055] = 131;
    exp_33_ram[1056] = 19;
    exp_33_ram[1057] = 19;
    exp_33_ram[1058] = 147;
    exp_33_ram[1059] = 179;
    exp_33_ram[1060] = 147;
    exp_33_ram[1061] = 179;
    exp_33_ram[1062] = 239;
    exp_33_ram[1063] = 163;
    exp_33_ram[1064] = 3;
    exp_33_ram[1065] = 147;
    exp_33_ram[1066] = 19;
    exp_33_ram[1067] = 239;
    exp_33_ram[1068] = 35;
    exp_33_ram[1069] = 131;
    exp_33_ram[1070] = 35;
    exp_33_ram[1071] = 35;
    exp_33_ram[1072] = 147;
    exp_33_ram[1073] = 35;
    exp_33_ram[1074] = 131;
    exp_33_ram[1075] = 147;
    exp_33_ram[1076] = 147;
    exp_33_ram[1077] = 163;
    exp_33_ram[1078] = 3;
    exp_33_ram[1079] = 239;
    exp_33_ram[1080] = 35;
    exp_33_ram[1081] = 131;
    exp_33_ram[1082] = 35;
    exp_33_ram[1083] = 163;
    exp_33_ram[1084] = 147;
    exp_33_ram[1085] = 163;
    exp_33_ram[1086] = 131;
    exp_33_ram[1087] = 147;
    exp_33_ram[1088] = 147;
    exp_33_ram[1089] = 35;
    exp_33_ram[1090] = 3;
    exp_33_ram[1091] = 239;
    exp_33_ram[1092] = 35;
    exp_33_ram[1093] = 131;
    exp_33_ram[1094] = 35;
    exp_33_ram[1095] = 35;
    exp_33_ram[1096] = 147;
    exp_33_ram[1097] = 35;
    exp_33_ram[1098] = 131;
    exp_33_ram[1099] = 147;
    exp_33_ram[1100] = 147;
    exp_33_ram[1101] = 163;
    exp_33_ram[1102] = 3;
    exp_33_ram[1103] = 239;
    exp_33_ram[1104] = 35;
    exp_33_ram[1105] = 131;
    exp_33_ram[1106] = 35;
    exp_33_ram[1107] = 163;
    exp_33_ram[1108] = 147;
    exp_33_ram[1109] = 163;
    exp_33_ram[1110] = 131;
    exp_33_ram[1111] = 147;
    exp_33_ram[1112] = 147;
    exp_33_ram[1113] = 35;
    exp_33_ram[1114] = 3;
    exp_33_ram[1115] = 19;
    exp_33_ram[1116] = 239;
    exp_33_ram[1117] = 35;
    exp_33_ram[1118] = 35;
    exp_33_ram[1119] = 131;
    exp_33_ram[1120] = 3;
    exp_33_ram[1121] = 147;
    exp_33_ram[1122] = 147;
    exp_33_ram[1123] = 35;
    exp_33_ram[1124] = 239;
    exp_33_ram[1125] = 35;
    exp_33_ram[1126] = 35;
    exp_33_ram[1127] = 131;
    exp_33_ram[1128] = 3;
    exp_33_ram[1129] = 147;
    exp_33_ram[1130] = 147;
    exp_33_ram[1131] = 163;
    exp_33_ram[1132] = 239;
    exp_33_ram[1133] = 35;
    exp_33_ram[1134] = 131;
    exp_33_ram[1135] = 35;
    exp_33_ram[1136] = 131;
    exp_33_ram[1137] = 147;
    exp_33_ram[1138] = 35;
    exp_33_ram[1139] = 131;
    exp_33_ram[1140] = 131;
    exp_33_ram[1141] = 3;
    exp_33_ram[1142] = 147;
    exp_33_ram[1143] = 163;
    exp_33_ram[1144] = 147;
    exp_33_ram[1145] = 35;
    exp_33_ram[1146] = 3;
    exp_33_ram[1147] = 3;
    exp_33_ram[1148] = 19;
    exp_33_ram[1149] = 131;
    exp_33_ram[1150] = 19;
    exp_33_ram[1151] = 103;
    exp_33_ram[1152] = 19;
    exp_33_ram[1153] = 35;
    exp_33_ram[1154] = 55;
    exp_33_ram[1155] = 35;
    exp_33_ram[1156] = 35;
    exp_33_ram[1157] = 35;
    exp_33_ram[1158] = 35;
    exp_33_ram[1159] = 35;
    exp_33_ram[1160] = 35;
    exp_33_ram[1161] = 35;
    exp_33_ram[1162] = 35;
    exp_33_ram[1163] = 35;
    exp_33_ram[1164] = 35;
    exp_33_ram[1165] = 19;
    exp_33_ram[1166] = 147;
    exp_33_ram[1167] = 19;
    exp_33_ram[1168] = 147;
    exp_33_ram[1169] = 147;
    exp_33_ram[1170] = 19;
    exp_33_ram[1171] = 19;
    exp_33_ram[1172] = 239;
    exp_33_ram[1173] = 51;
    exp_33_ram[1174] = 19;
    exp_33_ram[1175] = 147;
    exp_33_ram[1176] = 19;
    exp_33_ram[1177] = 239;
    exp_33_ram[1178] = 147;
    exp_33_ram[1179] = 99;
    exp_33_ram[1180] = 99;
    exp_33_ram[1181] = 51;
    exp_33_ram[1182] = 51;
    exp_33_ram[1183] = 179;
    exp_33_ram[1184] = 147;
    exp_33_ram[1185] = 51;
    exp_33_ram[1186] = 147;
    exp_33_ram[1187] = 111;
    exp_33_ram[1188] = 55;
    exp_33_ram[1189] = 147;
    exp_33_ram[1190] = 19;
    exp_33_ram[1191] = 19;
    exp_33_ram[1192] = 147;
    exp_33_ram[1193] = 19;
    exp_33_ram[1194] = 239;
    exp_33_ram[1195] = 147;
    exp_33_ram[1196] = 19;
    exp_33_ram[1197] = 147;
    exp_33_ram[1198] = 147;
    exp_33_ram[1199] = 239;
    exp_33_ram[1200] = 99;
    exp_33_ram[1201] = 99;
    exp_33_ram[1202] = 51;
    exp_33_ram[1203] = 179;
    exp_33_ram[1204] = 179;
    exp_33_ram[1205] = 51;
    exp_33_ram[1206] = 147;
    exp_33_ram[1207] = 51;
    exp_33_ram[1208] = 111;
    exp_33_ram[1209] = 183;
    exp_33_ram[1210] = 19;
    exp_33_ram[1211] = 147;
    exp_33_ram[1212] = 239;
    exp_33_ram[1213] = 35;
    exp_33_ram[1214] = 147;
    exp_33_ram[1215] = 35;
    exp_33_ram[1216] = 51;
    exp_33_ram[1217] = 3;
    exp_33_ram[1218] = 183;
    exp_33_ram[1219] = 147;
    exp_33_ram[1220] = 239;
    exp_33_ram[1221] = 35;
    exp_33_ram[1222] = 19;
    exp_33_ram[1223] = 35;
    exp_33_ram[1224] = 3;
    exp_33_ram[1225] = 147;
    exp_33_ram[1226] = 147;
    exp_33_ram[1227] = 239;
    exp_33_ram[1228] = 147;
    exp_33_ram[1229] = 35;
    exp_33_ram[1230] = 35;
    exp_33_ram[1231] = 35;
    exp_33_ram[1232] = 35;
    exp_33_ram[1233] = 35;
    exp_33_ram[1234] = 35;
    exp_33_ram[1235] = 35;
    exp_33_ram[1236] = 51;
    exp_33_ram[1237] = 35;
    exp_33_ram[1238] = 147;
    exp_33_ram[1239] = 239;
    exp_33_ram[1240] = 35;
    exp_33_ram[1241] = 35;
    exp_33_ram[1242] = 131;
    exp_33_ram[1243] = 19;
    exp_33_ram[1244] = 3;
    exp_33_ram[1245] = 131;
    exp_33_ram[1246] = 3;
    exp_33_ram[1247] = 131;
    exp_33_ram[1248] = 3;
    exp_33_ram[1249] = 131;
    exp_33_ram[1250] = 3;
    exp_33_ram[1251] = 131;
    exp_33_ram[1252] = 3;
    exp_33_ram[1253] = 131;
    exp_33_ram[1254] = 19;
    exp_33_ram[1255] = 103;
    exp_33_ram[1256] = 19;
    exp_33_ram[1257] = 35;
    exp_33_ram[1258] = 131;
    exp_33_ram[1259] = 147;
    exp_33_ram[1260] = 35;
    exp_33_ram[1261] = 35;
    exp_33_ram[1262] = 35;
    exp_33_ram[1263] = 147;
    exp_33_ram[1264] = 19;
    exp_33_ram[1265] = 19;
    exp_33_ram[1266] = 19;
    exp_33_ram[1267] = 147;
    exp_33_ram[1268] = 19;
    exp_33_ram[1269] = 35;
    exp_33_ram[1270] = 35;
    exp_33_ram[1271] = 35;
    exp_33_ram[1272] = 35;
    exp_33_ram[1273] = 35;
    exp_33_ram[1274] = 35;
    exp_33_ram[1275] = 35;
    exp_33_ram[1276] = 35;
    exp_33_ram[1277] = 35;
    exp_33_ram[1278] = 35;
    exp_33_ram[1279] = 239;
    exp_33_ram[1280] = 19;
    exp_33_ram[1281] = 239;
    exp_33_ram[1282] = 19;
    exp_33_ram[1283] = 147;
    exp_33_ram[1284] = 19;
    exp_33_ram[1285] = 239;
    exp_33_ram[1286] = 3;
    exp_33_ram[1287] = 131;
    exp_33_ram[1288] = 19;
    exp_33_ram[1289] = 147;
    exp_33_ram[1290] = 179;
    exp_33_ram[1291] = 19;
    exp_33_ram[1292] = 35;
    exp_33_ram[1293] = 239;
    exp_33_ram[1294] = 19;
    exp_33_ram[1295] = 239;
    exp_33_ram[1296] = 147;
    exp_33_ram[1297] = 19;
    exp_33_ram[1298] = 147;
    exp_33_ram[1299] = 19;
    exp_33_ram[1300] = 19;
    exp_33_ram[1301] = 147;
    exp_33_ram[1302] = 35;
    exp_33_ram[1303] = 35;
    exp_33_ram[1304] = 35;
    exp_33_ram[1305] = 35;
    exp_33_ram[1306] = 35;
    exp_33_ram[1307] = 35;
    exp_33_ram[1308] = 239;
    exp_33_ram[1309] = 19;
    exp_33_ram[1310] = 239;
    exp_33_ram[1311] = 19;
    exp_33_ram[1312] = 147;
    exp_33_ram[1313] = 19;
    exp_33_ram[1314] = 239;
    exp_33_ram[1315] = 3;
    exp_33_ram[1316] = 131;
    exp_33_ram[1317] = 19;
    exp_33_ram[1318] = 147;
    exp_33_ram[1319] = 179;
    exp_33_ram[1320] = 19;
    exp_33_ram[1321] = 35;
    exp_33_ram[1322] = 239;
    exp_33_ram[1323] = 19;
    exp_33_ram[1324] = 239;
    exp_33_ram[1325] = 147;
    exp_33_ram[1326] = 19;
    exp_33_ram[1327] = 19;
    exp_33_ram[1328] = 147;
    exp_33_ram[1329] = 19;
    exp_33_ram[1330] = 239;
    exp_33_ram[1331] = 19;
    exp_33_ram[1332] = 239;
    exp_33_ram[1333] = 99;
    exp_33_ram[1334] = 19;
    exp_33_ram[1335] = 147;
    exp_33_ram[1336] = 99;
    exp_33_ram[1337] = 99;
    exp_33_ram[1338] = 19;
    exp_33_ram[1339] = 99;
    exp_33_ram[1340] = 99;
    exp_33_ram[1341] = 99;
    exp_33_ram[1342] = 19;
    exp_33_ram[1343] = 131;
    exp_33_ram[1344] = 3;
    exp_33_ram[1345] = 131;
    exp_33_ram[1346] = 3;
    exp_33_ram[1347] = 131;
    exp_33_ram[1348] = 3;
    exp_33_ram[1349] = 131;
    exp_33_ram[1350] = 19;
    exp_33_ram[1351] = 103;
    exp_33_ram[1352] = 19;
    exp_33_ram[1353] = 147;
    exp_33_ram[1354] = 35;
    exp_33_ram[1355] = 19;
    exp_33_ram[1356] = 19;
    exp_33_ram[1357] = 19;
    exp_33_ram[1358] = 35;
    exp_33_ram[1359] = 35;
    exp_33_ram[1360] = 35;
    exp_33_ram[1361] = 35;
    exp_33_ram[1362] = 239;
    exp_33_ram[1363] = 19;
    exp_33_ram[1364] = 147;
    exp_33_ram[1365] = 19;
    exp_33_ram[1366] = 131;
    exp_33_ram[1367] = 239;
    exp_33_ram[1368] = 19;
    exp_33_ram[1369] = 239;
    exp_33_ram[1370] = 147;
    exp_33_ram[1371] = 19;
    exp_33_ram[1372] = 99;
    exp_33_ram[1373] = 183;
    exp_33_ram[1374] = 147;
    exp_33_ram[1375] = 179;
    exp_33_ram[1376] = 51;
    exp_33_ram[1377] = 19;
    exp_33_ram[1378] = 147;
    exp_33_ram[1379] = 51;
    exp_33_ram[1380] = 147;
    exp_33_ram[1381] = 19;
    exp_33_ram[1382] = 19;
    exp_33_ram[1383] = 239;
    exp_33_ram[1384] = 19;
    exp_33_ram[1385] = 147;
    exp_33_ram[1386] = 19;
    exp_33_ram[1387] = 239;
    exp_33_ram[1388] = 99;
    exp_33_ram[1389] = 147;
    exp_33_ram[1390] = 35;
    exp_33_ram[1391] = 131;
    exp_33_ram[1392] = 147;
    exp_33_ram[1393] = 3;
    exp_33_ram[1394] = 3;
    exp_33_ram[1395] = 131;
    exp_33_ram[1396] = 19;
    exp_33_ram[1397] = 131;
    exp_33_ram[1398] = 19;
    exp_33_ram[1399] = 103;
    exp_33_ram[1400] = 227;
    exp_33_ram[1401] = 19;
    exp_33_ram[1402] = 147;
    exp_33_ram[1403] = 19;
    exp_33_ram[1404] = 239;
    exp_33_ram[1405] = 19;
    exp_33_ram[1406] = 239;
    exp_33_ram[1407] = 147;
    exp_33_ram[1408] = 99;
    exp_33_ram[1409] = 183;
    exp_33_ram[1410] = 147;
    exp_33_ram[1411] = 179;
    exp_33_ram[1412] = 51;
    exp_33_ram[1413] = 51;
    exp_33_ram[1414] = 147;
    exp_33_ram[1415] = 111;
    exp_33_ram[1416] = 99;
    exp_33_ram[1417] = 19;
    exp_33_ram[1418] = 147;
    exp_33_ram[1419] = 19;
    exp_33_ram[1420] = 239;
    exp_33_ram[1421] = 19;
    exp_33_ram[1422] = 239;
    exp_33_ram[1423] = 35;
    exp_33_ram[1424] = 111;
    exp_33_ram[1425] = 35;
    exp_33_ram[1426] = 111;
    exp_33_ram[1427] = 19;
    exp_33_ram[1428] = 19;
    exp_33_ram[1429] = 147;
    exp_33_ram[1430] = 19;
    exp_33_ram[1431] = 35;
    exp_33_ram[1432] = 239;
    exp_33_ram[1433] = 147;
    exp_33_ram[1434] = 19;
    exp_33_ram[1435] = 19;
    exp_33_ram[1436] = 239;
    exp_33_ram[1437] = 19;
    exp_33_ram[1438] = 239;
    exp_33_ram[1439] = 131;
    exp_33_ram[1440] = 19;
    exp_33_ram[1441] = 103;
    exp_33_ram[1442] = 131;
    exp_33_ram[1443] = 3;
    exp_33_ram[1444] = 19;
    exp_33_ram[1445] = 19;
    exp_33_ram[1446] = 35;
    exp_33_ram[1447] = 35;
    exp_33_ram[1448] = 239;
    exp_33_ram[1449] = 55;
    exp_33_ram[1450] = 147;
    exp_33_ram[1451] = 19;
    exp_33_ram[1452] = 19;
    exp_33_ram[1453] = 239;
    exp_33_ram[1454] = 131;
    exp_33_ram[1455] = 19;
    exp_33_ram[1456] = 3;
    exp_33_ram[1457] = 19;
    exp_33_ram[1458] = 103;
    exp_33_ram[1459] = 19;
    exp_33_ram[1460] = 35;
    exp_33_ram[1461] = 35;
    exp_33_ram[1462] = 131;
    exp_33_ram[1463] = 3;
    exp_33_ram[1464] = 35;
    exp_33_ram[1465] = 147;
    exp_33_ram[1466] = 19;
    exp_33_ram[1467] = 35;
    exp_33_ram[1468] = 35;
    exp_33_ram[1469] = 239;
    exp_33_ram[1470] = 19;
    exp_33_ram[1471] = 99;
    exp_33_ram[1472] = 55;
    exp_33_ram[1473] = 19;
    exp_33_ram[1474] = 179;
    exp_33_ram[1475] = 51;
    exp_33_ram[1476] = 51;
    exp_33_ram[1477] = 19;
    exp_33_ram[1478] = 239;
    exp_33_ram[1479] = 55;
    exp_33_ram[1480] = 147;
    exp_33_ram[1481] = 19;
    exp_33_ram[1482] = 19;
    exp_33_ram[1483] = 239;
    exp_33_ram[1484] = 19;
    exp_33_ram[1485] = 147;
    exp_33_ram[1486] = 239;
    exp_33_ram[1487] = 147;
    exp_33_ram[1488] = 35;
    exp_33_ram[1489] = 131;
    exp_33_ram[1490] = 19;
    exp_33_ram[1491] = 3;
    exp_33_ram[1492] = 131;
    exp_33_ram[1493] = 3;
    exp_33_ram[1494] = 131;
    exp_33_ram[1495] = 19;
    exp_33_ram[1496] = 103;
    exp_33_ram[1497] = 19;
    exp_33_ram[1498] = 35;
    exp_33_ram[1499] = 239;
    exp_33_ram[1500] = 131;
    exp_33_ram[1501] = 19;
    exp_33_ram[1502] = 111;
    exp_33_ram[1503] = 19;
    exp_33_ram[1504] = 35;
    exp_33_ram[1505] = 35;
    exp_33_ram[1506] = 19;
    exp_33_ram[1507] = 183;
    exp_33_ram[1508] = 19;
    exp_33_ram[1509] = 239;
    exp_33_ram[1510] = 183;
    exp_33_ram[1511] = 19;
    exp_33_ram[1512] = 239;
    exp_33_ram[1513] = 131;
    exp_33_ram[1514] = 3;
    exp_33_ram[1515] = 19;
    exp_33_ram[1516] = 103;
    exp_33_ram[1517] = 19;
    exp_33_ram[1518] = 35;
    exp_33_ram[1519] = 35;
    exp_33_ram[1520] = 35;
    exp_33_ram[1521] = 35;
    exp_33_ram[1522] = 35;
    exp_33_ram[1523] = 35;
    exp_33_ram[1524] = 35;
    exp_33_ram[1525] = 35;
    exp_33_ram[1526] = 19;
    exp_33_ram[1527] = 183;
    exp_33_ram[1528] = 19;
    exp_33_ram[1529] = 239;
    exp_33_ram[1530] = 147;
    exp_33_ram[1531] = 35;
    exp_33_ram[1532] = 147;
    exp_33_ram[1533] = 35;
    exp_33_ram[1534] = 147;
    exp_33_ram[1535] = 35;
    exp_33_ram[1536] = 147;
    exp_33_ram[1537] = 35;
    exp_33_ram[1538] = 147;
    exp_33_ram[1539] = 35;
    exp_33_ram[1540] = 35;
    exp_33_ram[1541] = 147;
    exp_33_ram[1542] = 35;
    exp_33_ram[1543] = 147;
    exp_33_ram[1544] = 19;
    exp_33_ram[1545] = 239;
    exp_33_ram[1546] = 19;
    exp_33_ram[1547] = 147;
    exp_33_ram[1548] = 35;
    exp_33_ram[1549] = 35;
    exp_33_ram[1550] = 147;
    exp_33_ram[1551] = 19;
    exp_33_ram[1552] = 239;
    exp_33_ram[1553] = 19;
    exp_33_ram[1554] = 183;
    exp_33_ram[1555] = 147;
    exp_33_ram[1556] = 19;
    exp_33_ram[1557] = 239;
    exp_33_ram[1558] = 147;
    exp_33_ram[1559] = 99;
    exp_33_ram[1560] = 183;
    exp_33_ram[1561] = 19;
    exp_33_ram[1562] = 239;
    exp_33_ram[1563] = 111;
    exp_33_ram[1564] = 147;
    exp_33_ram[1565] = 19;
    exp_33_ram[1566] = 239;
    exp_33_ram[1567] = 147;
    exp_33_ram[1568] = 19;
    exp_33_ram[1569] = 239;
    exp_33_ram[1570] = 19;
    exp_33_ram[1571] = 183;
    exp_33_ram[1572] = 147;
    exp_33_ram[1573] = 19;
    exp_33_ram[1574] = 239;
    exp_33_ram[1575] = 147;
    exp_33_ram[1576] = 99;
    exp_33_ram[1577] = 183;
    exp_33_ram[1578] = 19;
    exp_33_ram[1579] = 239;
    exp_33_ram[1580] = 111;
    exp_33_ram[1581] = 147;
    exp_33_ram[1582] = 19;
    exp_33_ram[1583] = 239;
    exp_33_ram[1584] = 147;
    exp_33_ram[1585] = 19;
    exp_33_ram[1586] = 239;
    exp_33_ram[1587] = 19;
    exp_33_ram[1588] = 183;
    exp_33_ram[1589] = 147;
    exp_33_ram[1590] = 19;
    exp_33_ram[1591] = 239;
    exp_33_ram[1592] = 147;
    exp_33_ram[1593] = 99;
    exp_33_ram[1594] = 183;
    exp_33_ram[1595] = 19;
    exp_33_ram[1596] = 239;
    exp_33_ram[1597] = 111;
    exp_33_ram[1598] = 147;
    exp_33_ram[1599] = 19;
    exp_33_ram[1600] = 239;
    exp_33_ram[1601] = 19;
    exp_33_ram[1602] = 183;
    exp_33_ram[1603] = 147;
    exp_33_ram[1604] = 19;
    exp_33_ram[1605] = 239;
    exp_33_ram[1606] = 147;
    exp_33_ram[1607] = 99;
    exp_33_ram[1608] = 183;
    exp_33_ram[1609] = 19;
    exp_33_ram[1610] = 239;
    exp_33_ram[1611] = 111;
    exp_33_ram[1612] = 147;
    exp_33_ram[1613] = 35;
    exp_33_ram[1614] = 147;
    exp_33_ram[1615] = 35;
    exp_33_ram[1616] = 147;
    exp_33_ram[1617] = 35;
    exp_33_ram[1618] = 147;
    exp_33_ram[1619] = 35;
    exp_33_ram[1620] = 147;
    exp_33_ram[1621] = 35;
    exp_33_ram[1622] = 35;
    exp_33_ram[1623] = 147;
    exp_33_ram[1624] = 35;
    exp_33_ram[1625] = 147;
    exp_33_ram[1626] = 19;
    exp_33_ram[1627] = 239;
    exp_33_ram[1628] = 19;
    exp_33_ram[1629] = 147;
    exp_33_ram[1630] = 35;
    exp_33_ram[1631] = 35;
    exp_33_ram[1632] = 147;
    exp_33_ram[1633] = 19;
    exp_33_ram[1634] = 239;
    exp_33_ram[1635] = 19;
    exp_33_ram[1636] = 183;
    exp_33_ram[1637] = 147;
    exp_33_ram[1638] = 19;
    exp_33_ram[1639] = 239;
    exp_33_ram[1640] = 147;
    exp_33_ram[1641] = 99;
    exp_33_ram[1642] = 183;
    exp_33_ram[1643] = 19;
    exp_33_ram[1644] = 239;
    exp_33_ram[1645] = 111;
    exp_33_ram[1646] = 147;
    exp_33_ram[1647] = 19;
    exp_33_ram[1648] = 239;
    exp_33_ram[1649] = 147;
    exp_33_ram[1650] = 19;
    exp_33_ram[1651] = 239;
    exp_33_ram[1652] = 19;
    exp_33_ram[1653] = 183;
    exp_33_ram[1654] = 147;
    exp_33_ram[1655] = 19;
    exp_33_ram[1656] = 239;
    exp_33_ram[1657] = 147;
    exp_33_ram[1658] = 99;
    exp_33_ram[1659] = 183;
    exp_33_ram[1660] = 19;
    exp_33_ram[1661] = 239;
    exp_33_ram[1662] = 111;
    exp_33_ram[1663] = 147;
    exp_33_ram[1664] = 19;
    exp_33_ram[1665] = 239;
    exp_33_ram[1666] = 147;
    exp_33_ram[1667] = 19;
    exp_33_ram[1668] = 239;
    exp_33_ram[1669] = 19;
    exp_33_ram[1670] = 183;
    exp_33_ram[1671] = 147;
    exp_33_ram[1672] = 19;
    exp_33_ram[1673] = 239;
    exp_33_ram[1674] = 147;
    exp_33_ram[1675] = 99;
    exp_33_ram[1676] = 183;
    exp_33_ram[1677] = 19;
    exp_33_ram[1678] = 239;
    exp_33_ram[1679] = 111;
    exp_33_ram[1680] = 147;
    exp_33_ram[1681] = 19;
    exp_33_ram[1682] = 239;
    exp_33_ram[1683] = 19;
    exp_33_ram[1684] = 183;
    exp_33_ram[1685] = 147;
    exp_33_ram[1686] = 19;
    exp_33_ram[1687] = 239;
    exp_33_ram[1688] = 147;
    exp_33_ram[1689] = 99;
    exp_33_ram[1690] = 183;
    exp_33_ram[1691] = 19;
    exp_33_ram[1692] = 239;
    exp_33_ram[1693] = 111;
    exp_33_ram[1694] = 147;
    exp_33_ram[1695] = 35;
    exp_33_ram[1696] = 147;
    exp_33_ram[1697] = 35;
    exp_33_ram[1698] = 147;
    exp_33_ram[1699] = 35;
    exp_33_ram[1700] = 147;
    exp_33_ram[1701] = 35;
    exp_33_ram[1702] = 147;
    exp_33_ram[1703] = 35;
    exp_33_ram[1704] = 35;
    exp_33_ram[1705] = 35;
    exp_33_ram[1706] = 147;
    exp_33_ram[1707] = 19;
    exp_33_ram[1708] = 239;
    exp_33_ram[1709] = 19;
    exp_33_ram[1710] = 147;
    exp_33_ram[1711] = 35;
    exp_33_ram[1712] = 35;
    exp_33_ram[1713] = 147;
    exp_33_ram[1714] = 19;
    exp_33_ram[1715] = 239;
    exp_33_ram[1716] = 19;
    exp_33_ram[1717] = 183;
    exp_33_ram[1718] = 147;
    exp_33_ram[1719] = 19;
    exp_33_ram[1720] = 239;
    exp_33_ram[1721] = 147;
    exp_33_ram[1722] = 99;
    exp_33_ram[1723] = 183;
    exp_33_ram[1724] = 19;
    exp_33_ram[1725] = 239;
    exp_33_ram[1726] = 111;
    exp_33_ram[1727] = 147;
    exp_33_ram[1728] = 19;
    exp_33_ram[1729] = 239;
    exp_33_ram[1730] = 147;
    exp_33_ram[1731] = 19;
    exp_33_ram[1732] = 239;
    exp_33_ram[1733] = 19;
    exp_33_ram[1734] = 183;
    exp_33_ram[1735] = 147;
    exp_33_ram[1736] = 19;
    exp_33_ram[1737] = 239;
    exp_33_ram[1738] = 147;
    exp_33_ram[1739] = 99;
    exp_33_ram[1740] = 183;
    exp_33_ram[1741] = 19;
    exp_33_ram[1742] = 239;
    exp_33_ram[1743] = 111;
    exp_33_ram[1744] = 147;
    exp_33_ram[1745] = 19;
    exp_33_ram[1746] = 239;
    exp_33_ram[1747] = 147;
    exp_33_ram[1748] = 19;
    exp_33_ram[1749] = 239;
    exp_33_ram[1750] = 19;
    exp_33_ram[1751] = 183;
    exp_33_ram[1752] = 147;
    exp_33_ram[1753] = 19;
    exp_33_ram[1754] = 239;
    exp_33_ram[1755] = 147;
    exp_33_ram[1756] = 99;
    exp_33_ram[1757] = 183;
    exp_33_ram[1758] = 19;
    exp_33_ram[1759] = 239;
    exp_33_ram[1760] = 111;
    exp_33_ram[1761] = 147;
    exp_33_ram[1762] = 19;
    exp_33_ram[1763] = 239;
    exp_33_ram[1764] = 19;
    exp_33_ram[1765] = 183;
    exp_33_ram[1766] = 147;
    exp_33_ram[1767] = 19;
    exp_33_ram[1768] = 239;
    exp_33_ram[1769] = 147;
    exp_33_ram[1770] = 99;
    exp_33_ram[1771] = 183;
    exp_33_ram[1772] = 19;
    exp_33_ram[1773] = 239;
    exp_33_ram[1774] = 111;
    exp_33_ram[1775] = 183;
    exp_33_ram[1776] = 19;
    exp_33_ram[1777] = 239;
    exp_33_ram[1778] = 147;
    exp_33_ram[1779] = 35;
    exp_33_ram[1780] = 147;
    exp_33_ram[1781] = 35;
    exp_33_ram[1782] = 147;
    exp_33_ram[1783] = 35;
    exp_33_ram[1784] = 35;
    exp_33_ram[1785] = 147;
    exp_33_ram[1786] = 35;
    exp_33_ram[1787] = 147;
    exp_33_ram[1788] = 35;
    exp_33_ram[1789] = 147;
    exp_33_ram[1790] = 35;
    exp_33_ram[1791] = 147;
    exp_33_ram[1792] = 19;
    exp_33_ram[1793] = 239;
    exp_33_ram[1794] = 19;
    exp_33_ram[1795] = 147;
    exp_33_ram[1796] = 35;
    exp_33_ram[1797] = 35;
    exp_33_ram[1798] = 3;
    exp_33_ram[1799] = 131;
    exp_33_ram[1800] = 19;
    exp_33_ram[1801] = 147;
    exp_33_ram[1802] = 239;
    exp_33_ram[1803] = 239;
    exp_33_ram[1804] = 35;
    exp_33_ram[1805] = 35;
    exp_33_ram[1806] = 35;
    exp_33_ram[1807] = 111;
    exp_33_ram[1808] = 19;
    exp_33_ram[1809] = 239;
    exp_33_ram[1810] = 19;
    exp_33_ram[1811] = 147;
    exp_33_ram[1812] = 3;
    exp_33_ram[1813] = 131;
    exp_33_ram[1814] = 19;
    exp_33_ram[1815] = 147;
    exp_33_ram[1816] = 239;
    exp_33_ram[1817] = 19;
    exp_33_ram[1818] = 147;
    exp_33_ram[1819] = 183;
    exp_33_ram[1820] = 131;
    exp_33_ram[1821] = 19;
    exp_33_ram[1822] = 239;
    exp_33_ram[1823] = 19;
    exp_33_ram[1824] = 147;
    exp_33_ram[1825] = 19;
    exp_33_ram[1826] = 147;
    exp_33_ram[1827] = 19;
    exp_33_ram[1828] = 147;
    exp_33_ram[1829] = 239;
    exp_33_ram[1830] = 147;
    exp_33_ram[1831] = 227;
    exp_33_ram[1832] = 183;
    exp_33_ram[1833] = 131;
    exp_33_ram[1834] = 19;
    exp_33_ram[1835] = 147;
    exp_33_ram[1836] = 3;
    exp_33_ram[1837] = 131;
    exp_33_ram[1838] = 51;
    exp_33_ram[1839] = 147;
    exp_33_ram[1840] = 179;
    exp_33_ram[1841] = 179;
    exp_33_ram[1842] = 179;
    exp_33_ram[1843] = 147;
    exp_33_ram[1844] = 35;
    exp_33_ram[1845] = 35;
    exp_33_ram[1846] = 19;
    exp_33_ram[1847] = 239;
    exp_33_ram[1848] = 19;
    exp_33_ram[1849] = 147;
    exp_33_ram[1850] = 35;
    exp_33_ram[1851] = 35;
    exp_33_ram[1852] = 147;
    exp_33_ram[1853] = 19;
    exp_33_ram[1854] = 239;
    exp_33_ram[1855] = 147;
    exp_33_ram[1856] = 19;
    exp_33_ram[1857] = 239;
    exp_33_ram[1858] = 131;
    exp_33_ram[1859] = 147;
    exp_33_ram[1860] = 35;
    exp_33_ram[1861] = 3;
    exp_33_ram[1862] = 147;
    exp_33_ram[1863] = 227;
    exp_33_ram[1864] = 147;
    exp_33_ram[1865] = 35;
    exp_33_ram[1866] = 147;
    exp_33_ram[1867] = 35;
    exp_33_ram[1868] = 147;
    exp_33_ram[1869] = 35;
    exp_33_ram[1870] = 147;
    exp_33_ram[1871] = 35;
    exp_33_ram[1872] = 147;
    exp_33_ram[1873] = 35;
    exp_33_ram[1874] = 147;
    exp_33_ram[1875] = 35;
    exp_33_ram[1876] = 147;
    exp_33_ram[1877] = 35;
    exp_33_ram[1878] = 147;
    exp_33_ram[1879] = 19;
    exp_33_ram[1880] = 239;
    exp_33_ram[1881] = 19;
    exp_33_ram[1882] = 147;
    exp_33_ram[1883] = 35;
    exp_33_ram[1884] = 35;
    exp_33_ram[1885] = 147;
    exp_33_ram[1886] = 19;
    exp_33_ram[1887] = 239;
    exp_33_ram[1888] = 147;
    exp_33_ram[1889] = 19;
    exp_33_ram[1890] = 239;
    exp_33_ram[1891] = 147;
    exp_33_ram[1892] = 19;
    exp_33_ram[1893] = 239;
    exp_33_ram[1894] = 147;
    exp_33_ram[1895] = 19;
    exp_33_ram[1896] = 239;
    exp_33_ram[1897] = 3;
    exp_33_ram[1898] = 131;
    exp_33_ram[1899] = 19;
    exp_33_ram[1900] = 147;
    exp_33_ram[1901] = 239;
    exp_33_ram[1902] = 19;
    exp_33_ram[1903] = 239;
    exp_33_ram[1904] = 19;
    exp_33_ram[1905] = 147;
    exp_33_ram[1906] = 35;
    exp_33_ram[1907] = 35;
    exp_33_ram[1908] = 147;
    exp_33_ram[1909] = 19;
    exp_33_ram[1910] = 239;
    exp_33_ram[1911] = 147;
    exp_33_ram[1912] = 19;
    exp_33_ram[1913] = 239;
    exp_33_ram[1914] = 239;
    exp_33_ram[1915] = 35;
    exp_33_ram[1916] = 35;
    exp_33_ram[1917] = 35;
    exp_33_ram[1918] = 111;
    exp_33_ram[1919] = 19;
    exp_33_ram[1920] = 239;
    exp_33_ram[1921] = 19;
    exp_33_ram[1922] = 147;
    exp_33_ram[1923] = 3;
    exp_33_ram[1924] = 131;
    exp_33_ram[1925] = 19;
    exp_33_ram[1926] = 147;
    exp_33_ram[1927] = 239;
    exp_33_ram[1928] = 19;
    exp_33_ram[1929] = 147;
    exp_33_ram[1930] = 183;
    exp_33_ram[1931] = 131;
    exp_33_ram[1932] = 19;
    exp_33_ram[1933] = 239;
    exp_33_ram[1934] = 19;
    exp_33_ram[1935] = 147;
    exp_33_ram[1936] = 19;
    exp_33_ram[1937] = 147;
    exp_33_ram[1938] = 19;
    exp_33_ram[1939] = 147;
    exp_33_ram[1940] = 239;
    exp_33_ram[1941] = 147;
    exp_33_ram[1942] = 227;
    exp_33_ram[1943] = 183;
    exp_33_ram[1944] = 131;
    exp_33_ram[1945] = 19;
    exp_33_ram[1946] = 147;
    exp_33_ram[1947] = 3;
    exp_33_ram[1948] = 131;
    exp_33_ram[1949] = 51;
    exp_33_ram[1950] = 147;
    exp_33_ram[1951] = 179;
    exp_33_ram[1952] = 179;
    exp_33_ram[1953] = 179;
    exp_33_ram[1954] = 147;
    exp_33_ram[1955] = 35;
    exp_33_ram[1956] = 35;
    exp_33_ram[1957] = 19;
    exp_33_ram[1958] = 239;
    exp_33_ram[1959] = 19;
    exp_33_ram[1960] = 147;
    exp_33_ram[1961] = 35;
    exp_33_ram[1962] = 35;
    exp_33_ram[1963] = 147;
    exp_33_ram[1964] = 19;
    exp_33_ram[1965] = 239;
    exp_33_ram[1966] = 147;
    exp_33_ram[1967] = 19;
    exp_33_ram[1968] = 239;
    exp_33_ram[1969] = 131;
    exp_33_ram[1970] = 147;
    exp_33_ram[1971] = 35;
    exp_33_ram[1972] = 3;
    exp_33_ram[1973] = 147;
    exp_33_ram[1974] = 227;
    exp_33_ram[1975] = 131;
    exp_33_ram[1976] = 3;
    exp_33_ram[1977] = 3;
    exp_33_ram[1978] = 131;
    exp_33_ram[1979] = 3;
    exp_33_ram[1980] = 131;
    exp_33_ram[1981] = 3;
    exp_33_ram[1982] = 131;
    exp_33_ram[1983] = 19;
    exp_33_ram[1984] = 103;
    exp_33_ram[1985] = 19;
    exp_33_ram[1986] = 35;
    exp_33_ram[1987] = 35;
    exp_33_ram[1988] = 19;
    exp_33_ram[1989] = 239;
    exp_33_ram[1990] = 239;
    exp_33_ram[1991] = 19;
    exp_33_ram[1992] = 131;
    exp_33_ram[1993] = 3;
    exp_33_ram[1994] = 19;
    exp_33_ram[1995] = 103;
    exp_33_ram[1996] = 19;
    exp_33_ram[1997] = 147;
    exp_33_ram[1998] = 51;
    exp_33_ram[1999] = 19;
    exp_33_ram[2000] = 179;
    exp_33_ram[2001] = 99;
    exp_33_ram[2002] = 99;
    exp_33_ram[2003] = 19;
    exp_33_ram[2004] = 179;
    exp_33_ram[2005] = 19;
    exp_33_ram[2006] = 103;
    exp_33_ram[2007] = 227;
    exp_33_ram[2008] = 19;
    exp_33_ram[2009] = 179;
    exp_33_ram[2010] = 111;
    exp_33_ram[2011] = 128;
    exp_33_ram[2012] = 8;
    exp_33_ram[2013] = 83;
    exp_33_ram[2014] = 111;
    exp_33_ram[2015] = 101;
    exp_33_ram[2016] = 84;
    exp_33_ram[2017] = 114;
    exp_33_ram[2018] = 116;
    exp_33_ram[2019] = 74;
    exp_33_ram[2020] = 101;
    exp_33_ram[2021] = 114;
    exp_33_ram[2022] = 77;
    exp_33_ram[2023] = 117;
    exp_33_ram[2024] = 108;
    exp_33_ram[2025] = 83;
    exp_33_ram[2026] = 99;
    exp_33_ram[2027] = 118;
    exp_33_ram[2028] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_31) begin
      exp_33_ram[exp_27] <= exp_29;
    end
  end
  assign exp_33 = exp_33_ram[exp_28];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_59) begin
        exp_33_ram[exp_55] <= exp_57;
    end
  end
  assign exp_61 = exp_33_ram[exp_56];
  assign exp_60 = exp_92;
  assign exp_92 = 1;
  assign exp_56 = exp_91;
  assign exp_91 = exp_8[31:2];
  assign exp_59 = exp_84;
  assign exp_55 = exp_83;
  assign exp_57 = exp_83;
  assign exp_32 = exp_127;
  assign exp_127 = 1;
  assign exp_28 = exp_126;
  assign exp_126 = exp_10[31:2];
  assign exp_31 = exp_101;
  assign exp_101 = exp_99 & exp_100;
  assign exp_99 = exp_14 & exp_15;
  assign exp_100 = exp_16[0:0];
  assign exp_27 = exp_97;
  assign exp_97 = exp_10[31:2];
  assign exp_29 = exp_98;
  assign exp_98 = exp_11[7:0];
  assign exp_118 = 1;
  assign exp_141 = exp_179;

  reg [31:0] exp_179_reg;
  always@(*) begin
    case (exp_177)
      0:exp_179_reg <= exp_157;
      1:exp_179_reg <= exp_167;
      default:exp_179_reg <= exp_178;
    endcase
  end
  assign exp_179 = exp_179_reg;
  assign exp_177 = exp_139[2:2];
  assign exp_139 = exp_1;
  assign exp_178 = 0;

      reg [31:0] exp_157_reg = 0;
      always@(posedge clk) begin
        if (exp_156) begin
          exp_157_reg <= exp_164;
        end
      end
      assign exp_157 = exp_157_reg;
    
  reg [31:0] exp_164_reg;
  always@(*) begin
    case (exp_159)
      0:exp_164_reg <= exp_161;
      1:exp_164_reg <= exp_162;
      default:exp_164_reg <= exp_163;
    endcase
  end
  assign exp_164 = exp_164_reg;
  assign exp_159 = exp_157 == exp_158;
  assign exp_158 = 4294967295;
  assign exp_163 = 0;
  assign exp_161 = exp_157 + exp_160;
  assign exp_160 = 1;
  assign exp_162 = 0;
  assign exp_156 = 1;

      reg [31:0] exp_167_reg = 0;
      always@(posedge clk) begin
        if (exp_166) begin
          exp_167_reg <= exp_174;
        end
      end
      assign exp_167 = exp_167_reg;
    
  reg [31:0] exp_174_reg;
  always@(*) begin
    case (exp_169)
      0:exp_174_reg <= exp_171;
      1:exp_174_reg <= exp_172;
      default:exp_174_reg <= exp_173;
    endcase
  end
  assign exp_174 = exp_174_reg;
  assign exp_169 = exp_167 == exp_168;
  assign exp_168 = 4294967295;
  assign exp_173 = 0;
  assign exp_171 = exp_167 + exp_170;
  assign exp_170 = 1;
  assign exp_172 = 0;
  assign exp_166 = exp_159 & exp_165;
  assign exp_165 = 1;
  assign exp_182 = exp_201;
  assign exp_201 = 0;
  assign exp_204 = exp_222;
  assign exp_222 = 0;
  assign exp_226 = exp_241;
  assign exp_241 = stdin_in;
  assign exp_461 = exp_248[15:8];
  assign exp_462 = exp_248[23:16];
  assign exp_463 = exp_248[31:24];
  assign exp_475 = $signed(exp_474);
  assign exp_474 = exp_473 + exp_469;
  assign exp_473 = 0;

  reg [15:0] exp_469_reg;
  always@(*) begin
    case (exp_459)
      0:exp_469_reg <= exp_466;
      1:exp_469_reg <= exp_467;
      default:exp_469_reg <= exp_468;
    endcase
  end
  assign exp_469 = exp_469_reg;
  assign exp_468 = 0;
  assign exp_466 = exp_248[15:0];
  assign exp_467 = exp_248[31:16];
  assign exp_476 = 0;
  assign exp_477 = exp_465;
  assign exp_478 = exp_469;
  assign exp_479 = 0;
  assign exp_480 = 0;

  reg [31:0] exp_839_reg;
  always@(*) begin
    case (exp_629)
      0:exp_839_reg <= exp_835;
      1:exp_839_reg <= exp_837;
      default:exp_839_reg <= exp_838;
    endcase
  end
  assign exp_839 = exp_839_reg;
  assign exp_838 = 0;

  reg [31:0] exp_835_reg;
  always@(*) begin
    case (exp_606)
      0:exp_835_reg <= exp_830;
      1:exp_835_reg <= exp_831;
      default:exp_835_reg <= exp_834;
    endcase
  end
  assign exp_835 = exp_835_reg;
  assign exp_606 = exp_605 & exp_603;
  assign exp_605 = exp_598 == exp_604;
  assign exp_604 = 0;
  assign exp_834 = 0;
  assign exp_830 = exp_829[63:32];

  reg [63:0] exp_829_reg;
  always@(*) begin
    case (exp_826)
      0:exp_829_reg <= exp_825;
      1:exp_829_reg <= exp_827;
      default:exp_829_reg <= exp_828;
    endcase
  end
  assign exp_829 = exp_829_reg;

      reg [0:0] exp_826_reg = 0;
      always@(posedge clk) begin
        if (exp_811) begin
          exp_826_reg <= exp_809;
        end
      end
      assign exp_826 = exp_826_reg;
    
      reg [0:0] exp_809_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_809_reg <= exp_786;
        end
      end
      assign exp_809 = exp_809_reg;
    
      reg [0:0] exp_786_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_786_reg <= exp_783;
        end
      end
      assign exp_786 = exp_786_reg;
      assign exp_783 = exp_781 ^ exp_782;
  assign exp_781 = exp_763 & exp_746;
  assign exp_763 = exp_762 + exp_761;
  assign exp_762 = 0;
  assign exp_761 = exp_759[31:31];

      reg [31:0] exp_759_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_759_reg <= exp_376;
        end
      end
      assign exp_759 = exp_759_reg;
      assign exp_758 = exp_748 == exp_757;
  assign exp_757 = 0;
  assign exp_746 = exp_745 | exp_612;
  assign exp_745 = exp_606 | exp_609;
  assign exp_609 = exp_608 & exp_603;
  assign exp_608 = exp_598 == exp_607;
  assign exp_607 = 1;
  assign exp_612 = exp_611 & exp_603;
  assign exp_611 = exp_598 == exp_610;
  assign exp_610 = 2;
  assign exp_782 = exp_766 & exp_747;
  assign exp_766 = exp_765 + exp_764;
  assign exp_765 = 0;
  assign exp_764 = exp_760[31:31];

      reg [31:0] exp_760_reg = 0;
      always@(posedge clk) begin
        if (exp_758) begin
          exp_760_reg <= exp_377;
        end
      end
      assign exp_760 = exp_760_reg;
      assign exp_747 = exp_606 | exp_609;
  assign exp_768 = exp_748 == exp_767;
  assign exp_767 = 1;
  assign exp_788 = exp_748 == exp_787;
  assign exp_787 = 2;
  assign exp_811 = exp_748 == exp_810;
  assign exp_810 = 3;
  assign exp_828 = 0;

      reg [63:0] exp_825_reg = 0;
      always@(posedge clk) begin
        if (exp_811) begin
          exp_825_reg <= exp_824;
        end
      end
      assign exp_825 = exp_825_reg;
      assign exp_824 = exp_820 + exp_823;
  assign exp_820 = exp_816 + exp_819;
  assign exp_816 = exp_812 + exp_815;
  assign exp_812 = exp_805;

      reg [31:0] exp_805_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_805_reg <= exp_792;
        end
      end
      assign exp_805 = exp_805_reg;
      assign exp_792 = exp_790 * exp_791;
  assign exp_790 = exp_789;
  assign exp_789 = exp_784[15:0];

      reg [31:0] exp_784_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_784_reg <= exp_774;
        end
      end
      assign exp_784 = exp_784_reg;
      assign exp_774 = exp_773 + exp_772;
  assign exp_773 = 0;

  reg [31:0] exp_772_reg;
  always@(*) begin
    case (exp_769)
      0:exp_772_reg <= exp_759;
      1:exp_772_reg <= exp_770;
      default:exp_772_reg <= exp_771;
    endcase
  end
  assign exp_772 = exp_772_reg;
  assign exp_769 = exp_763 & exp_746;
  assign exp_771 = 0;
  assign exp_770 = -exp_759;
  assign exp_791 = exp_785[15:0];

      reg [31:0] exp_785_reg = 0;
      always@(posedge clk) begin
        if (exp_768) begin
          exp_785_reg <= exp_780;
        end
      end
      assign exp_785 = exp_785_reg;
      assign exp_780 = exp_779 + exp_778;
  assign exp_779 = 0;

  reg [31:0] exp_778_reg;
  always@(*) begin
    case (exp_775)
      0:exp_778_reg <= exp_760;
      1:exp_778_reg <= exp_776;
      default:exp_778_reg <= exp_777;
    endcase
  end
  assign exp_778 = exp_778_reg;
  assign exp_775 = exp_766 & exp_747;
  assign exp_777 = 0;
  assign exp_776 = -exp_760;
  assign exp_815 = exp_813 << exp_814;
  assign exp_813 = exp_806;

      reg [31:0] exp_806_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_806_reg <= exp_796;
        end
      end
      assign exp_806 = exp_806_reg;
      assign exp_796 = exp_794 * exp_795;
  assign exp_794 = exp_793;
  assign exp_793 = exp_784[15:0];
  assign exp_795 = exp_785[31:16];
  assign exp_814 = 16;
  assign exp_819 = exp_817 << exp_818;
  assign exp_817 = exp_807;

      reg [31:0] exp_807_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_807_reg <= exp_800;
        end
      end
      assign exp_807 = exp_807_reg;
      assign exp_800 = exp_798 * exp_799;
  assign exp_798 = exp_797;
  assign exp_797 = exp_784[31:16];
  assign exp_799 = exp_785[15:0];
  assign exp_818 = 16;
  assign exp_823 = exp_821 << exp_822;
  assign exp_821 = exp_808;

      reg [31:0] exp_808_reg = 0;
      always@(posedge clk) begin
        if (exp_788) begin
          exp_808_reg <= exp_804;
        end
      end
      assign exp_808 = exp_808_reg;
      assign exp_804 = exp_802 * exp_803;
  assign exp_802 = exp_801;
  assign exp_801 = exp_784[31:16];
  assign exp_803 = exp_785[31:16];
  assign exp_822 = 32;
  assign exp_827 = -exp_825;
  assign exp_831 = exp_829[31:0];

  reg [31:0] exp_837_reg;
  always@(*) begin
    case (exp_630)
      0:exp_837_reg <= exp_740;
      1:exp_837_reg <= exp_741;
      default:exp_837_reg <= exp_836;
    endcase
  end
  assign exp_837 = exp_837_reg;
  assign exp_630 = exp_598[1:1];
  assign exp_836 = 0;

      reg [31:0] exp_740_reg = 0;
      always@(posedge clk) begin
        if (exp_649) begin
          exp_740_reg <= exp_734;
        end
      end
      assign exp_740 = exp_740_reg;
    
  reg [31:0] exp_734_reg;
  always@(*) begin
    case (exp_730)
      0:exp_734_reg <= exp_721;
      1:exp_734_reg <= exp_732;
      default:exp_734_reg <= exp_733;
    endcase
  end
  assign exp_734 = exp_734_reg;
  assign exp_730 = exp_729 & exp_632;
  assign exp_729 = exp_678 == exp_728;

      reg [31:0] exp_678_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_678_reg <= exp_675;
        end
      end
      assign exp_678 = exp_678_reg;
      assign exp_675 = exp_674 + exp_673;
  assign exp_674 = 0;

  reg [31:0] exp_673_reg;
  always@(*) begin
    case (exp_670)
      0:exp_673_reg <= exp_655;
      1:exp_673_reg <= exp_671;
      default:exp_673_reg <= exp_672;
    endcase
  end
  assign exp_673 = exp_673_reg;
  assign exp_670 = exp_661 & exp_632;
  assign exp_661 = exp_660 + exp_659;
  assign exp_660 = 0;
  assign exp_659 = exp_655[31:31];

      reg [31:0] exp_655_reg = 0;
      always@(posedge clk) begin
        if (exp_653) begin
          exp_655_reg <= exp_377;
        end
      end
      assign exp_655 = exp_655_reg;
      assign exp_653 = exp_635 == exp_652;
  assign exp_652 = 0;
  assign exp_632 = ~exp_631;
  assign exp_631 = exp_598[0:0];
  assign exp_672 = 0;
  assign exp_671 = -exp_655;
  assign exp_663 = exp_635 == exp_662;
  assign exp_662 = 1;
  assign exp_728 = 0;
  assign exp_733 = 0;
  assign exp_721 = exp_720 + exp_719;
  assign exp_720 = 0;

  reg [31:0] exp_719_reg;
  always@(*) begin
    case (exp_716)
      0:exp_719_reg <= exp_714;
      1:exp_719_reg <= exp_717;
      default:exp_719_reg <= exp_718;
    endcase
  end
  assign exp_719 = exp_719_reg;
  assign exp_716 = exp_680 & exp_632;

      reg [0:0] exp_680_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_680_reg <= exp_676;
        end
      end
      assign exp_680 = exp_680_reg;
      assign exp_676 = exp_658 ^ exp_661;
  assign exp_658 = exp_657 + exp_656;
  assign exp_657 = 0;
  assign exp_656 = exp_654[31:31];

      reg [31:0] exp_654_reg = 0;
      always@(posedge clk) begin
        if (exp_653) begin
          exp_654_reg <= exp_376;
        end
      end
      assign exp_654 = exp_654_reg;
      assign exp_718 = 0;

      reg [31:0] exp_714_reg = 0;
      always@(posedge clk) begin
        if (exp_647) begin
          exp_714_reg <= exp_684;
        end
      end
      assign exp_714 = exp_714_reg;
    
      reg [31:0] exp_684_reg = 0;
      always@(posedge clk) begin
        if (exp_683) begin
          exp_684_reg <= exp_711;
        end
      end
      assign exp_684 = exp_684_reg;
    
  reg [31:0] exp_711_reg;
  always@(*) begin
    case (exp_645)
      0:exp_711_reg <= exp_703;
      1:exp_711_reg <= exp_709;
      default:exp_711_reg <= exp_710;
    endcase
  end
  assign exp_711 = exp_711_reg;
  assign exp_645 = exp_635 == exp_644;
  assign exp_644 = 2;
  assign exp_710 = 0;

  reg [31:0] exp_703_reg;
  always@(*) begin
    case (exp_693)
      0:exp_703_reg <= exp_697;
      1:exp_703_reg <= exp_701;
      default:exp_703_reg <= exp_702;
    endcase
  end
  assign exp_703 = exp_703_reg;
  assign exp_693 = ~exp_692;
  assign exp_692 = exp_691[32:32];
  assign exp_691 = exp_690 - exp_678;
  assign exp_690 = exp_689;
  assign exp_689 = {exp_687, exp_688};  assign exp_687 = exp_682[31:0];

      reg [31:0] exp_682_reg = 0;
      always@(posedge clk) begin
        if (exp_681) begin
          exp_682_reg <= exp_708;
        end
      end
      assign exp_682 = exp_682_reg;
    
  reg [32:0] exp_708_reg;
  always@(*) begin
    case (exp_645)
      0:exp_708_reg <= exp_695;
      1:exp_708_reg <= exp_706;
      default:exp_708_reg <= exp_707;
    endcase
  end
  assign exp_708 = exp_708_reg;
  assign exp_707 = 0;

  reg [32:0] exp_695_reg;
  always@(*) begin
    case (exp_693)
      0:exp_695_reg <= exp_689;
      1:exp_695_reg <= exp_691;
      default:exp_695_reg <= exp_694;
    endcase
  end
  assign exp_695 = exp_695_reg;
  assign exp_694 = 0;
  assign exp_706 = 0;
  assign exp_681 = 1;
  assign exp_688 = exp_686[31:31];

      reg [31:0] exp_686_reg = 0;
      always@(posedge clk) begin
        if (exp_685) begin
          exp_686_reg <= exp_713;
        end
      end
      assign exp_686 = exp_686_reg;
    
  reg [31:0] exp_713_reg;
  always@(*) begin
    case (exp_645)
      0:exp_713_reg <= exp_705;
      1:exp_713_reg <= exp_677;
      default:exp_713_reg <= exp_712;
    endcase
  end
  assign exp_713 = exp_713_reg;
  assign exp_712 = 0;
  assign exp_705 = exp_686 << exp_704;
  assign exp_704 = 1;

      reg [31:0] exp_677_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_677_reg <= exp_669;
        end
      end
      assign exp_677 = exp_677_reg;
      assign exp_669 = exp_668 + exp_667;
  assign exp_668 = 0;

  reg [31:0] exp_667_reg;
  always@(*) begin
    case (exp_664)
      0:exp_667_reg <= exp_654;
      1:exp_667_reg <= exp_665;
      default:exp_667_reg <= exp_666;
    endcase
  end
  assign exp_667 = exp_667_reg;
  assign exp_664 = exp_658 & exp_632;
  assign exp_666 = 0;
  assign exp_665 = -exp_654;
  assign exp_685 = 1;
  assign exp_702 = 0;
  assign exp_697 = exp_684 << exp_696;
  assign exp_696 = 1;
  assign exp_701 = exp_699 | exp_700;
  assign exp_699 = exp_684 << exp_698;
  assign exp_698 = 1;
  assign exp_700 = 1;
  assign exp_709 = 0;
  assign exp_683 = 1;
  assign exp_647 = exp_635 == exp_646;
  assign exp_646 = 35;
  assign exp_717 = -exp_714;
  assign exp_732 = $signed(exp_731);
  assign exp_731 = -1;
  assign exp_649 = exp_635 == exp_648;
  assign exp_648 = 36;

      reg [31:0] exp_741_reg = 0;
      always@(posedge clk) begin
        if (exp_649) begin
          exp_741_reg <= exp_739;
        end
      end
      assign exp_741 = exp_741_reg;
    
  reg [31:0] exp_739_reg;
  always@(*) begin
    case (exp_737)
      0:exp_739_reg <= exp_727;
      1:exp_739_reg <= exp_654;
      default:exp_739_reg <= exp_738;
    endcase
  end
  assign exp_739 = exp_739_reg;
  assign exp_737 = exp_736 & exp_632;
  assign exp_736 = exp_678 == exp_735;
  assign exp_735 = 0;
  assign exp_738 = 0;
  assign exp_727 = exp_726 + exp_725;
  assign exp_726 = 0;

  reg [31:0] exp_725_reg;
  always@(*) begin
    case (exp_722)
      0:exp_725_reg <= exp_715;
      1:exp_725_reg <= exp_723;
      default:exp_725_reg <= exp_724;
    endcase
  end
  assign exp_725 = exp_725_reg;
  assign exp_722 = exp_679 & exp_632;

      reg [0:0] exp_679_reg = 0;
      always@(posedge clk) begin
        if (exp_663) begin
          exp_679_reg <= exp_658;
        end
      end
      assign exp_679 = exp_679_reg;
      assign exp_724 = 0;

      reg [31:0] exp_715_reg = 0;
      always@(posedge clk) begin
        if (exp_647) begin
          exp_715_reg <= exp_682;
        end
      end
      assign exp_715 = exp_715_reg;
      assign exp_723 = -exp_715;
  assign exp_310 = $signed(exp_309);
  assign exp_309 = 0;
  assign exp_539 = exp_374 != exp_375;
  assign exp_552 = 0;
  assign exp_553 = 0;
  assign exp_540 = $signed(exp_374) < $signed(exp_375);
  assign exp_541 = $signed(exp_374) >= $signed(exp_375);
  assign exp_546 = exp_543 < exp_545;
  assign exp_543 = exp_542 + exp_374;
  assign exp_542 = 0;
  assign exp_545 = exp_544 + exp_375;
  assign exp_544 = 0;
  assign exp_551 = exp_548 >= exp_550;
  assign exp_548 = exp_547 + exp_374;
  assign exp_547 = 0;
  assign exp_550 = exp_549 + exp_375;
  assign exp_549 = 0;
  assign exp_866 = 0;
  assign exp_865 = exp_264 + exp_864;
  assign exp_864 = 4;

  reg [32:0] exp_596_reg;
  always@(*) begin
    case (exp_397)
      0:exp_596_reg <= exp_586;
      1:exp_596_reg <= exp_594;
      default:exp_596_reg <= exp_595;
    endcase
  end
  assign exp_596 = exp_596_reg;
  assign exp_595 = 0;
  assign exp_586 = exp_585 + exp_383;

  reg [31:0] exp_585_reg;
  always@(*) begin
    case (exp_395)
      0:exp_585_reg <= exp_571;
      1:exp_585_reg <= exp_583;
      default:exp_585_reg <= exp_584;
    endcase
  end
  assign exp_585 = exp_585_reg;
  assign exp_584 = 0;
  assign exp_571 = $signed(exp_570);
  assign exp_570 = exp_569 + exp_568;
  assign exp_569 = 0;
  assign exp_568 = {exp_567, exp_564};  assign exp_567 = {exp_566, exp_563};  assign exp_566 = {exp_565, exp_562};  assign exp_565 = {exp_560, exp_561};  assign exp_560 = exp_382[31:31];
  assign exp_561 = exp_382[7:7];
  assign exp_562 = exp_382[30:25];
  assign exp_563 = exp_382[11:8];
  assign exp_564 = 0;
  assign exp_583 = $signed(exp_582);
  assign exp_582 = exp_581 + exp_580;
  assign exp_581 = 0;
  assign exp_580 = {exp_579, exp_576};  assign exp_579 = {exp_578, exp_575};  assign exp_578 = {exp_577, exp_574};  assign exp_577 = {exp_572, exp_573};  assign exp_572 = exp_382[31:31];
  assign exp_573 = exp_382[19:12];
  assign exp_574 = exp_382[20:20];
  assign exp_575 = exp_382[30:21];
  assign exp_576 = 0;

      reg [31:0] exp_383_reg = 0;
      always@(posedge clk) begin
        if (exp_373) begin
          exp_383_reg <= exp_266;
        end
      end
      assign exp_383 = exp_383_reg;
      assign exp_594 = exp_593 & exp_592;
  assign exp_593 = $signed(exp_591);
  assign exp_591 = exp_374 + exp_590;
  assign exp_590 = $signed(exp_589);
  assign exp_589 = exp_588 + exp_587;
  assign exp_588 = 0;
  assign exp_587 = exp_382[31:20];
  assign exp_592 = 4294967294;
  assign exp_263 = exp_256 & exp_254;
  assign exp_80 = exp_84;
  assign exp_76 = exp_83;
  assign exp_78 = exp_83;
  assign exp_9 = exp_265;
  assign exp_398 = 3;
  assign exp_244 = ~exp_229;
  assign exp_229 = exp_6;
  assign exp_200 = exp_184 & exp_185;
  assign exp_184 = exp_192;
  assign exp_192 = exp_5 & exp_191;
  assign exp_185 = exp_6;
  assign exp_181 = exp_2;

      reg [31:0] exp_221_reg = 0;
      always@(posedge clk) begin
        if (exp_220) begin
          exp_221_reg <= exp_203;
        end
      end
      assign exp_221 = exp_221_reg;
      assign exp_203 = exp_2;
  assign exp_220 = exp_206 & exp_207;
  assign exp_206 = exp_214;
  assign exp_214 = exp_5 & exp_213;
  assign exp_207 = exp_6;
  assign stdin_ready_out = exp_245;
  assign stdout_valid_out = exp_200;
  assign stdout_out = exp_181;
  assign leds_out = exp_221;

endmodule