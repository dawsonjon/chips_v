
module soc(clk, stdin_rx, stdout_tx, leds_out, pwm_pwm_out);
  input [0:0] stdin_rx;
  input [0:0] clk;
  output [0:0] stdout_tx;
  output [31:0] leds_out;
  output [0:0] pwm_pwm_out;
  wire [0:0] exp_333;
  wire [0:0] exp_429;
  wire [0:0] exp_427;
  wire [0:0] exp_426;
  wire [0:0] exp_416;
  wire [0:0] exp_370;
  wire [0:0] exp_415;
  wire [2:0] exp_325;
  wire [2:0] exp_447;
  wire [0:0] exp_445;
  wire [0:0] exp_444;
  wire [0:0] exp_443;
  wire [2:0] exp_442;
  wire [0:0] exp_365;
  wire [8:0] exp_335;
  wire [8:0] exp_454;
  wire [0:0] exp_452;
  wire [0:0] exp_451;
  wire [0:0] exp_453;
  wire [8:0] exp_440;
  wire [0:0] exp_438;
  wire [0:0] exp_437;
  wire [0:0] exp_351;
  wire [0:0] exp_350;
  wire [0:0] exp_439;
  wire [8:0] exp_425;
  wire [0:0] exp_423;
  wire [0:0] exp_424;
  wire [8:0] exp_412;
  wire [0:0] exp_410;
  wire [0:0] exp_393;
  wire [0:0] exp_392;
  wire [0:0] exp_391;
  wire [0:0] exp_409;
  wire [0:0] exp_341;
  wire [0:0] exp_340;
  wire [0:0] exp_411;
  wire [8:0] exp_399;
  wire [0:0] exp_397;
  wire [0:0] exp_398;
  wire [8:0] exp_383;
  wire [0:0] exp_381;
  wire [0:0] exp_374;
  wire [0:0] exp_373;
  wire [0:0] exp_372;
  wire [0:0] exp_323;
  wire [0:0] exp_309;
  wire [0:0] exp_315;
  wire [0:0] exp_11;
  wire [0:0] exp_534;
  wire [0:0] exp_531;
  wire [0:0] exp_525;
  wire [0:0] exp_882;
  wire [0:0] exp_819;
  wire [0:0] exp_684;
  wire [6:0] exp_669;
  wire [31:0] exp_667;
  wire [31:0] exp_104;
  wire [31:0] exp_103;
  wire [23:0] exp_102;
  wire [15:0] exp_101;
  wire [7:0] exp_90;
  wire [0:0] exp_89;
  wire [0:0] exp_94;
  wire [12:0] exp_85;
  wire [29:0] exp_93;
  wire [31:0] exp_16;
  wire [31:0] exp_549;
  wire [32:0] exp_1152;
  wire [0:0] exp_1148;
  wire [0:0] exp_844;
  wire [0:0] exp_822;
  wire [0:0] exp_680;
  wire [6:0] exp_679;
  wire [0:0] exp_682;
  wire [6:0] exp_681;
  wire [0:0] exp_843;
  wire [0:0] exp_688;
  wire [6:0] exp_687;
  wire [0:0] exp_842;
  wire [0:0] exp_841;
  wire [0:0] exp_840;
  wire [2:0] exp_670;
  wire [0:0] exp_839;
  wire [0:0] exp_823;
  wire [31:0] exp_659;
  wire [31:0] exp_597;
  wire [0:0] exp_593;
  wire [4:0] exp_573;
  wire [0:0] exp_592;
  wire [0:0] exp_596;
  wire [31:0] exp_589;
  wire [0:0] exp_570;
  wire [0:0] exp_1143;
  wire [0:0] exp_1142;
  wire [0:0] exp_1141;
  wire [0:0] exp_1140;
  wire [4:0] exp_552;
  wire [4:0] exp_1135;
  wire [0:0] exp_1134;
  wire [0:0] exp_726;
  wire [0:0] exp_725;
  wire [0:0] exp_724;
  wire [0:0] exp_723;
  wire [0:0] exp_722;
  wire [0:0] exp_721;
  wire [0:0] exp_672;
  wire [4:0] exp_671;
  wire [0:0] exp_674;
  wire [5:0] exp_673;
  wire [0:0] exp_676;
  wire [5:0] exp_675;
  wire [0:0] exp_678;
  wire [4:0] exp_677;
  wire [0:0] exp_1129;
  wire [0:0] exp_1128;
  wire [0:0] exp_914;
  wire [0:0] exp_888;
  wire [0:0] exp_886;
  wire [6:0] exp_884;
  wire [5:0] exp_885;
  wire [0:0] exp_887;
  wire [0:0] exp_913;
  wire [2:0] exp_883;
  wire [0:0] exp_1127;
  wire [0:0] exp_1125;
  wire [0:0] exp_1118;
  wire [2:0] exp_1033;
  wire [2:0] exp_1040;
  wire [0:0] exp_1035;
  wire [2:0] exp_1034;
  wire [0:0] exp_1039;
  wire [2:0] exp_1037;
  wire [0:0] exp_1036;
  wire [0:0] exp_1038;
  wire [0:0] exp_1029;
  wire [0:0] exp_1028;
  wire [0:0] exp_1027;
  wire [2:0] exp_1117;
  wire [0:0] exp_1126;
  wire [0:0] exp_936;
  wire [5:0] exp_920;
  wire [5:0] exp_927;
  wire [0:0] exp_922;
  wire [5:0] exp_921;
  wire [0:0] exp_926;
  wire [5:0] exp_924;
  wire [0:0] exp_923;
  wire [0:0] exp_925;
  wire [5:0] exp_935;
  wire [0:0] exp_547;
  wire [0:0] exp_546;
  wire [0:0] exp_544;
  wire [0:0] exp_543;
  wire [0:0] exp_541;
  wire [0:0] exp_542;
  wire [0:0] exp_540;
  wire [0:0] exp_1153;
  wire [0:0] exp_539;
  wire [0:0] exp_538;
  wire [0:0] exp_1157;
  wire [0:0] exp_1156;
  wire [0:0] exp_1155;
  wire [0:0] exp_1154;
  wire [0:0] exp_524;
  wire [0:0] exp_528;
  wire [0:0] exp_537;
  wire [0:0] exp_494;
  wire [0:0] exp_473;
  wire [0:0] exp_321;
  wire [0:0] exp_204;
  wire [0:0] exp_163;
  wire [0:0] exp_34;
  wire [0:0] exp_15;
  wire [0:0] exp_33;
  wire [0:0] exp_27;
  wire [7:0] exp_25;
  wire [31:0] exp_9;
  wire [31:0] exp_532;
  wire [31:0] exp_521;
  wire [31:0] exp_738;
  wire [31:0] exp_737;
  wire [31:0] exp_736;
  wire [31:0] exp_735;
  wire [11:0] exp_734;
  wire [11:0] exp_733;
  wire [11:0] exp_732;
  wire [0:0] exp_686;
  wire [5:0] exp_685;
  wire [0:0] exp_731;
  wire [11:0] exp_727;
  wire [11:0] exp_730;
  wire [6:0] exp_728;
  wire [4:0] exp_729;
  wire [0:0] exp_529;
  wire [0:0] exp_26;
  wire [0:0] exp_21;
  wire [0:0] exp_146;
  wire [0:0] exp_23;
  wire [0:0] exp_12;
  wire [0:0] exp_535;
  wire [0:0] exp_526;
  wire [0:0] exp_821;
  wire [0:0] exp_820;
  wire [0:0] exp_145;
  wire [0:0] exp_140;
  wire [0:0] exp_144;
  wire [0:0] exp_142;
  wire [0:0] exp_22;
  wire [0:0] exp_28;
  wire [0:0] exp_141;
  wire [0:0] exp_143;
  wire [0:0] exp_139;
  wire [0:0] exp_125;
  wire [0:0] exp_162;
  wire [0:0] exp_156;
  wire [7:0] exp_154;
  wire [0:0] exp_155;
  wire [0:0] exp_150;
  wire [0:0] exp_184;
  wire [0:0] exp_203;
  wire [0:0] exp_197;
  wire [7:0] exp_195;
  wire [1:0] exp_196;
  wire [0:0] exp_191;
  wire [0:0] exp_220;
  wire [0:0] exp_302;
  wire [0:0] exp_300;
  wire [0:0] exp_296;
  wire [0:0] exp_244;
  wire [0:0] exp_295;
  wire [2:0] exp_214;
  wire [2:0] exp_299;
  wire [0:0] exp_297;
  wire [0:0] exp_206;
  wire [0:0] exp_192;
  wire [0:0] exp_198;
  wire [0:0] exp_205;
  wire [0:0] exp_193;
  wire [0:0] exp_298;
  wire [2:0] exp_289;
  wire [0:0] exp_287;
  wire [0:0] exp_286;
  wire [0:0] exp_285;
  wire [1:0] exp_284;
  wire [0:0] exp_212;
  wire [0:0] exp_210;
  wire [0:0] exp_208;
  wire [0:0] exp_7;
  wire [0:0] exp_207;
  wire [0:0] exp_209;
  wire [0:0] exp_211;
  wire [0:0] exp_288;
  wire [2:0] exp_274;
  wire [0:0] exp_272;
  wire [0:0] exp_268;
  wire [0:0] exp_261;
  wire [0:0] exp_260;
  wire [0:0] exp_259;
  wire [0:0] exp_228;
  wire [9:0] exp_222;
  wire [9:0] exp_282;
  wire [0:0] exp_280;
  wire [0:0] exp_279;
  wire [0:0] exp_281;
  wire [9:0] exp_271;
  wire [0:0] exp_269;
  wire [0:0] exp_233;
  wire [2:0] exp_216;
  wire [2:0] exp_278;
  wire [0:0] exp_276;
  wire [0:0] exp_275;
  wire [0:0] exp_277;
  wire [2:0] exp_257;
  wire [0:0] exp_255;
  wire [0:0] exp_248;
  wire [0:0] exp_247;
  wire [0:0] exp_246;
  wire [0:0] exp_223;
  wire [0:0] exp_256;
  wire [2:0] exp_226;
  wire [2:0] exp_237;
  wire [0:0] exp_236;
  wire [0:0] exp_215;
  wire [2:0] exp_232;
  wire [0:0] exp_270;
  wire [9:0] exp_267;
  wire [0:0] exp_265;
  wire [0:0] exp_266;
  wire [9:0] exp_254;
  wire [0:0] exp_252;
  wire [0:0] exp_253;
  wire [9:0] exp_225;
  wire [9:0] exp_231;
  wire [9:0] exp_234;
  wire [9:0] exp_239;
  wire [0:0] exp_238;
  wire [0:0] exp_221;
  wire [0:0] exp_227;
  wire [0:0] exp_273;
  wire [2:0] exp_251;
  wire [0:0] exp_249;
  wire [0:0] exp_250;
  wire [2:0] exp_224;
  wire [2:0] exp_235;
  wire [2:0] exp_240;
  wire [2:0] exp_242;
  wire [0:0] exp_213;
  wire [2:0] exp_294;
  wire [0:0] exp_301;
  wire [0:0] exp_292;
  wire [0:0] exp_290;
  wire [0:0] exp_291;
  wire [0:0] exp_241;
  wire [0:0] exp_243;
  wire [0:0] exp_219;
  wire [0:0] exp_320;
  wire [0:0] exp_314;
  wire [7:0] exp_312;
  wire [1:0] exp_313;
  wire [0:0] exp_308;
  wire [0:0] exp_331;
  wire [0:0] exp_450;
  wire [0:0] exp_448;
  wire [0:0] exp_449;
  wire [0:0] exp_386;
  wire [0:0] exp_384;
  wire [0:0] exp_385;
  wire [0:0] exp_338;
  wire [0:0] exp_367;
  wire [0:0] exp_330;
  wire [0:0] exp_472;
  wire [0:0] exp_466;
  wire [7:0] exp_464;
  wire [2:0] exp_465;
  wire [0:0] exp_460;
  wire [0:0] exp_477;
  wire [0:0] exp_493;
  wire [0:0] exp_487;
  wire [7:0] exp_485;
  wire [2:0] exp_486;
  wire [0:0] exp_481;
  wire [0:0] exp_520;
  wire [0:0] exp_1131;
  wire [0:0] exp_1130;
  wire [0:0] exp_545;
  wire [0:0] exp_588;
  wire [31:0] exp_560;
  wire [0:0] exp_559;
  wire [1:0] exp_568;
  wire [4:0] exp_555;
  wire [0:0] exp_558;
  wire [0:0] exp_1137;
  wire [0:0] exp_1136;
  wire [4:0] exp_554;
  wire [31:0] exp_556;
  wire [31:0] exp_1133;
  wire [0:0] exp_1132;
  wire [31:0] exp_769;
  wire [0:0] exp_768;
  wire [31:0] exp_720;
  wire [2:0] exp_663;
  wire [2:0] exp_654;
  wire [0:0] exp_651;
  wire [0:0] exp_585;
  wire [6:0] exp_575;
  wire [6:0] exp_584;
  wire [0:0] exp_587;
  wire [6:0] exp_586;
  wire [0:0] exp_653;
  wire [2:0] exp_641;
  wire [0:0] exp_583;
  wire [4:0] exp_582;
  wire [0:0] exp_640;
  wire [2:0] exp_628;
  wire [0:0] exp_581;
  wire [5:0] exp_580;
  wire [0:0] exp_627;
  wire [2:0] exp_577;
  wire [0:0] exp_626;
  wire [0:0] exp_639;
  wire [0:0] exp_652;
  wire [0:0] exp_658;
  wire [0:0] exp_719;
  wire [31:0] exp_699;
  wire [0:0] exp_665;
  wire [0:0] exp_657;
  wire [0:0] exp_643;
  wire [0:0] exp_630;
  wire [0:0] exp_616;
  wire [0:0] exp_614;
  wire [0:0] exp_615;
  wire [0:0] exp_579;
  wire [4:0] exp_578;
  wire [0:0] exp_629;
  wire [0:0] exp_642;
  wire [0:0] exp_656;
  wire [0:0] exp_655;
  wire [0:0] exp_698;
  wire [31:0] exp_696;
  wire [31:0] exp_661;
  wire [31:0] exp_647;
  wire [0:0] exp_644;
  wire [0:0] exp_646;
  wire [31:0] exp_636;
  wire [0:0] exp_635;
  wire [31:0] exp_622;
  wire [0:0] exp_621;
  wire [31:0] exp_620;
  wire [31:0] exp_618;
  wire [19:0] exp_617;
  wire [3:0] exp_619;
  wire [31:0] exp_634;
  wire [31:0] exp_632;
  wire [19:0] exp_631;
  wire [3:0] exp_633;
  wire [31:0] exp_645;
  wire [31:0] exp_662;
  wire [31:0] exp_650;
  wire [0:0] exp_648;
  wire [0:0] exp_649;
  wire [31:0] exp_638;
  wire [0:0] exp_637;
  wire [31:0] exp_625;
  wire [0:0] exp_624;
  wire [31:0] exp_609;
  wire [0:0] exp_608;
  wire [31:0] exp_603;
  wire [0:0] exp_599;
  wire [4:0] exp_574;
  wire [0:0] exp_598;
  wire [0:0] exp_602;
  wire [31:0] exp_591;
  wire [0:0] exp_571;
  wire [0:0] exp_1147;
  wire [0:0] exp_1146;
  wire [0:0] exp_1145;
  wire [0:0] exp_1144;
  wire [4:0] exp_553;
  wire [0:0] exp_590;
  wire [31:0] exp_567;
  wire [0:0] exp_566;
  wire [1:0] exp_569;
  wire [4:0] exp_562;
  wire [0:0] exp_565;
  wire [0:0] exp_1139;
  wire [0:0] exp_1138;
  wire [4:0] exp_561;
  wire [31:0] exp_563;
  wire [31:0] exp_572;
  wire [31:0] exp_601;
  wire [0:0] exp_600;
  wire [31:0] exp_607;
  wire [31:0] exp_604;
  wire [31:0] exp_606;
  wire [11:0] exp_605;
  wire [31:0] exp_623;
  wire [31:0] exp_551;
  wire [0:0] exp_550;
  wire [31:0] exp_697;
  wire [31:0] exp_701;
  wire [31:0] exp_700;
  wire [5:0] exp_695;
  wire [5:0] exp_694;
  wire [5:0] exp_693;
  wire [4:0] exp_664;
  wire [4:0] exp_613;
  wire [0:0] exp_612;
  wire [4:0] exp_611;
  wire [4:0] exp_576;
  wire [31:0] exp_717;
  wire [1:0] exp_703;
  wire [0:0] exp_702;
  wire [31:0] exp_718;
  wire [1:0] exp_709;
  wire [0:0] exp_708;
  wire [31:0] exp_705;
  wire [31:0] exp_704;
  wire [31:0] exp_707;
  wire [31:0] exp_706;
  wire [31:0] exp_710;
  wire [31:0] exp_714;
  wire [32:0] exp_713;
  wire [32:0] exp_711;
  wire [0:0] exp_692;
  wire [0:0] exp_666;
  wire [0:0] exp_610;
  wire [0:0] exp_691;
  wire [0:0] exp_690;
  wire [0:0] exp_689;
  wire [32:0] exp_712;
  wire [31:0] exp_715;
  wire [31:0] exp_716;
  wire [31:0] exp_767;
  wire [0:0] exp_766;
  wire [31:0] exp_757;
  wire [7:0] exp_756;
  wire [7:0] exp_755;
  wire [7:0] exp_750;
  wire [1:0] exp_741;
  wire [1:0] exp_740;
  wire [1:0] exp_739;
  wire [0:0] exp_749;
  wire [7:0] exp_745;
  wire [31:0] exp_523;
  wire [31:0] exp_492;
  wire [31:0] exp_471;
  wire [31:0] exp_319;
  wire [31:0] exp_202;
  wire [31:0] exp_161;
  wire [31:0] exp_32;
  wire [31:0] exp_14;
  wire [31:0] exp_31;
  wire [0:0] exp_30;
  wire [31:0] exp_29;
  wire [31:0] exp_20;
  wire [31:0] exp_127;
  wire [31:0] exp_138;
  wire [23:0] exp_137;
  wire [15:0] exp_136;
  wire [7:0] exp_62;
  wire [0:0] exp_61;
  wire [0:0] exp_129;
  wire [12:0] exp_57;
  wire [29:0] exp_128;
  wire [31:0] exp_18;
  wire [0:0] exp_60;
  wire [0:0] exp_124;
  wire [0:0] exp_122;
  wire [0:0] exp_123;
  wire [3:0] exp_24;
  wire [3:0] exp_13;
  wire [3:0] exp_536;
  wire [3:0] exp_527;
  wire [3:0] exp_818;
  wire [0:0] exp_817;
  wire [3:0] exp_805;
  wire [3:0] exp_801;
  wire [1:0] exp_804;
  wire [1:0] exp_803;
  wire [1:0] exp_802;
  wire [3:0] exp_810;
  wire [3:0] exp_806;
  wire [0:0] exp_809;
  wire [0:0] exp_808;
  wire [0:0] exp_807;
  wire [3:0] exp_811;
  wire [3:0] exp_812;
  wire [3:0] exp_813;
  wire [3:0] exp_814;
  wire [3:0] exp_815;
  wire [3:0] exp_816;
  wire [12:0] exp_56;
  wire [29:0] exp_120;
  wire [7:0] exp_58;
  wire [7:0] exp_121;
  wire [31:0] exp_19;
  wire [31:0] exp_10;
  wire [31:0] exp_533;
  wire [31:0] exp_522;
  wire [31:0] exp_800;
  wire [0:0] exp_799;
  wire [31:0] exp_787;
  wire [0:0] exp_786;
  wire [31:0] exp_773;
  wire [7:0] exp_772;
  wire [7:0] exp_771;
  wire [7:0] exp_770;
  wire [31:0] exp_660;
  wire [31:0] exp_781;
  wire [3:0] exp_780;
  wire [31:0] exp_783;
  wire [4:0] exp_782;
  wire [31:0] exp_785;
  wire [4:0] exp_784;
  wire [31:0] exp_791;
  wire [0:0] exp_744;
  wire [0:0] exp_743;
  wire [0:0] exp_742;
  wire [0:0] exp_790;
  wire [31:0] exp_777;
  wire [15:0] exp_776;
  wire [15:0] exp_775;
  wire [15:0] exp_774;
  wire [31:0] exp_789;
  wire [4:0] exp_788;
  wire [31:0] exp_793;
  wire [31:0] exp_792;
  wire [31:0] exp_779;
  wire [31:0] exp_778;
  wire [31:0] exp_794;
  wire [31:0] exp_795;
  wire [31:0] exp_796;
  wire [31:0] exp_797;
  wire [31:0] exp_798;
  wire [7:0] exp_55;
  wire [7:0] exp_83;
  wire [0:0] exp_82;
  wire [0:0] exp_96;
  wire [12:0] exp_78;
  wire [29:0] exp_95;
  wire [0:0] exp_81;
  wire [0:0] exp_92;
  wire [12:0] exp_77;
  wire [31:0] exp_91;
  wire [7:0] exp_79;
  wire [0:0] exp_54;
  wire [0:0] exp_131;
  wire [12:0] exp_50;
  wire [29:0] exp_130;
  wire [0:0] exp_53;
  wire [0:0] exp_119;
  wire [0:0] exp_117;
  wire [0:0] exp_118;
  wire [12:0] exp_49;
  wire [29:0] exp_115;
  wire [7:0] exp_51;
  wire [7:0] exp_116;
  wire [7:0] exp_48;
  wire [7:0] exp_76;
  wire [0:0] exp_75;
  wire [0:0] exp_98;
  wire [12:0] exp_71;
  wire [29:0] exp_97;
  wire [0:0] exp_74;
  wire [12:0] exp_70;
  wire [7:0] exp_72;
  wire [0:0] exp_47;
  wire [0:0] exp_133;
  wire [12:0] exp_43;
  wire [29:0] exp_132;
  wire [0:0] exp_46;
  wire [0:0] exp_114;
  wire [0:0] exp_112;
  wire [0:0] exp_113;
  wire [12:0] exp_42;
  wire [29:0] exp_110;
  wire [7:0] exp_44;
  wire [7:0] exp_111;
  wire [7:0] exp_41;
  wire [7:0] exp_69;
  wire [0:0] exp_68;
  wire [0:0] exp_100;
  wire [12:0] exp_64;
  wire [29:0] exp_99;
  wire [0:0] exp_67;
  wire [12:0] exp_63;
  wire [7:0] exp_65;
  wire [0:0] exp_40;
  wire [0:0] exp_135;
  wire [12:0] exp_36;
  wire [29:0] exp_134;
  wire [0:0] exp_39;
  wire [0:0] exp_109;
  wire [0:0] exp_107;
  wire [0:0] exp_108;
  wire [12:0] exp_35;
  wire [29:0] exp_105;
  wire [7:0] exp_37;
  wire [7:0] exp_106;
  wire [0:0] exp_126;
  wire [31:0] exp_160;
  wire [0:0] exp_159;
  wire [31:0] exp_158;
  wire [31:0] exp_149;
  wire [31:0] exp_187;
  wire [0:0] exp_185;
  wire [31:0] exp_147;
  wire [0:0] exp_186;
  wire [31:0] exp_165;
  wire [31:0] exp_172;
  wire [0:0] exp_167;
  wire [31:0] exp_166;
  wire [0:0] exp_171;
  wire [31:0] exp_169;
  wire [0:0] exp_168;
  wire [0:0] exp_170;
  wire [0:0] exp_164;
  wire [31:0] exp_175;
  wire [31:0] exp_182;
  wire [0:0] exp_177;
  wire [31:0] exp_176;
  wire [0:0] exp_181;
  wire [31:0] exp_179;
  wire [0:0] exp_178;
  wire [0:0] exp_180;
  wire [0:0] exp_174;
  wire [0:0] exp_173;
  wire [31:0] exp_201;
  wire [0:0] exp_200;
  wire [31:0] exp_199;
  wire [31:0] exp_190;
  wire [31:0] exp_304;
  wire [7:0] exp_218;
  wire [7:0] exp_264;
  wire [0:0] exp_262;
  wire [0:0] exp_263;
  wire [7:0] exp_230;
  wire [6:0] exp_229;
  wire [0:0] exp_217;
  wire [31:0] exp_318;
  wire [0:0] exp_317;
  wire [31:0] exp_316;
  wire [31:0] exp_307;
  wire [31:0] exp_456;
  wire [31:0] exp_470;
  wire [0:0] exp_469;
  wire [31:0] exp_468;
  wire [31:0] exp_459;
  wire [31:0] exp_476;
  wire [31:0] exp_491;
  wire [0:0] exp_490;
  wire [31:0] exp_489;
  wire [31:0] exp_480;
  wire [31:0] exp_519;
  wire [7:0] exp_746;
  wire [7:0] exp_747;
  wire [7:0] exp_748;
  wire [31:0] exp_760;
  wire [15:0] exp_759;
  wire [15:0] exp_758;
  wire [15:0] exp_754;
  wire [0:0] exp_753;
  wire [15:0] exp_751;
  wire [15:0] exp_752;
  wire [31:0] exp_761;
  wire [31:0] exp_762;
  wire [31:0] exp_763;
  wire [31:0] exp_764;
  wire [31:0] exp_765;
  wire [31:0] exp_1124;
  wire [0:0] exp_1123;
  wire [31:0] exp_1120;
  wire [0:0] exp_891;
  wire [0:0] exp_890;
  wire [0:0] exp_889;
  wire [0:0] exp_1119;
  wire [31:0] exp_1115;
  wire [63:0] exp_1114;
  wire [0:0] exp_1111;
  wire [0:0] exp_1094;
  wire [0:0] exp_1071;
  wire [0:0] exp_1068;
  wire [0:0] exp_1066;
  wire [0:0] exp_1048;
  wire [0:0] exp_1047;
  wire [0:0] exp_1046;
  wire [31:0] exp_1044;
  wire [0:0] exp_1043;
  wire [0:0] exp_1042;
  wire [0:0] exp_1031;
  wire [0:0] exp_1030;
  wire [0:0] exp_894;
  wire [0:0] exp_893;
  wire [0:0] exp_892;
  wire [0:0] exp_897;
  wire [0:0] exp_896;
  wire [1:0] exp_895;
  wire [0:0] exp_1067;
  wire [0:0] exp_1051;
  wire [0:0] exp_1050;
  wire [0:0] exp_1049;
  wire [31:0] exp_1045;
  wire [0:0] exp_1032;
  wire [0:0] exp_1053;
  wire [0:0] exp_1052;
  wire [0:0] exp_1073;
  wire [1:0] exp_1072;
  wire [0:0] exp_1096;
  wire [1:0] exp_1095;
  wire [0:0] exp_1113;
  wire [63:0] exp_1110;
  wire [63:0] exp_1109;
  wire [63:0] exp_1105;
  wire [63:0] exp_1101;
  wire [63:0] exp_1097;
  wire [31:0] exp_1090;
  wire [31:0] exp_1077;
  wire [31:0] exp_1075;
  wire [15:0] exp_1074;
  wire [31:0] exp_1069;
  wire [31:0] exp_1059;
  wire [31:0] exp_1058;
  wire [31:0] exp_1057;
  wire [0:0] exp_1054;
  wire [0:0] exp_1056;
  wire [31:0] exp_1055;
  wire [15:0] exp_1076;
  wire [31:0] exp_1070;
  wire [31:0] exp_1065;
  wire [31:0] exp_1064;
  wire [31:0] exp_1063;
  wire [0:0] exp_1060;
  wire [0:0] exp_1062;
  wire [31:0] exp_1061;
  wire [63:0] exp_1100;
  wire [63:0] exp_1098;
  wire [31:0] exp_1091;
  wire [31:0] exp_1081;
  wire [31:0] exp_1079;
  wire [15:0] exp_1078;
  wire [15:0] exp_1080;
  wire [4:0] exp_1099;
  wire [63:0] exp_1104;
  wire [63:0] exp_1102;
  wire [31:0] exp_1092;
  wire [31:0] exp_1085;
  wire [31:0] exp_1083;
  wire [15:0] exp_1082;
  wire [15:0] exp_1084;
  wire [4:0] exp_1103;
  wire [63:0] exp_1108;
  wire [63:0] exp_1106;
  wire [31:0] exp_1093;
  wire [31:0] exp_1089;
  wire [31:0] exp_1087;
  wire [15:0] exp_1086;
  wire [15:0] exp_1088;
  wire [5:0] exp_1107;
  wire [63:0] exp_1112;
  wire [31:0] exp_1116;
  wire [31:0] exp_1122;
  wire [0:0] exp_915;
  wire [0:0] exp_1121;
  wire [31:0] exp_1025;
  wire [31:0] exp_1019;
  wire [0:0] exp_1015;
  wire [0:0] exp_1014;
  wire [31:0] exp_963;
  wire [31:0] exp_960;
  wire [31:0] exp_959;
  wire [31:0] exp_958;
  wire [0:0] exp_955;
  wire [0:0] exp_946;
  wire [0:0] exp_945;
  wire [0:0] exp_944;
  wire [31:0] exp_940;
  wire [0:0] exp_938;
  wire [0:0] exp_937;
  wire [0:0] exp_917;
  wire [0:0] exp_916;
  wire [0:0] exp_957;
  wire [31:0] exp_956;
  wire [0:0] exp_948;
  wire [0:0] exp_947;
  wire [0:0] exp_1013;
  wire [0:0] exp_1018;
  wire [31:0] exp_1006;
  wire [31:0] exp_1005;
  wire [31:0] exp_1004;
  wire [0:0] exp_1001;
  wire [0:0] exp_965;
  wire [0:0] exp_961;
  wire [0:0] exp_943;
  wire [0:0] exp_942;
  wire [0:0] exp_941;
  wire [31:0] exp_939;
  wire [0:0] exp_1003;
  wire [31:0] exp_999;
  wire [31:0] exp_969;
  wire [31:0] exp_996;
  wire [0:0] exp_930;
  wire [1:0] exp_929;
  wire [0:0] exp_995;
  wire [31:0] exp_988;
  wire [0:0] exp_978;
  wire [0:0] exp_977;
  wire [32:0] exp_976;
  wire [32:0] exp_975;
  wire [32:0] exp_974;
  wire [31:0] exp_972;
  wire [31:0] exp_967;
  wire [32:0] exp_993;
  wire [0:0] exp_992;
  wire [32:0] exp_980;
  wire [0:0] exp_979;
  wire [0:0] exp_991;
  wire [0:0] exp_966;
  wire [0:0] exp_973;
  wire [31:0] exp_971;
  wire [31:0] exp_998;
  wire [0:0] exp_997;
  wire [31:0] exp_990;
  wire [0:0] exp_989;
  wire [31:0] exp_962;
  wire [31:0] exp_954;
  wire [31:0] exp_953;
  wire [31:0] exp_952;
  wire [0:0] exp_949;
  wire [0:0] exp_951;
  wire [31:0] exp_950;
  wire [0:0] exp_970;
  wire [0:0] exp_987;
  wire [31:0] exp_982;
  wire [0:0] exp_981;
  wire [31:0] exp_986;
  wire [31:0] exp_984;
  wire [0:0] exp_983;
  wire [0:0] exp_985;
  wire [0:0] exp_994;
  wire [0:0] exp_968;
  wire [0:0] exp_932;
  wire [5:0] exp_931;
  wire [31:0] exp_1002;
  wire [31:0] exp_1017;
  wire [0:0] exp_1016;
  wire [0:0] exp_934;
  wire [5:0] exp_933;
  wire [31:0] exp_1026;
  wire [31:0] exp_1024;
  wire [0:0] exp_1022;
  wire [0:0] exp_1021;
  wire [0:0] exp_1020;
  wire [0:0] exp_1023;
  wire [31:0] exp_1012;
  wire [31:0] exp_1011;
  wire [31:0] exp_1010;
  wire [0:0] exp_1007;
  wire [0:0] exp_964;
  wire [0:0] exp_1009;
  wire [31:0] exp_1000;
  wire [31:0] exp_1008;
  wire [31:0] exp_595;
  wire [0:0] exp_594;
  wire [0:0] exp_824;
  wire [0:0] exp_837;
  wire [0:0] exp_838;
  wire [0:0] exp_825;
  wire [0:0] exp_826;
  wire [0:0] exp_831;
  wire [31:0] exp_828;
  wire [31:0] exp_827;
  wire [31:0] exp_830;
  wire [31:0] exp_829;
  wire [0:0] exp_836;
  wire [31:0] exp_833;
  wire [31:0] exp_832;
  wire [31:0] exp_835;
  wire [31:0] exp_834;
  wire [0:0] exp_1151;
  wire [31:0] exp_1150;
  wire [2:0] exp_1149;
  wire [32:0] exp_881;
  wire [0:0] exp_880;
  wire [31:0] exp_871;
  wire [31:0] exp_870;
  wire [0:0] exp_869;
  wire [31:0] exp_856;
  wire [12:0] exp_855;
  wire [12:0] exp_854;
  wire [12:0] exp_853;
  wire [11:0] exp_852;
  wire [7:0] exp_851;
  wire [1:0] exp_850;
  wire [0:0] exp_845;
  wire [0:0] exp_846;
  wire [5:0] exp_847;
  wire [3:0] exp_848;
  wire [0:0] exp_849;
  wire [31:0] exp_868;
  wire [20:0] exp_867;
  wire [20:0] exp_866;
  wire [20:0] exp_865;
  wire [19:0] exp_864;
  wire [9:0] exp_863;
  wire [8:0] exp_862;
  wire [0:0] exp_857;
  wire [7:0] exp_858;
  wire [0:0] exp_859;
  wire [9:0] exp_860;
  wire [0:0] exp_861;
  wire [31:0] exp_668;
  wire [32:0] exp_879;
  wire [32:0] exp_878;
  wire [31:0] exp_876;
  wire [31:0] exp_875;
  wire [11:0] exp_874;
  wire [11:0] exp_873;
  wire [11:0] exp_872;
  wire [32:0] exp_877;
  wire [0:0] exp_548;
  wire [0:0] exp_88;
  wire [12:0] exp_84;
  wire [7:0] exp_86;
  wire [0:0] exp_17;
  wire [1:0] exp_683;
  wire [0:0] exp_530;
  wire [0:0] exp_310;
  wire [0:0] exp_382;
  wire [8:0] exp_337;
  wire [8:0] exp_343;
  wire [8:0] exp_349;
  wire [0:0] exp_348;
  wire [8:0] exp_355;
  wire [8:0] exp_363;
  wire [0:0] exp_362;
  wire [8:0] exp_369;
  wire [0:0] exp_368;
  wire [0:0] exp_334;
  wire [0:0] exp_364;
  wire [0:0] exp_446;
  wire [2:0] exp_432;
  wire [0:0] exp_430;
  wire [0:0] exp_357;
  wire [2:0] exp_327;
  wire [2:0] exp_436;
  wire [0:0] exp_434;
  wire [0:0] exp_433;
  wire [0:0] exp_435;
  wire [2:0] exp_402;
  wire [0:0] exp_400;
  wire [0:0] exp_401;
  wire [2:0] exp_344;
  wire [2:0] exp_361;
  wire [0:0] exp_360;
  wire [0:0] exp_326;
  wire [2:0] exp_356;
  wire [0:0] exp_431;
  wire [2:0] exp_396;
  wire [0:0] exp_394;
  wire [0:0] exp_395;
  wire [2:0] exp_380;
  wire [0:0] exp_378;
  wire [0:0] exp_379;
  wire [2:0] exp_336;
  wire [2:0] exp_342;
  wire [2:0] exp_359;
  wire [2:0] exp_366;
  wire [0:0] exp_324;
  wire [1:0] exp_414;
  wire [0:0] exp_428;
  wire [0:0] exp_422;
  wire [0:0] exp_420;
  wire [0:0] exp_421;
  wire [0:0] exp_405;
  wire [0:0] exp_403;
  wire [0:0] exp_404;
  wire [0:0] exp_389;
  wire [0:0] exp_387;
  wire [0:0] exp_388;
  wire [0:0] exp_339;
  wire [0:0] exp_345;
  wire [7:0] exp_329;
  wire [7:0] exp_419;
  wire [0:0] exp_417;
  wire [0:0] exp_418;
  wire [7:0] exp_408;
  wire [0:0] exp_406;
  wire [0:0] exp_407;
  wire [7:0] exp_377;
  wire [0:0] exp_375;
  wire [0:0] exp_376;
  wire [7:0] exp_322;
  wire [31:0] exp_306;
  wire [7:0] exp_347;
  wire [0:0] exp_346;
  wire [7:0] exp_353;
  wire [0:0] exp_352;
  wire [0:0] exp_328;
  wire [0:0] exp_354;
  wire [0:0] exp_358;
  wire [0:0] exp_332;
  wire [31:0] exp_475;
  wire [31:0] exp_458;
  wire [0:0] exp_474;
  wire [0:0] exp_461;
  wire [0:0] exp_467;
  wire [0:0] exp_462;
  wire [0:0] exp_518;
  wire [10:0] exp_517;
  wire [31:0] exp_479;
  wire [0:0] exp_495;
  wire [0:0] exp_482;
  wire [0:0] exp_488;
  wire [0:0] exp_483;
  wire [9:0] exp_507;
  wire [9:0] exp_514;
  wire [0:0] exp_509;
  wire [9:0] exp_508;
  wire [0:0] exp_513;
  wire [9:0] exp_511;
  wire [0:0] exp_510;
  wire [0:0] exp_512;
  wire [0:0] exp_506;
  wire [0:0] exp_499;
  wire [1:0] exp_497;
  wire [1:0] exp_504;
  wire [0:0] exp_503;
  wire [1:0] exp_501;
  wire [0:0] exp_500;
  wire [0:0] exp_502;
  wire [0:0] exp_496;
  wire [1:0] exp_498;
  wire [0:0] exp_505;


      reg [0:0] exp_333_reg = 1;
      always@(posedge clk) begin
        if (exp_332) begin
          exp_333_reg <= exp_429;
        end
      end
      assign exp_333 = exp_333_reg;
    
  reg [0:0] exp_429_reg;
  always@(*) begin
    case (exp_427)
      0:exp_429_reg <= exp_422;
      1:exp_429_reg <= exp_358;
      default:exp_429_reg <= exp_428;
    endcase
  end
  assign exp_429 = exp_429_reg;
  assign exp_427 = exp_426 & exp_357;
  assign exp_426 = exp_416 & exp_351;
  assign exp_416 = exp_370 & exp_415;
  assign exp_370 = 1;
  assign exp_415 = exp_325 == exp_414;

      reg [2:0] exp_325_reg = 0;
      always@(posedge clk) begin
        if (exp_324) begin
          exp_325_reg <= exp_447;
        end
      end
      assign exp_325 = exp_325_reg;
    
  reg [2:0] exp_447_reg;
  always@(*) begin
    case (exp_445)
      0:exp_447_reg <= exp_432;
      1:exp_447_reg <= exp_366;
      default:exp_447_reg <= exp_446;
    endcase
  end
  assign exp_447 = exp_447_reg;
  assign exp_445 = exp_444 & exp_365;
  assign exp_444 = exp_370 & exp_443;
  assign exp_443 = exp_325 == exp_442;
  assign exp_442 = 4;
  assign exp_365 = exp_335 == exp_364;

      reg [8:0] exp_335_reg = 0;
      always@(posedge clk) begin
        if (exp_334) begin
          exp_335_reg <= exp_454;
        end
      end
      assign exp_335 = exp_335_reg;
    
  reg [8:0] exp_454_reg;
  always@(*) begin
    case (exp_452)
      0:exp_454_reg <= exp_440;
      1:exp_454_reg <= exp_369;
      default:exp_454_reg <= exp_453;
    endcase
  end
  assign exp_454 = exp_454_reg;
  assign exp_452 = exp_444 & exp_451;
  assign exp_451 = ~exp_365;
  assign exp_453 = 0;

  reg [8:0] exp_440_reg;
  always@(*) begin
    case (exp_438)
      0:exp_440_reg <= exp_425;
      1:exp_440_reg <= exp_363;
      default:exp_440_reg <= exp_439;
    endcase
  end
  assign exp_440 = exp_440_reg;
  assign exp_438 = exp_416 & exp_437;
  assign exp_437 = ~exp_351;
  assign exp_351 = exp_335 == exp_350;
  assign exp_350 = 0;
  assign exp_439 = 0;

  reg [8:0] exp_425_reg;
  always@(*) begin
    case (exp_423)
      0:exp_425_reg <= exp_412;
      1:exp_425_reg <= exp_355;
      default:exp_425_reg <= exp_424;
    endcase
  end
  assign exp_425 = exp_425_reg;
  assign exp_423 = exp_416 & exp_351;
  assign exp_424 = 0;

  reg [8:0] exp_412_reg;
  always@(*) begin
    case (exp_410)
      0:exp_412_reg <= exp_399;
      1:exp_412_reg <= exp_349;
      default:exp_412_reg <= exp_411;
    endcase
  end
  assign exp_412 = exp_412_reg;
  assign exp_410 = exp_393 & exp_409;
  assign exp_393 = exp_370 & exp_392;
  assign exp_392 = exp_325 == exp_391;
  assign exp_391 = 1;
  assign exp_409 = ~exp_341;
  assign exp_341 = exp_335 == exp_340;
  assign exp_340 = 0;
  assign exp_411 = 0;

  reg [8:0] exp_399_reg;
  always@(*) begin
    case (exp_397)
      0:exp_399_reg <= exp_383;
      1:exp_399_reg <= exp_343;
      default:exp_399_reg <= exp_398;
    endcase
  end
  assign exp_399 = exp_399_reg;
  assign exp_397 = exp_393 & exp_341;
  assign exp_398 = 0;

  reg [8:0] exp_383_reg;
  always@(*) begin
    case (exp_381)
      0:exp_383_reg <= exp_335;
      1:exp_383_reg <= exp_337;
      default:exp_383_reg <= exp_382;
    endcase
  end
  assign exp_383 = exp_383_reg;
  assign exp_381 = exp_374 & exp_323;
  assign exp_374 = exp_370 & exp_373;
  assign exp_373 = exp_325 == exp_372;
  assign exp_372 = 0;
  assign exp_323 = exp_309 & exp_310;
  assign exp_309 = exp_315;
  assign exp_315 = exp_11 & exp_314;
  assign exp_11 = exp_534;

      reg [0:0] exp_534_reg = 0;
      always@(posedge clk) begin
        if (exp_529) begin
          exp_534_reg <= exp_531;
        end
      end
      assign exp_534 = exp_534_reg;
      assign exp_531 = exp_525 & exp_530;
  assign exp_525 = exp_882;
  assign exp_882 = exp_819 & exp_547;
  assign exp_819 = exp_684 | exp_686;
  assign exp_684 = exp_669 == exp_683;
  assign exp_669 = exp_667[6:0];

      reg [31:0] exp_667_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_667_reg <= exp_104;
        end
      end
      assign exp_667 = exp_667_reg;
    
      reg [31:0] exp_104_reg = 0;
      always@(posedge clk) begin
        if (exp_17) begin
          exp_104_reg <= exp_103;
        end
      end
      assign exp_104 = exp_104_reg;
      assign exp_103 = {exp_102, exp_69};  assign exp_102 = {exp_101, exp_76};  assign exp_101 = {exp_90, exp_83};  assign exp_89 = exp_94;
  assign exp_94 = 1;
  assign exp_85 = exp_93;
  assign exp_93 = exp_16[31:2];
  assign exp_16 = exp_549;

      reg [31:0] exp_549_reg = 0;
      always@(posedge clk) begin
        if (exp_548) begin
          exp_549_reg <= exp_1152;
        end
      end
      assign exp_549 = exp_549_reg;
    
  reg [32:0] exp_1152_reg;
  always@(*) begin
    case (exp_1148)
      0:exp_1152_reg <= exp_1150;
      1:exp_1152_reg <= exp_881;
      default:exp_1152_reg <= exp_1151;
    endcase
  end
  assign exp_1152 = exp_1152_reg;
  assign exp_1148 = exp_844 & exp_547;
  assign exp_844 = exp_822 | exp_843;
  assign exp_822 = exp_680 | exp_682;
  assign exp_680 = exp_669 == exp_679;
  assign exp_679 = 111;
  assign exp_682 = exp_669 == exp_681;
  assign exp_681 = 103;

  reg [0:0] exp_843_reg;
  always@(*) begin
    case (exp_688)
      0:exp_843_reg <= exp_841;
      1:exp_843_reg <= exp_840;
      default:exp_843_reg <= exp_842;
    endcase
  end
  assign exp_843 = exp_843_reg;
  assign exp_688 = exp_669 == exp_687;
  assign exp_687 = 99;
  assign exp_842 = 0;
  assign exp_841 = 0;

  reg [0:0] exp_840_reg;
  always@(*) begin
    case (exp_670)
      0:exp_840_reg <= exp_823;
      1:exp_840_reg <= exp_824;
      2:exp_840_reg <= exp_837;
      3:exp_840_reg <= exp_838;
      4:exp_840_reg <= exp_825;
      5:exp_840_reg <= exp_826;
      6:exp_840_reg <= exp_831;
      7:exp_840_reg <= exp_836;
      default:exp_840_reg <= exp_839;
    endcase
  end
  assign exp_840 = exp_840_reg;
  assign exp_670 = exp_667[14:12];
  assign exp_839 = 0;
  assign exp_823 = exp_659 == exp_660;

      reg [31:0] exp_659_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_659_reg <= exp_597;
        end
      end
      assign exp_659 = exp_659_reg;
    
  reg [31:0] exp_597_reg;
  always@(*) begin
    case (exp_593)
      0:exp_597_reg <= exp_589;
      1:exp_597_reg <= exp_595;
      default:exp_597_reg <= exp_596;
    endcase
  end
  assign exp_597 = exp_597_reg;
  assign exp_593 = exp_573 == exp_592;
  assign exp_573 = exp_104[19:15];
  assign exp_592 = 0;
  assign exp_596 = 0;

  reg [31:0] exp_589_reg;
  always@(*) begin
    case (exp_570)
      0:exp_589_reg <= exp_560;
      1:exp_589_reg <= exp_572;
      default:exp_589_reg <= exp_588;
    endcase
  end
  assign exp_589 = exp_589_reg;
  assign exp_570 = exp_1143;
  assign exp_1143 = exp_1142 & exp_539;
  assign exp_1142 = exp_1141 & exp_547;
  assign exp_1141 = exp_1140 & exp_1134;
  assign exp_1140 = exp_552 == exp_1135;
  assign exp_552 = exp_104[19:15];
  assign exp_1135 = exp_667[11:7];
  assign exp_1134 = exp_726 | exp_1129;
  assign exp_726 = exp_725 | exp_684;
  assign exp_725 = exp_724 | exp_678;
  assign exp_724 = exp_723 | exp_676;
  assign exp_723 = exp_722 | exp_682;
  assign exp_722 = exp_721 | exp_680;
  assign exp_721 = exp_672 | exp_674;
  assign exp_672 = exp_669 == exp_671;
  assign exp_671 = 19;
  assign exp_674 = exp_669 == exp_673;
  assign exp_673 = 51;
  assign exp_676 = exp_669 == exp_675;
  assign exp_675 = 55;
  assign exp_678 = exp_669 == exp_677;
  assign exp_677 = 23;
  assign exp_1129 = exp_1128 & exp_888;

  reg [0:0] exp_1128_reg;
  always@(*) begin
    case (exp_914)
      0:exp_1128_reg <= exp_1125;
      1:exp_1128_reg <= exp_1126;
      default:exp_1128_reg <= exp_1127;
    endcase
  end
  assign exp_1128 = exp_1128_reg;
  assign exp_914 = exp_888 & exp_913;
  assign exp_888 = exp_886 & exp_887;
  assign exp_886 = exp_884 == exp_885;
  assign exp_884 = exp_667[6:0];
  assign exp_885 = 51;
  assign exp_887 = exp_667[25:25];
  assign exp_913 = exp_883[2:2];
  assign exp_883 = exp_667[14:12];
  assign exp_1127 = 0;
  assign exp_1125 = exp_1118 & exp_888;
  assign exp_1118 = exp_1033 == exp_1117;

      reg [2:0] exp_1033_reg = 0;
      always@(posedge clk) begin
        if (exp_1029) begin
          exp_1033_reg <= exp_1040;
        end
      end
      assign exp_1033 = exp_1033_reg;
    
  reg [2:0] exp_1040_reg;
  always@(*) begin
    case (exp_1035)
      0:exp_1040_reg <= exp_1037;
      1:exp_1040_reg <= exp_1038;
      default:exp_1040_reg <= exp_1039;
    endcase
  end
  assign exp_1040 = exp_1040_reg;
  assign exp_1035 = exp_1033 == exp_1034;
  assign exp_1034 = 4;
  assign exp_1039 = 0;
  assign exp_1037 = exp_1033 + exp_1036;
  assign exp_1036 = 1;
  assign exp_1038 = 0;
  assign exp_1029 = exp_888 & exp_1028;
  assign exp_1028 = ~exp_1027;
  assign exp_1027 = exp_883[2:2];
  assign exp_1117 = 4;
  assign exp_1126 = exp_936 & exp_888;
  assign exp_936 = exp_920 == exp_935;

      reg [5:0] exp_920_reg = 0;
      always@(posedge clk) begin
        if (exp_914) begin
          exp_920_reg <= exp_927;
        end
      end
      assign exp_920 = exp_920_reg;
    
  reg [5:0] exp_927_reg;
  always@(*) begin
    case (exp_922)
      0:exp_927_reg <= exp_924;
      1:exp_927_reg <= exp_925;
      default:exp_927_reg <= exp_926;
    endcase
  end
  assign exp_927 = exp_927_reg;
  assign exp_922 = exp_920 == exp_921;
  assign exp_921 = 37;
  assign exp_926 = 0;
  assign exp_924 = exp_920 + exp_923;
  assign exp_923 = 1;
  assign exp_925 = 0;
  assign exp_935 = 37;

      reg [0:0] exp_547_reg = 0;
      always@(posedge clk) begin
        if (exp_539) begin
          exp_547_reg <= exp_546;
        end
      end
      assign exp_547 = exp_547_reg;
      assign exp_546 = exp_544 & exp_545;

      reg [0:0] exp_544_reg = 0;
      always@(posedge clk) begin
        if (exp_539) begin
          exp_544_reg <= exp_543;
        end
      end
      assign exp_544 = exp_544_reg;
      assign exp_543 = exp_541 & exp_542;
  assign exp_541 = 1;
  assign exp_542 = ~exp_540;
  assign exp_540 = exp_1153;
  assign exp_1153 = exp_547 & exp_844;
  assign exp_539 = ~exp_538;
  assign exp_538 = exp_1157;
  assign exp_1157 = exp_547 & exp_1156;
  assign exp_1156 = exp_1155 | exp_1131;
  assign exp_1155 = exp_525 & exp_1154;
  assign exp_1154 = ~exp_524;
  assign exp_524 = exp_528;
  assign exp_528 = exp_537;
  assign exp_537 = exp_494 & exp_534;
  assign exp_494 = exp_473 | exp_493;
  assign exp_473 = exp_321 | exp_472;
  assign exp_321 = exp_204 | exp_320;
  assign exp_204 = exp_163 | exp_203;
  assign exp_163 = exp_34 | exp_162;
  assign exp_34 = exp_15 | exp_33;
  assign exp_15 = 0;
  assign exp_33 = exp_27 & exp_21;
  assign exp_27 = exp_25 == exp_26;
  assign exp_25 = exp_9[31:24];
  assign exp_9 = exp_532;

      reg [31:0] exp_532_reg = 0;
      always@(posedge clk) begin
        if (exp_529) begin
          exp_532_reg <= exp_521;
        end
      end
      assign exp_532 = exp_532_reg;
      assign exp_521 = exp_738;
  assign exp_738 = exp_737 + exp_736;
  assign exp_737 = 0;
  assign exp_736 = exp_659 + exp_735;
  assign exp_735 = $signed(exp_734);
  assign exp_734 = exp_733 + exp_732;
  assign exp_733 = 0;

  reg [11:0] exp_732_reg;
  always@(*) begin
    case (exp_686)
      0:exp_732_reg <= exp_727;
      1:exp_732_reg <= exp_730;
      default:exp_732_reg <= exp_731;
    endcase
  end
  assign exp_732 = exp_732_reg;
  assign exp_686 = exp_669 == exp_685;
  assign exp_685 = 35;
  assign exp_731 = 0;
  assign exp_727 = exp_667[31:20];
  assign exp_730 = {exp_728, exp_729};  assign exp_728 = exp_667[31:25];
  assign exp_729 = exp_667[11:7];
  assign exp_529 = 1;
  assign exp_26 = 0;
  assign exp_21 = exp_146;

  reg [0:0] exp_146_reg;
  always@(*) begin
    case (exp_23)
      0:exp_146_reg <= exp_140;
      1:exp_146_reg <= exp_125;
      default:exp_146_reg <= exp_145;
    endcase
  end
  assign exp_146 = exp_146_reg;
  assign exp_23 = exp_12;
  assign exp_12 = exp_535;

      reg [0:0] exp_535_reg = 0;
      always@(posedge clk) begin
        if (exp_529) begin
          exp_535_reg <= exp_526;
        end
      end
      assign exp_535 = exp_535_reg;
      assign exp_526 = exp_821;
  assign exp_821 = exp_820 + exp_686;
  assign exp_820 = 0;
  assign exp_145 = 0;

      reg [0:0] exp_140_reg = 0;
      always@(posedge clk) begin
        if (exp_139) begin
          exp_140_reg <= exp_144;
        end
      end
      assign exp_140 = exp_140_reg;
      assign exp_144 = exp_142 & exp_143;
  assign exp_142 = exp_22 & exp_141;
  assign exp_22 = exp_28;
  assign exp_28 = exp_11 & exp_27;
  assign exp_141 = ~exp_23;
  assign exp_143 = ~exp_140;
  assign exp_139 = 1;
  assign exp_125 = 1;
  assign exp_162 = exp_156 & exp_150;
  assign exp_156 = exp_154 == exp_155;
  assign exp_154 = exp_9[31:24];
  assign exp_155 = 1;
  assign exp_150 = exp_184;
  assign exp_184 = 1;
  assign exp_203 = exp_197 & exp_191;
  assign exp_197 = exp_195 == exp_196;
  assign exp_195 = exp_9[31:24];
  assign exp_196 = 2;
  assign exp_191 = exp_220;

      reg [0:0] exp_220_reg = 0;
      always@(posedge clk) begin
        if (exp_219) begin
          exp_220_reg <= exp_302;
        end
      end
      assign exp_220 = exp_220_reg;
    
  reg [0:0] exp_302_reg;
  always@(*) begin
    case (exp_300)
      0:exp_302_reg <= exp_292;
      1:exp_302_reg <= exp_243;
      default:exp_302_reg <= exp_301;
    endcase
  end
  assign exp_302 = exp_302_reg;
  assign exp_300 = exp_296 & exp_206;
  assign exp_296 = exp_244 & exp_295;
  assign exp_244 = 1;
  assign exp_295 = exp_214 == exp_294;

      reg [2:0] exp_214_reg = 0;
      always@(posedge clk) begin
        if (exp_213) begin
          exp_214_reg <= exp_299;
        end
      end
      assign exp_214 = exp_214_reg;
    
  reg [2:0] exp_299_reg;
  always@(*) begin
    case (exp_297)
      0:exp_299_reg <= exp_289;
      1:exp_299_reg <= exp_242;
      default:exp_299_reg <= exp_298;
    endcase
  end
  assign exp_299 = exp_299_reg;
  assign exp_297 = exp_296 & exp_206;
  assign exp_206 = exp_192 & exp_205;
  assign exp_192 = exp_198;
  assign exp_198 = exp_11 & exp_197;
  assign exp_205 = ~exp_193;
  assign exp_193 = exp_12;
  assign exp_298 = 0;

  reg [2:0] exp_289_reg;
  always@(*) begin
    case (exp_287)
      0:exp_289_reg <= exp_274;
      1:exp_289_reg <= exp_240;
      default:exp_289_reg <= exp_288;
    endcase
  end
  assign exp_289 = exp_289_reg;
  assign exp_287 = exp_286 & exp_212;
  assign exp_286 = exp_244 & exp_285;
  assign exp_285 = exp_214 == exp_284;
  assign exp_284 = 2;

      reg [0:0] exp_212_reg = 1;
      always@(posedge clk) begin
        if (exp_211) begin
          exp_212_reg <= exp_210;
        end
      end
      assign exp_212 = exp_212_reg;
    
      reg [0:0] exp_210_reg = 1;
      always@(posedge clk) begin
        if (exp_209) begin
          exp_210_reg <= exp_208;
        end
      end
      assign exp_210 = exp_210_reg;
    
      reg [0:0] exp_208_reg = 1;
      always@(posedge clk) begin
        if (exp_207) begin
          exp_208_reg <= exp_7;
        end
      end
      assign exp_208 = exp_208_reg;
      assign exp_7 = stdin_rx;
  assign exp_207 = 1;
  assign exp_209 = 1;
  assign exp_211 = 1;
  assign exp_288 = 0;

  reg [2:0] exp_274_reg;
  always@(*) begin
    case (exp_272)
      0:exp_274_reg <= exp_251;
      1:exp_274_reg <= exp_235;
      default:exp_274_reg <= exp_273;
    endcase
  end
  assign exp_274 = exp_274_reg;
  assign exp_272 = exp_268 & exp_233;
  assign exp_268 = exp_261 & exp_228;
  assign exp_261 = exp_244 & exp_260;
  assign exp_260 = exp_214 == exp_259;
  assign exp_259 = 1;
  assign exp_228 = exp_222 == exp_227;

      reg [9:0] exp_222_reg = 0;
      always@(posedge clk) begin
        if (exp_221) begin
          exp_222_reg <= exp_282;
        end
      end
      assign exp_222 = exp_222_reg;
    
  reg [9:0] exp_282_reg;
  always@(*) begin
    case (exp_280)
      0:exp_282_reg <= exp_271;
      1:exp_282_reg <= exp_239;
      default:exp_282_reg <= exp_281;
    endcase
  end
  assign exp_282 = exp_282_reg;
  assign exp_280 = exp_261 & exp_279;
  assign exp_279 = ~exp_228;
  assign exp_281 = 0;

  reg [9:0] exp_271_reg;
  always@(*) begin
    case (exp_269)
      0:exp_271_reg <= exp_267;
      1:exp_271_reg <= exp_234;
      default:exp_271_reg <= exp_270;
    endcase
  end
  assign exp_271 = exp_271_reg;
  assign exp_269 = exp_268 & exp_233;
  assign exp_233 = exp_216 == exp_232;

      reg [2:0] exp_216_reg = 0;
      always@(posedge clk) begin
        if (exp_215) begin
          exp_216_reg <= exp_278;
        end
      end
      assign exp_216 = exp_216_reg;
    
  reg [2:0] exp_278_reg;
  always@(*) begin
    case (exp_276)
      0:exp_278_reg <= exp_257;
      1:exp_278_reg <= exp_237;
      default:exp_278_reg <= exp_277;
    endcase
  end
  assign exp_278 = exp_278_reg;
  assign exp_276 = exp_268 & exp_275;
  assign exp_275 = ~exp_233;
  assign exp_277 = 0;

  reg [2:0] exp_257_reg;
  always@(*) begin
    case (exp_255)
      0:exp_257_reg <= exp_216;
      1:exp_257_reg <= exp_226;
      default:exp_257_reg <= exp_256;
    endcase
  end
  assign exp_257 = exp_257_reg;
  assign exp_255 = exp_248 & exp_223;
  assign exp_248 = exp_244 & exp_247;
  assign exp_247 = exp_214 == exp_246;
  assign exp_246 = 0;
  assign exp_223 = ~exp_212;
  assign exp_256 = 0;
  assign exp_226 = 0;
  assign exp_237 = exp_216 + exp_236;
  assign exp_236 = 1;
  assign exp_215 = 1;
  assign exp_232 = 7;
  assign exp_270 = 0;

  reg [9:0] exp_267_reg;
  always@(*) begin
    case (exp_265)
      0:exp_267_reg <= exp_254;
      1:exp_267_reg <= exp_231;
      default:exp_267_reg <= exp_266;
    endcase
  end
  assign exp_267 = exp_267_reg;
  assign exp_265 = exp_261 & exp_228;
  assign exp_266 = 0;

  reg [9:0] exp_254_reg;
  always@(*) begin
    case (exp_252)
      0:exp_254_reg <= exp_222;
      1:exp_254_reg <= exp_225;
      default:exp_254_reg <= exp_253;
    endcase
  end
  assign exp_254 = exp_254_reg;
  assign exp_252 = exp_248 & exp_223;
  assign exp_253 = 0;
  assign exp_225 = 650;
  assign exp_231 = 433;
  assign exp_234 = 433;
  assign exp_239 = exp_222 - exp_238;
  assign exp_238 = 1;
  assign exp_221 = 1;
  assign exp_227 = 0;
  assign exp_273 = 0;

  reg [2:0] exp_251_reg;
  always@(*) begin
    case (exp_249)
      0:exp_251_reg <= exp_214;
      1:exp_251_reg <= exp_224;
      default:exp_251_reg <= exp_250;
    endcase
  end
  assign exp_251 = exp_251_reg;
  assign exp_249 = exp_248 & exp_223;
  assign exp_250 = 0;
  assign exp_224 = 1;
  assign exp_235 = 2;
  assign exp_240 = 4;
  assign exp_242 = 0;
  assign exp_213 = 1;
  assign exp_294 = 4;
  assign exp_301 = 0;

  reg [0:0] exp_292_reg;
  always@(*) begin
    case (exp_290)
      0:exp_292_reg <= exp_220;
      1:exp_292_reg <= exp_241;
      default:exp_292_reg <= exp_291;
    endcase
  end
  assign exp_292 = exp_292_reg;
  assign exp_290 = exp_286 & exp_212;
  assign exp_291 = 0;
  assign exp_241 = 1;
  assign exp_243 = 0;
  assign exp_219 = 1;
  assign exp_320 = exp_314 & exp_308;
  assign exp_314 = exp_312 == exp_313;
  assign exp_312 = exp_9[31:24];
  assign exp_313 = 3;
  assign exp_308 = exp_331;

      reg [0:0] exp_331_reg = 1;
      always@(posedge clk) begin
        if (exp_330) begin
          exp_331_reg <= exp_450;
        end
      end
      assign exp_331 = exp_331_reg;
    
  reg [0:0] exp_450_reg;
  always@(*) begin
    case (exp_448)
      0:exp_450_reg <= exp_386;
      1:exp_450_reg <= exp_367;
      default:exp_450_reg <= exp_449;
    endcase
  end
  assign exp_450 = exp_450_reg;
  assign exp_448 = exp_444 & exp_365;
  assign exp_449 = 0;

  reg [0:0] exp_386_reg;
  always@(*) begin
    case (exp_384)
      0:exp_386_reg <= exp_331;
      1:exp_386_reg <= exp_338;
      default:exp_386_reg <= exp_385;
    endcase
  end
  assign exp_386 = exp_386_reg;
  assign exp_384 = exp_374 & exp_323;
  assign exp_385 = 0;
  assign exp_338 = 0;
  assign exp_367 = 1;
  assign exp_330 = 1;
  assign exp_472 = exp_466 & exp_460;
  assign exp_466 = exp_464 == exp_465;
  assign exp_464 = exp_9[31:24];
  assign exp_465 = 4;
  assign exp_460 = exp_477;
  assign exp_477 = 1;
  assign exp_493 = exp_487 & exp_481;
  assign exp_487 = exp_485 == exp_486;
  assign exp_485 = exp_9[31:24];
  assign exp_486 = 5;
  assign exp_481 = exp_520;
  assign exp_520 = 1;
  assign exp_1131 = exp_888 & exp_1130;
  assign exp_1130 = ~exp_1128;
  assign exp_545 = ~exp_540;
  assign exp_588 = 0;

  //Create RAM
  reg [31:0] exp_560_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_558) begin
      exp_560_ram[exp_554] <= exp_556;
    end
  end
  assign exp_560 = exp_560_ram[exp_555];
  assign exp_559 = exp_568;
  assign exp_568 = 1;
  assign exp_555 = exp_552;
  assign exp_558 = exp_1137;
  assign exp_1137 = exp_1136 & exp_539;
  assign exp_1136 = exp_1134 & exp_547;
  assign exp_554 = exp_1135;
  assign exp_556 = exp_1133;

  reg [31:0] exp_1133_reg;
  always@(*) begin
    case (exp_1129)
      0:exp_1133_reg <= exp_769;
      1:exp_1133_reg <= exp_1124;
      default:exp_1133_reg <= exp_1132;
    endcase
  end
  assign exp_1133 = exp_1133_reg;
  assign exp_1132 = 0;

  reg [31:0] exp_769_reg;
  always@(*) begin
    case (exp_684)
      0:exp_769_reg <= exp_720;
      1:exp_769_reg <= exp_767;
      default:exp_769_reg <= exp_768;
    endcase
  end
  assign exp_769 = exp_769_reg;
  assign exp_768 = 0;

  reg [31:0] exp_720_reg;
  always@(*) begin
    case (exp_663)
      0:exp_720_reg <= exp_699;
      1:exp_720_reg <= exp_701;
      2:exp_720_reg <= exp_717;
      3:exp_720_reg <= exp_718;
      4:exp_720_reg <= exp_710;
      5:exp_720_reg <= exp_714;
      6:exp_720_reg <= exp_715;
      7:exp_720_reg <= exp_716;
      default:exp_720_reg <= exp_719;
    endcase
  end
  assign exp_720 = exp_720_reg;

      reg [2:0] exp_663_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_663_reg <= exp_654;
        end
      end
      assign exp_663 = exp_663_reg;
    
  reg [2:0] exp_654_reg;
  always@(*) begin
    case (exp_651)
      0:exp_654_reg <= exp_641;
      1:exp_654_reg <= exp_652;
      default:exp_654_reg <= exp_653;
    endcase
  end
  assign exp_654 = exp_654_reg;
  assign exp_651 = exp_585 | exp_587;
  assign exp_585 = exp_575 == exp_584;
  assign exp_575 = exp_104[6:0];
  assign exp_584 = 111;
  assign exp_587 = exp_575 == exp_586;
  assign exp_586 = 103;
  assign exp_653 = 0;

  reg [2:0] exp_641_reg;
  always@(*) begin
    case (exp_583)
      0:exp_641_reg <= exp_628;
      1:exp_641_reg <= exp_639;
      default:exp_641_reg <= exp_640;
    endcase
  end
  assign exp_641 = exp_641_reg;
  assign exp_583 = exp_575 == exp_582;
  assign exp_582 = 23;
  assign exp_640 = 0;

  reg [2:0] exp_628_reg;
  always@(*) begin
    case (exp_581)
      0:exp_628_reg <= exp_577;
      1:exp_628_reg <= exp_626;
      default:exp_628_reg <= exp_627;
    endcase
  end
  assign exp_628 = exp_628_reg;
  assign exp_581 = exp_575 == exp_580;
  assign exp_580 = 55;
  assign exp_627 = 0;
  assign exp_577 = exp_104[14:12];
  assign exp_626 = 0;
  assign exp_639 = 0;
  assign exp_652 = 0;
  assign exp_658 = exp_539 & exp_544;
  assign exp_719 = 0;

  reg [31:0] exp_699_reg;
  always@(*) begin
    case (exp_665)
      0:exp_699_reg <= exp_696;
      1:exp_699_reg <= exp_697;
      default:exp_699_reg <= exp_698;
    endcase
  end
  assign exp_699 = exp_699_reg;

      reg [0:0] exp_665_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_665_reg <= exp_657;
        end
      end
      assign exp_665 = exp_665_reg;
      assign exp_657 = exp_643 & exp_656;
  assign exp_643 = exp_630 & exp_642;
  assign exp_630 = exp_616 & exp_629;
  assign exp_616 = exp_614 & exp_615;
  assign exp_614 = exp_104[30:30];
  assign exp_615 = ~exp_579;
  assign exp_579 = exp_575 == exp_578;
  assign exp_578 = 19;
  assign exp_629 = ~exp_581;
  assign exp_642 = ~exp_583;
  assign exp_656 = ~exp_655;
  assign exp_655 = exp_585 | exp_587;
  assign exp_698 = 0;
  assign exp_696 = exp_661 + exp_662;

      reg [31:0] exp_661_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_661_reg <= exp_647;
        end
      end
      assign exp_661 = exp_661_reg;
    
  reg [31:0] exp_647_reg;
  always@(*) begin
    case (exp_644)
      0:exp_647_reg <= exp_636;
      1:exp_647_reg <= exp_645;
      default:exp_647_reg <= exp_646;
    endcase
  end
  assign exp_647 = exp_647_reg;
  assign exp_644 = exp_585 | exp_587;
  assign exp_646 = 0;

  reg [31:0] exp_636_reg;
  always@(*) begin
    case (exp_583)
      0:exp_636_reg <= exp_622;
      1:exp_636_reg <= exp_634;
      default:exp_636_reg <= exp_635;
    endcase
  end
  assign exp_636 = exp_636_reg;
  assign exp_635 = 0;

  reg [31:0] exp_622_reg;
  always@(*) begin
    case (exp_581)
      0:exp_622_reg <= exp_597;
      1:exp_622_reg <= exp_620;
      default:exp_622_reg <= exp_621;
    endcase
  end
  assign exp_622 = exp_622_reg;
  assign exp_621 = 0;
  assign exp_620 = exp_618 << exp_619;
  assign exp_618 = exp_617;
  assign exp_617 = exp_104[31:12];
  assign exp_619 = 12;
  assign exp_634 = exp_632 << exp_633;
  assign exp_632 = exp_631;
  assign exp_631 = exp_104[31:12];
  assign exp_633 = 12;
  assign exp_645 = 4;

      reg [31:0] exp_662_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_662_reg <= exp_650;
        end
      end
      assign exp_662 = exp_662_reg;
    
  reg [31:0] exp_650_reg;
  always@(*) begin
    case (exp_648)
      0:exp_650_reg <= exp_638;
      1:exp_650_reg <= exp_551;
      default:exp_650_reg <= exp_649;
    endcase
  end
  assign exp_650 = exp_650_reg;
  assign exp_648 = exp_585 | exp_587;
  assign exp_649 = 0;

  reg [31:0] exp_638_reg;
  always@(*) begin
    case (exp_583)
      0:exp_638_reg <= exp_625;
      1:exp_638_reg <= exp_551;
      default:exp_638_reg <= exp_637;
    endcase
  end
  assign exp_638 = exp_638_reg;
  assign exp_637 = 0;

  reg [31:0] exp_625_reg;
  always@(*) begin
    case (exp_581)
      0:exp_625_reg <= exp_609;
      1:exp_625_reg <= exp_623;
      default:exp_625_reg <= exp_624;
    endcase
  end
  assign exp_625 = exp_625_reg;
  assign exp_624 = 0;

  reg [31:0] exp_609_reg;
  always@(*) begin
    case (exp_579)
      0:exp_609_reg <= exp_603;
      1:exp_609_reg <= exp_607;
      default:exp_609_reg <= exp_608;
    endcase
  end
  assign exp_609 = exp_609_reg;
  assign exp_608 = 0;

  reg [31:0] exp_603_reg;
  always@(*) begin
    case (exp_599)
      0:exp_603_reg <= exp_591;
      1:exp_603_reg <= exp_601;
      default:exp_603_reg <= exp_602;
    endcase
  end
  assign exp_603 = exp_603_reg;
  assign exp_599 = exp_574 == exp_598;
  assign exp_574 = exp_104[24:20];
  assign exp_598 = 0;
  assign exp_602 = 0;

  reg [31:0] exp_591_reg;
  always@(*) begin
    case (exp_571)
      0:exp_591_reg <= exp_567;
      1:exp_591_reg <= exp_572;
      default:exp_591_reg <= exp_590;
    endcase
  end
  assign exp_591 = exp_591_reg;
  assign exp_571 = exp_1147;
  assign exp_1147 = exp_1146 & exp_539;
  assign exp_1146 = exp_1145 & exp_547;
  assign exp_1145 = exp_1144 & exp_1134;
  assign exp_1144 = exp_553 == exp_1135;
  assign exp_553 = exp_104[24:20];
  assign exp_590 = 0;

  //Create RAM
  reg [31:0] exp_567_ram [31:0];

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_565) begin
      exp_567_ram[exp_561] <= exp_563;
    end
  end
  assign exp_567 = exp_567_ram[exp_562];
  assign exp_566 = exp_569;
  assign exp_569 = 1;
  assign exp_562 = exp_553;
  assign exp_565 = exp_1139;
  assign exp_1139 = exp_1138 & exp_539;
  assign exp_1138 = exp_1134 & exp_547;
  assign exp_561 = exp_1135;
  assign exp_563 = exp_1133;
  assign exp_572 = exp_1133;
  assign exp_601 = $signed(exp_600);
  assign exp_600 = 0;
  assign exp_607 = exp_604 + exp_606;
  assign exp_604 = 0;
  assign exp_606 = $signed(exp_605);
  assign exp_605 = exp_104[31:20];
  assign exp_623 = 0;

      reg [31:0] exp_551_reg = 0;
      always@(posedge clk) begin
        if (exp_550) begin
          exp_551_reg <= exp_549;
        end
      end
      assign exp_551 = exp_551_reg;
      assign exp_550 = exp_541 & exp_539;
  assign exp_697 = exp_661 - exp_662;
  assign exp_701 = exp_661 << exp_700;
  assign exp_700 = $signed(exp_695);
  assign exp_695 = exp_694 + exp_693;
  assign exp_694 = 0;
  assign exp_693 = exp_664;

      reg [4:0] exp_664_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_664_reg <= exp_613;
        end
      end
      assign exp_664 = exp_664_reg;
    
  reg [4:0] exp_613_reg;
  always@(*) begin
    case (exp_579)
      0:exp_613_reg <= exp_611;
      1:exp_613_reg <= exp_576;
      default:exp_613_reg <= exp_612;
    endcase
  end
  assign exp_613 = exp_613_reg;
  assign exp_612 = 0;
  assign exp_611 = exp_609[4:0];
  assign exp_576 = exp_104[24:20];
  assign exp_717 = $signed(exp_703);
  assign exp_703 = exp_702;
  assign exp_702 = $signed(exp_661) < $signed(exp_662);
  assign exp_718 = $signed(exp_709);
  assign exp_709 = exp_708;
  assign exp_708 = exp_705 < exp_707;
  assign exp_705 = exp_704 + exp_661;
  assign exp_704 = 0;
  assign exp_707 = exp_706 + exp_662;
  assign exp_706 = 0;
  assign exp_710 = exp_661 ^ exp_662;
  assign exp_714 = exp_713[31:0];
  assign exp_713 = $signed(exp_711) >>> $signed(exp_712);
  assign exp_711 = {exp_692, exp_661};
  reg [0:0] exp_692_reg;
  always@(*) begin
    case (exp_666)
      0:exp_692_reg <= exp_690;
      1:exp_692_reg <= exp_689;
      default:exp_692_reg <= exp_691;
    endcase
  end
  assign exp_692 = exp_692_reg;

      reg [0:0] exp_666_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_666_reg <= exp_610;
        end
      end
      assign exp_666 = exp_666_reg;
      assign exp_610 = exp_104[30:30];
  assign exp_691 = 0;
  assign exp_690 = 0;
  assign exp_689 = exp_661[31:31];
  assign exp_712 = $signed(exp_695);
  assign exp_715 = exp_661 | exp_662;
  assign exp_716 = exp_661 & exp_662;

  reg [31:0] exp_767_reg;
  always@(*) begin
    case (exp_670)
      0:exp_767_reg <= exp_757;
      1:exp_767_reg <= exp_760;
      2:exp_767_reg <= exp_523;
      3:exp_767_reg <= exp_761;
      4:exp_767_reg <= exp_762;
      5:exp_767_reg <= exp_763;
      6:exp_767_reg <= exp_764;
      7:exp_767_reg <= exp_765;
      default:exp_767_reg <= exp_766;
    endcase
  end
  assign exp_767 = exp_767_reg;
  assign exp_766 = 0;
  assign exp_757 = $signed(exp_756);
  assign exp_756 = exp_755 + exp_750;
  assign exp_755 = 0;

  reg [7:0] exp_750_reg;
  always@(*) begin
    case (exp_741)
      0:exp_750_reg <= exp_745;
      1:exp_750_reg <= exp_746;
      2:exp_750_reg <= exp_747;
      3:exp_750_reg <= exp_748;
      default:exp_750_reg <= exp_749;
    endcase
  end
  assign exp_750 = exp_750_reg;
  assign exp_741 = exp_740 + exp_739;
  assign exp_740 = 0;
  assign exp_739 = exp_738[1:0];
  assign exp_749 = 0;
  assign exp_745 = exp_523[7:0];
  assign exp_523 = exp_492;
  assign exp_492 = exp_471 | exp_491;
  assign exp_471 = exp_319 | exp_470;
  assign exp_319 = exp_202 | exp_318;
  assign exp_202 = exp_161 | exp_201;
  assign exp_161 = exp_32 | exp_160;
  assign exp_32 = exp_14 | exp_31;
  assign exp_14 = 0;

  reg [31:0] exp_31_reg;
  always@(*) begin
    case (exp_27)
      0:exp_31_reg <= exp_29;
      1:exp_31_reg <= exp_20;
      default:exp_31_reg <= exp_30;
    endcase
  end
  assign exp_31 = exp_31_reg;
  assign exp_30 = 0;
  assign exp_29 = 0;
  assign exp_20 = exp_127;

      reg [31:0] exp_127_reg = 0;
      always@(posedge clk) begin
        if (exp_126) begin
          exp_127_reg <= exp_138;
        end
      end
      assign exp_127 = exp_127_reg;
      assign exp_138 = {exp_137, exp_41};  assign exp_137 = {exp_136, exp_48};  assign exp_136 = {exp_62, exp_55};
  //Create RAM
  reg [7:0] exp_62_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_62_ram[0] = 0;
    exp_62_ram[1] = 0;
    exp_62_ram[2] = 0;
    exp_62_ram[3] = 0;
    exp_62_ram[4] = 0;
    exp_62_ram[5] = 0;
    exp_62_ram[6] = 0;
    exp_62_ram[7] = 0;
    exp_62_ram[8] = 0;
    exp_62_ram[9] = 0;
    exp_62_ram[10] = 0;
    exp_62_ram[11] = 0;
    exp_62_ram[12] = 0;
    exp_62_ram[13] = 0;
    exp_62_ram[14] = 0;
    exp_62_ram[15] = 0;
    exp_62_ram[16] = 0;
    exp_62_ram[17] = 0;
    exp_62_ram[18] = 0;
    exp_62_ram[19] = 0;
    exp_62_ram[20] = 0;
    exp_62_ram[21] = 0;
    exp_62_ram[22] = 0;
    exp_62_ram[23] = 0;
    exp_62_ram[24] = 0;
    exp_62_ram[25] = 0;
    exp_62_ram[26] = 0;
    exp_62_ram[27] = 0;
    exp_62_ram[28] = 0;
    exp_62_ram[29] = 0;
    exp_62_ram[30] = 0;
    exp_62_ram[31] = 0;
    exp_62_ram[32] = 252;
    exp_62_ram[33] = 22;
    exp_62_ram[34] = 0;
    exp_62_ram[35] = 0;
    exp_62_ram[36] = 0;
    exp_62_ram[37] = 0;
    exp_62_ram[38] = 0;
    exp_62_ram[39] = 0;
    exp_62_ram[40] = 40;
    exp_62_ram[41] = 0;
    exp_62_ram[42] = 185;
    exp_62_ram[43] = 14;
    exp_62_ram[44] = 0;
    exp_62_ram[45] = 12;
    exp_62_ram[46] = 15;
    exp_62_ram[47] = 0;
    exp_62_ram[48] = 0;
    exp_62_ram[49] = 0;
    exp_62_ram[50] = 0;
    exp_62_ram[51] = 0;
    exp_62_ram[52] = 2;
    exp_62_ram[53] = 0;
    exp_62_ram[54] = 64;
    exp_62_ram[55] = 0;
    exp_62_ram[56] = 0;
    exp_62_ram[57] = 0;
    exp_62_ram[58] = 0;
    exp_62_ram[59] = 0;
    exp_62_ram[60] = 0;
    exp_62_ram[61] = 1;
    exp_62_ram[62] = 3;
    exp_62_ram[63] = 1;
    exp_62_ram[64] = 1;
    exp_62_ram[65] = 1;
    exp_62_ram[66] = 3;
    exp_62_ram[67] = 0;
    exp_62_ram[68] = 2;
    exp_62_ram[69] = 1;
    exp_62_ram[70] = 0;
    exp_62_ram[71] = 0;
    exp_62_ram[72] = 1;
    exp_62_ram[73] = 255;
    exp_62_ram[74] = 1;
    exp_62_ram[75] = 0;
    exp_62_ram[76] = 255;
    exp_62_ram[77] = 1;
    exp_62_ram[78] = 64;
    exp_62_ram[79] = 3;
    exp_62_ram[80] = 1;
    exp_62_ram[81] = 1;
    exp_62_ram[82] = 3;
    exp_62_ram[83] = 1;
    exp_62_ram[84] = 0;
    exp_62_ram[85] = 2;
    exp_62_ram[86] = 0;
    exp_62_ram[87] = 0;
    exp_62_ram[88] = 0;
    exp_62_ram[89] = 255;
    exp_62_ram[90] = 1;
    exp_62_ram[91] = 0;
    exp_62_ram[92] = 255;
    exp_62_ram[93] = 1;
    exp_62_ram[94] = 0;
    exp_62_ram[95] = 0;
    exp_62_ram[96] = 14;
    exp_62_ram[97] = 1;
    exp_62_ram[98] = 1;
    exp_62_ram[99] = 242;
    exp_62_ram[100] = 1;
    exp_62_ram[101] = 243;
    exp_62_ram[102] = 0;
    exp_62_ram[103] = 0;
    exp_62_ram[104] = 2;
    exp_62_ram[105] = 0;
    exp_62_ram[106] = 12;
    exp_62_ram[107] = 15;
    exp_62_ram[108] = 1;
    exp_62_ram[109] = 0;
    exp_62_ram[110] = 0;
    exp_62_ram[111] = 0;
    exp_62_ram[112] = 0;
    exp_62_ram[113] = 2;
    exp_62_ram[114] = 0;
    exp_62_ram[115] = 64;
    exp_62_ram[116] = 10;
    exp_62_ram[117] = 65;
    exp_62_ram[118] = 0;
    exp_62_ram[119] = 1;
    exp_62_ram[120] = 1;
    exp_62_ram[121] = 1;
    exp_62_ram[122] = 1;
    exp_62_ram[123] = 3;
    exp_62_ram[124] = 3;
    exp_62_ram[125] = 1;
    exp_62_ram[126] = 0;
    exp_62_ram[127] = 2;
    exp_62_ram[128] = 0;
    exp_62_ram[129] = 1;
    exp_62_ram[130] = 1;
    exp_62_ram[131] = 255;
    exp_62_ram[132] = 1;
    exp_62_ram[133] = 1;
    exp_62_ram[134] = 255;
    exp_62_ram[135] = 1;
    exp_62_ram[136] = 65;
    exp_62_ram[137] = 3;
    exp_62_ram[138] = 1;
    exp_62_ram[139] = 1;
    exp_62_ram[140] = 3;
    exp_62_ram[141] = 1;
    exp_62_ram[142] = 0;
    exp_62_ram[143] = 2;
    exp_62_ram[144] = 0;
    exp_62_ram[145] = 0;
    exp_62_ram[146] = 0;
    exp_62_ram[147] = 255;
    exp_62_ram[148] = 1;
    exp_62_ram[149] = 0;
    exp_62_ram[150] = 255;
    exp_62_ram[151] = 1;
    exp_62_ram[152] = 0;
    exp_62_ram[153] = 0;
    exp_62_ram[154] = 1;
    exp_62_ram[155] = 1;
    exp_62_ram[156] = 244;
    exp_62_ram[157] = 1;
    exp_62_ram[158] = 244;
    exp_62_ram[159] = 0;
    exp_62_ram[160] = 0;
    exp_62_ram[161] = 0;
    exp_62_ram[162] = 0;
    exp_62_ram[163] = 0;
    exp_62_ram[164] = 1;
    exp_62_ram[165] = 0;
    exp_62_ram[166] = 3;
    exp_62_ram[167] = 1;
    exp_62_ram[168] = 1;
    exp_62_ram[169] = 1;
    exp_62_ram[170] = 3;
    exp_62_ram[171] = 1;
    exp_62_ram[172] = 0;
    exp_62_ram[173] = 2;
    exp_62_ram[174] = 0;
    exp_62_ram[175] = 0;
    exp_62_ram[176] = 1;
    exp_62_ram[177] = 255;
    exp_62_ram[178] = 1;
    exp_62_ram[179] = 0;
    exp_62_ram[180] = 255;
    exp_62_ram[181] = 1;
    exp_62_ram[182] = 64;
    exp_62_ram[183] = 3;
    exp_62_ram[184] = 1;
    exp_62_ram[185] = 1;
    exp_62_ram[186] = 3;
    exp_62_ram[187] = 1;
    exp_62_ram[188] = 2;
    exp_62_ram[189] = 0;
    exp_62_ram[190] = 0;
    exp_62_ram[191] = 0;
    exp_62_ram[192] = 1;
    exp_62_ram[193] = 255;
    exp_62_ram[194] = 1;
    exp_62_ram[195] = 0;
    exp_62_ram[196] = 255;
    exp_62_ram[197] = 1;
    exp_62_ram[198] = 1;
    exp_62_ram[199] = 64;
    exp_62_ram[200] = 0;
    exp_62_ram[201] = 235;
    exp_62_ram[202] = 24;
    exp_62_ram[203] = 0;
    exp_62_ram[204] = 4;
    exp_62_ram[205] = 15;
    exp_62_ram[206] = 0;
    exp_62_ram[207] = 0;
    exp_62_ram[208] = 0;
    exp_62_ram[209] = 0;
    exp_62_ram[210] = 185;
    exp_62_ram[211] = 0;
    exp_62_ram[212] = 0;
    exp_62_ram[213] = 2;
    exp_62_ram[214] = 0;
    exp_62_ram[215] = 64;
    exp_62_ram[216] = 2;
    exp_62_ram[217] = 0;
    exp_62_ram[218] = 238;
    exp_62_ram[219] = 0;
    exp_62_ram[220] = 0;
    exp_62_ram[221] = 239;
    exp_62_ram[222] = 1;
    exp_62_ram[223] = 1;
    exp_62_ram[224] = 252;
    exp_62_ram[225] = 1;
    exp_62_ram[226] = 251;
    exp_62_ram[227] = 0;
    exp_62_ram[228] = 0;
    exp_62_ram[229] = 0;
    exp_62_ram[230] = 0;
    exp_62_ram[231] = 1;
    exp_62_ram[232] = 3;
    exp_62_ram[233] = 0;
    exp_62_ram[234] = 0;
    exp_62_ram[235] = 0;
    exp_62_ram[236] = 0;
    exp_62_ram[237] = 1;
    exp_62_ram[238] = 1;
    exp_62_ram[239] = 1;
    exp_62_ram[240] = 3;
    exp_62_ram[241] = 1;
    exp_62_ram[242] = 0;
    exp_62_ram[243] = 3;
    exp_62_ram[244] = 0;
    exp_62_ram[245] = 1;
    exp_62_ram[246] = 1;
    exp_62_ram[247] = 255;
    exp_62_ram[248] = 1;
    exp_62_ram[249] = 1;
    exp_62_ram[250] = 255;
    exp_62_ram[251] = 1;
    exp_62_ram[252] = 65;
    exp_62_ram[253] = 3;
    exp_62_ram[254] = 3;
    exp_62_ram[255] = 1;
    exp_62_ram[256] = 2;
    exp_62_ram[257] = 1;
    exp_62_ram[258] = 1;
    exp_62_ram[259] = 0;
    exp_62_ram[260] = 0;
    exp_62_ram[261] = 1;
    exp_62_ram[262] = 1;
    exp_62_ram[263] = 255;
    exp_62_ram[264] = 1;
    exp_62_ram[265] = 1;
    exp_62_ram[266] = 255;
    exp_62_ram[267] = 1;
    exp_62_ram[268] = 1;
    exp_62_ram[269] = 0;
    exp_62_ram[270] = 0;
    exp_62_ram[271] = 255;
    exp_62_ram[272] = 0;
    exp_62_ram[273] = 1;
    exp_62_ram[274] = 0;
    exp_62_ram[275] = 1;
    exp_62_ram[276] = 65;
    exp_62_ram[277] = 2;
    exp_62_ram[278] = 2;
    exp_62_ram[279] = 1;
    exp_62_ram[280] = 2;
    exp_62_ram[281] = 0;
    exp_62_ram[282] = 1;
    exp_62_ram[283] = 2;
    exp_62_ram[284] = 0;
    exp_62_ram[285] = 1;
    exp_62_ram[286] = 1;
    exp_62_ram[287] = 0;
    exp_62_ram[288] = 2;
    exp_62_ram[289] = 206;
    exp_62_ram[290] = 0;
    exp_62_ram[291] = 255;
    exp_62_ram[292] = 0;
    exp_62_ram[293] = 1;
    exp_62_ram[294] = 0;
    exp_62_ram[295] = 0;
    exp_62_ram[296] = 1;
    exp_62_ram[297] = 0;
    exp_62_ram[298] = 218;
    exp_62_ram[299] = 255;
    exp_62_ram[300] = 204;
    exp_62_ram[301] = 0;
    exp_62_ram[302] = 0;
    exp_62_ram[303] = 218;
    exp_62_ram[304] = 0;
    exp_62_ram[305] = 255;
    exp_62_ram[306] = 1;
    exp_62_ram[307] = 0;
    exp_62_ram[308] = 0;
    exp_62_ram[309] = 0;
    exp_62_ram[310] = 127;
    exp_62_ram[311] = 1;
    exp_62_ram[312] = 127;
    exp_62_ram[313] = 1;
    exp_62_ram[314] = 0;
    exp_62_ram[315] = 0;
    exp_62_ram[316] = 127;
    exp_62_ram[317] = 1;
    exp_62_ram[318] = 1;
    exp_62_ram[319] = 0;
    exp_62_ram[320] = 8;
    exp_62_ram[321] = 0;
    exp_62_ram[322] = 0;
    exp_62_ram[323] = 1;
    exp_62_ram[324] = 0;
    exp_62_ram[325] = 254;
    exp_62_ram[326] = 8;
    exp_62_ram[327] = 0;
    exp_62_ram[328] = 0;
    exp_62_ram[329] = 0;
    exp_62_ram[330] = 0;
    exp_62_ram[331] = 4;
    exp_62_ram[332] = 0;
    exp_62_ram[333] = 0;
    exp_62_ram[334] = 3;
    exp_62_ram[335] = 4;
    exp_62_ram[336] = 255;
    exp_62_ram[337] = 0;
    exp_62_ram[338] = 255;
    exp_62_ram[339] = 0;
    exp_62_ram[340] = 0;
    exp_62_ram[341] = 0;
    exp_62_ram[342] = 0;
    exp_62_ram[343] = 254;
    exp_62_ram[344] = 0;
    exp_62_ram[345] = 253;
    exp_62_ram[346] = 2;
    exp_62_ram[347] = 252;
    exp_62_ram[348] = 255;
    exp_62_ram[349] = 0;
    exp_62_ram[350] = 0;
    exp_62_ram[351] = 0;
    exp_62_ram[352] = 0;
    exp_62_ram[353] = 254;
    exp_62_ram[354] = 251;
    exp_62_ram[355] = 252;
    exp_62_ram[356] = 254;
    exp_62_ram[357] = 247;
    exp_62_ram[358] = 248;
    exp_62_ram[359] = 0;
    exp_62_ram[360] = 248;
    exp_62_ram[361] = 255;
    exp_62_ram[362] = 0;
    exp_62_ram[363] = 0;
    exp_62_ram[364] = 0;
    exp_62_ram[365] = 6;
    exp_62_ram[366] = 42;
    exp_62_ram[367] = 65;
    exp_62_ram[368] = 0;
    exp_62_ram[369] = 64;
    exp_62_ram[370] = 4;
    exp_62_ram[371] = 0;
    exp_62_ram[372] = 64;
    exp_62_ram[373] = 1;
    exp_62_ram[374] = 0;
    exp_62_ram[375] = 0;
    exp_62_ram[376] = 0;
    exp_62_ram[377] = 0;
    exp_62_ram[378] = 0;
    exp_62_ram[379] = 0;
    exp_62_ram[380] = 1;
    exp_62_ram[381] = 0;
    exp_62_ram[382] = 0;
    exp_62_ram[383] = 0;
    exp_62_ram[384] = 1;
    exp_62_ram[385] = 0;
    exp_62_ram[386] = 255;
    exp_62_ram[387] = 0;
    exp_62_ram[388] = 0;
    exp_62_ram[389] = 252;
    exp_62_ram[390] = 0;
    exp_62_ram[391] = 0;
    exp_62_ram[392] = 252;
    exp_62_ram[393] = 254;
    exp_62_ram[394] = 0;
    exp_62_ram[395] = 0;
    exp_62_ram[396] = 0;
    exp_62_ram[397] = 1;
    exp_62_ram[398] = 1;
    exp_62_ram[399] = 1;
    exp_62_ram[400] = 0;
    exp_62_ram[401] = 24;
    exp_62_ram[402] = 0;
    exp_62_ram[403] = 0;
    exp_62_ram[404] = 0;
    exp_62_ram[405] = 8;
    exp_62_ram[406] = 0;
    exp_62_ram[407] = 32;
    exp_62_ram[408] = 0;
    exp_62_ram[409] = 67;
    exp_62_ram[410] = 65;
    exp_62_ram[411] = 67;
    exp_62_ram[412] = 9;
    exp_62_ram[413] = 0;
    exp_62_ram[414] = 0;
    exp_62_ram[415] = 3;
    exp_62_ram[416] = 2;
    exp_62_ram[417] = 7;
    exp_62_ram[418] = 2;
    exp_62_ram[419] = 255;
    exp_62_ram[420] = 65;
    exp_62_ram[421] = 0;
    exp_62_ram[422] = 0;
    exp_62_ram[423] = 0;
    exp_62_ram[424] = 0;
    exp_62_ram[425] = 1;
    exp_62_ram[426] = 1;
    exp_62_ram[427] = 0;
    exp_62_ram[428] = 1;
    exp_62_ram[429] = 0;
    exp_62_ram[430] = 0;
    exp_62_ram[431] = 1;
    exp_62_ram[432] = 1;
    exp_62_ram[433] = 0;
    exp_62_ram[434] = 0;
    exp_62_ram[435] = 0;
    exp_62_ram[436] = 0;
    exp_62_ram[437] = 2;
    exp_62_ram[438] = 0;
    exp_62_ram[439] = 24;
    exp_62_ram[440] = 2;
    exp_62_ram[441] = 248;
    exp_62_ram[442] = 253;
    exp_62_ram[443] = 0;
    exp_62_ram[444] = 0;
    exp_62_ram[445] = 251;
    exp_62_ram[446] = 67;
    exp_62_ram[447] = 3;
    exp_62_ram[448] = 3;
    exp_62_ram[449] = 0;
    exp_62_ram[450] = 0;
    exp_62_ram[451] = 17;
    exp_62_ram[452] = 0;
    exp_62_ram[453] = 0;
    exp_62_ram[454] = 0;
    exp_62_ram[455] = 0;
    exp_62_ram[456] = 0;
    exp_62_ram[457] = 65;
    exp_62_ram[458] = 12;
    exp_62_ram[459] = 0;
    exp_62_ram[460] = 0;
    exp_62_ram[461] = 0;
    exp_62_ram[462] = 0;
    exp_62_ram[463] = 0;
    exp_62_ram[464] = 3;
    exp_62_ram[465] = 2;
    exp_62_ram[466] = 9;
    exp_62_ram[467] = 255;
    exp_62_ram[468] = 0;
    exp_62_ram[469] = 2;
    exp_62_ram[470] = 65;
    exp_62_ram[471] = 1;
    exp_62_ram[472] = 0;
    exp_62_ram[473] = 0;
    exp_62_ram[474] = 255;
    exp_62_ram[475] = 255;
    exp_62_ram[476] = 0;
    exp_62_ram[477] = 0;
    exp_62_ram[478] = 2;
    exp_62_ram[479] = 0;
    exp_62_ram[480] = 0;
    exp_62_ram[481] = 0;
    exp_62_ram[482] = 0;
    exp_62_ram[483] = 0;
    exp_62_ram[484] = 0;
    exp_62_ram[485] = 0;
    exp_62_ram[486] = 0;
    exp_62_ram[487] = 0;
    exp_62_ram[488] = 0;
    exp_62_ram[489] = 255;
    exp_62_ram[490] = 255;
    exp_62_ram[491] = 67;
    exp_62_ram[492] = 0;
    exp_62_ram[493] = 65;
    exp_62_ram[494] = 0;
    exp_62_ram[495] = 1;
    exp_62_ram[496] = 0;
    exp_62_ram[497] = 0;
    exp_62_ram[498] = 237;
    exp_62_ram[499] = 253;
    exp_62_ram[500] = 0;
    exp_62_ram[501] = 0;
    exp_62_ram[502] = 249;
    exp_62_ram[503] = 0;
    exp_62_ram[504] = 0;
    exp_62_ram[505] = 0;
    exp_62_ram[506] = 235;
    exp_62_ram[507] = 2;
    exp_62_ram[508] = 2;
    exp_62_ram[509] = 64;
    exp_62_ram[510] = 0;
    exp_62_ram[511] = 254;
    exp_62_ram[512] = 0;
    exp_62_ram[513] = 0;
    exp_62_ram[514] = 0;
    exp_62_ram[515] = 0;
    exp_62_ram[516] = 0;
    exp_62_ram[517] = 0;
    exp_62_ram[518] = 0;
    exp_62_ram[519] = 0;
    exp_62_ram[520] = 254;
    exp_62_ram[521] = 2;
    exp_62_ram[522] = 2;
    exp_62_ram[523] = 64;
    exp_62_ram[524] = 0;
    exp_62_ram[525] = 254;
    exp_62_ram[526] = 0;
    exp_62_ram[527] = 0;
    exp_62_ram[528] = 0;
    exp_62_ram[529] = 0;
    exp_62_ram[530] = 0;
    exp_62_ram[531] = 0;
    exp_62_ram[532] = 0;
    exp_62_ram[533] = 0;
    exp_62_ram[534] = 254;
    exp_62_ram[535] = 0;
    exp_62_ram[536] = 2;
    exp_62_ram[537] = 15;
    exp_62_ram[538] = 0;
    exp_62_ram[539] = 0;
    exp_62_ram[540] = 0;
    exp_62_ram[541] = 2;
    exp_62_ram[542] = 64;
    exp_62_ram[543] = 0;
    exp_62_ram[544] = 185;
    exp_62_ram[545] = 0;
    exp_62_ram[546] = 0;
    exp_62_ram[547] = 64;
    exp_62_ram[548] = 0;
    exp_62_ram[549] = 1;
    exp_62_ram[550] = 1;
    exp_62_ram[551] = 252;
    exp_62_ram[552] = 1;
    exp_62_ram[553] = 252;
    exp_62_ram[554] = 77;
    exp_62_ram[555] = 117;
    exp_62_ram[556] = 100;
    exp_62_ram[557] = 70;
    exp_62_ram[558] = 97;
    exp_62_ram[559] = 0;
    exp_62_ram[560] = 70;
    exp_62_ram[561] = 97;
    exp_62_ram[562] = 114;
    exp_62_ram[563] = 74;
    exp_62_ram[564] = 117;
    exp_62_ram[565] = 103;
    exp_62_ram[566] = 79;
    exp_62_ram[567] = 111;
    exp_62_ram[568] = 99;
    exp_62_ram[569] = 0;
    exp_62_ram[570] = 108;
    exp_62_ram[571] = 111;
    exp_62_ram[572] = 33;
    exp_62_ram[573] = 0;
    exp_62_ram[574] = 110;
    exp_62_ram[575] = 32;
    exp_62_ram[576] = 103;
    exp_62_ram[577] = 114;
    exp_62_ram[578] = 114;
    exp_62_ram[579] = 109;
    exp_62_ram[580] = 46;
    exp_62_ram[581] = 0;
    exp_62_ram[582] = 110;
    exp_62_ram[583] = 32;
    exp_62_ram[584] = 32;
    exp_62_ram[585] = 111;
    exp_62_ram[586] = 0;
    exp_62_ram[587] = 45;
    exp_62_ram[588] = 32;
    exp_62_ram[589] = 101;
    exp_62_ram[590] = 32;
    exp_62_ram[591] = 116;
    exp_62_ram[592] = 105;
    exp_62_ram[593] = 105;
    exp_62_ram[594] = 32;
    exp_62_ram[595] = 111;
    exp_62_ram[596] = 0;
    exp_62_ram[597] = 45;
    exp_62_ram[598] = 32;
    exp_62_ram[599] = 101;
    exp_62_ram[600] = 32;
    exp_62_ram[601] = 116;
    exp_62_ram[602] = 105;
    exp_62_ram[603] = 105;
    exp_62_ram[604] = 32;
    exp_62_ram[605] = 111;
    exp_62_ram[606] = 0;
    exp_62_ram[607] = 45;
    exp_62_ram[608] = 32;
    exp_62_ram[609] = 101;
    exp_62_ram[610] = 32;
    exp_62_ram[611] = 105;
    exp_62_ram[612] = 32;
    exp_62_ram[613] = 49;
    exp_62_ram[614] = 99;
    exp_62_ram[615] = 0;
    exp_62_ram[616] = 45;
    exp_62_ram[617] = 32;
    exp_62_ram[618] = 101;
    exp_62_ram[619] = 32;
    exp_62_ram[620] = 105;
    exp_62_ram[621] = 32;
    exp_62_ram[622] = 49;
    exp_62_ram[623] = 99;
    exp_62_ram[624] = 0;
    exp_62_ram[625] = 114;
    exp_62_ram[626] = 0;
    exp_62_ram[627] = 116;
    exp_62_ram[628] = 0;
    exp_62_ram[629] = 58;
    exp_62_ram[630] = 0;
    exp_62_ram[631] = 114;
    exp_62_ram[632] = 0;
    exp_62_ram[633] = 117;
    exp_62_ram[634] = 0;
    exp_62_ram[635] = 105;
    exp_62_ram[636] = 86;
    exp_62_ram[637] = 109;
    exp_62_ram[638] = 0;
    exp_62_ram[639] = 32;
    exp_62_ram[640] = 108;
    exp_62_ram[641] = 111;
    exp_62_ram[642] = 0;
    exp_62_ram[643] = 75;
    exp_62_ram[644] = 104;
    exp_62_ram[645] = 105;
    exp_62_ram[646] = 0;
    exp_62_ram[647] = 84;
    exp_62_ram[648] = 32;
    exp_62_ram[649] = 116;
    exp_62_ram[650] = 105;
    exp_62_ram[651] = 105;
    exp_62_ram[652] = 0;
    exp_62_ram[653] = 87;
    exp_62_ram[654] = 32;
    exp_62_ram[655] = 99;
    exp_62_ram[656] = 0;
    exp_62_ram[657] = 69;
    exp_62_ram[658] = 109;
    exp_62_ram[659] = 97;
    exp_62_ram[660] = 110;
    exp_62_ram[661] = 0;
    exp_62_ram[662] = 80;
    exp_62_ram[663] = 68;
    exp_62_ram[664] = 0;
    exp_62_ram[665] = 111;
    exp_62_ram[666] = 111;
    exp_62_ram[667] = 105;
    exp_62_ram[668] = 58;
    exp_62_ram[669] = 0;
    exp_62_ram[670] = 0;
    exp_62_ram[671] = 103;
    exp_62_ram[672] = 77;
    exp_62_ram[673] = 105;
    exp_62_ram[674] = 0;
    exp_62_ram[675] = 61;
    exp_62_ram[676] = 61;
    exp_62_ram[677] = 61;
    exp_62_ram[678] = 10;
    exp_62_ram[679] = 0;
    exp_62_ram[680] = 87;
    exp_62_ram[681] = 108;
    exp_62_ram[682] = 116;
    exp_62_ram[683] = 103;
    exp_62_ram[684] = 87;
    exp_62_ram[685] = 101;
    exp_62_ram[686] = 103;
    exp_62_ram[687] = 40;
    exp_62_ram[688] = 53;
    exp_62_ram[689] = 101;
    exp_62_ram[690] = 32;
    exp_62_ram[691] = 100;
    exp_62_ram[692] = 32;
    exp_62_ram[693] = 104;
    exp_62_ram[694] = 46;
    exp_62_ram[695] = 49;
    exp_62_ram[696] = 0;
    exp_62_ram[697] = 82;
    exp_62_ram[698] = 101;
    exp_62_ram[699] = 114;
    exp_62_ram[700] = 45;
    exp_62_ram[701] = 32;
    exp_62_ram[702] = 46;
    exp_62_ram[703] = 0;
    exp_62_ram[704] = 82;
    exp_62_ram[705] = 32;
    exp_62_ram[706] = 116;
    exp_62_ram[707] = 115;
    exp_62_ram[708] = 105;
    exp_62_ram[709] = 116;
    exp_62_ram[710] = 117;
    exp_62_ram[711] = 32;
    exp_62_ram[712] = 62;
    exp_62_ram[713] = 108;
    exp_62_ram[714] = 44;
    exp_62_ram[715] = 100;
    exp_62_ram[716] = 44;
    exp_62_ram[717] = 103;
    exp_62_ram[718] = 101;
    exp_62_ram[719] = 32;
    exp_62_ram[720] = 10;
    exp_62_ram[721] = 0;
    exp_62_ram[722] = 82;
    exp_62_ram[723] = 114;
    exp_62_ram[724] = 115;
    exp_62_ram[725] = 111;
    exp_62_ram[726] = 40;
    exp_62_ram[727] = 122;
    exp_62_ram[728] = 101;
    exp_62_ram[729] = 32;
    exp_62_ram[730] = 100;
    exp_62_ram[731] = 32;
    exp_62_ram[732] = 104;
    exp_62_ram[733] = 46;
    exp_62_ram[734] = 97;
    exp_62_ram[735] = 0;
    exp_62_ram[736] = 100;
    exp_62_ram[737] = 46;
    exp_62_ram[738] = 0;
    exp_62_ram[739] = 0;
    exp_62_ram[740] = 0;
    exp_62_ram[741] = 2;
    exp_62_ram[742] = 3;
    exp_62_ram[743] = 4;
    exp_62_ram[744] = 4;
    exp_62_ram[745] = 5;
    exp_62_ram[746] = 5;
    exp_62_ram[747] = 5;
    exp_62_ram[748] = 5;
    exp_62_ram[749] = 6;
    exp_62_ram[750] = 6;
    exp_62_ram[751] = 6;
    exp_62_ram[752] = 6;
    exp_62_ram[753] = 6;
    exp_62_ram[754] = 6;
    exp_62_ram[755] = 6;
    exp_62_ram[756] = 6;
    exp_62_ram[757] = 7;
    exp_62_ram[758] = 7;
    exp_62_ram[759] = 7;
    exp_62_ram[760] = 7;
    exp_62_ram[761] = 7;
    exp_62_ram[762] = 7;
    exp_62_ram[763] = 7;
    exp_62_ram[764] = 7;
    exp_62_ram[765] = 7;
    exp_62_ram[766] = 7;
    exp_62_ram[767] = 7;
    exp_62_ram[768] = 7;
    exp_62_ram[769] = 7;
    exp_62_ram[770] = 7;
    exp_62_ram[771] = 7;
    exp_62_ram[772] = 7;
    exp_62_ram[773] = 8;
    exp_62_ram[774] = 8;
    exp_62_ram[775] = 8;
    exp_62_ram[776] = 8;
    exp_62_ram[777] = 8;
    exp_62_ram[778] = 8;
    exp_62_ram[779] = 8;
    exp_62_ram[780] = 8;
    exp_62_ram[781] = 8;
    exp_62_ram[782] = 8;
    exp_62_ram[783] = 8;
    exp_62_ram[784] = 8;
    exp_62_ram[785] = 8;
    exp_62_ram[786] = 8;
    exp_62_ram[787] = 8;
    exp_62_ram[788] = 8;
    exp_62_ram[789] = 8;
    exp_62_ram[790] = 8;
    exp_62_ram[791] = 8;
    exp_62_ram[792] = 8;
    exp_62_ram[793] = 8;
    exp_62_ram[794] = 8;
    exp_62_ram[795] = 8;
    exp_62_ram[796] = 8;
    exp_62_ram[797] = 8;
    exp_62_ram[798] = 8;
    exp_62_ram[799] = 8;
    exp_62_ram[800] = 8;
    exp_62_ram[801] = 8;
    exp_62_ram[802] = 8;
    exp_62_ram[803] = 8;
    exp_62_ram[804] = 8;
    exp_62_ram[805] = 253;
    exp_62_ram[806] = 2;
    exp_62_ram[807] = 3;
    exp_62_ram[808] = 252;
    exp_62_ram[809] = 253;
    exp_62_ram[810] = 254;
    exp_62_ram[811] = 254;
    exp_62_ram[812] = 0;
    exp_62_ram[813] = 0;
    exp_62_ram[814] = 2;
    exp_62_ram[815] = 3;
    exp_62_ram[816] = 0;
    exp_62_ram[817] = 253;
    exp_62_ram[818] = 2;
    exp_62_ram[819] = 3;
    exp_62_ram[820] = 252;
    exp_62_ram[821] = 252;
    exp_62_ram[822] = 253;
    exp_62_ram[823] = 254;
    exp_62_ram[824] = 253;
    exp_62_ram[825] = 254;
    exp_62_ram[826] = 0;
    exp_62_ram[827] = 253;
    exp_62_ram[828] = 0;
    exp_62_ram[829] = 2;
    exp_62_ram[830] = 3;
    exp_62_ram[831] = 0;
    exp_62_ram[832] = 254;
    exp_62_ram[833] = 0;
    exp_62_ram[834] = 0;
    exp_62_ram[835] = 2;
    exp_62_ram[836] = 254;
    exp_62_ram[837] = 0;
    exp_62_ram[838] = 238;
    exp_62_ram[839] = 0;
    exp_62_ram[840] = 254;
    exp_62_ram[841] = 250;
    exp_62_ram[842] = 0;
    exp_62_ram[843] = 0;
    exp_62_ram[844] = 1;
    exp_62_ram[845] = 1;
    exp_62_ram[846] = 2;
    exp_62_ram[847] = 0;
    exp_62_ram[848] = 255;
    exp_62_ram[849] = 0;
    exp_62_ram[850] = 0;
    exp_62_ram[851] = 1;
    exp_62_ram[852] = 0;
    exp_62_ram[853] = 237;
    exp_62_ram[854] = 0;
    exp_62_ram[855] = 243;
    exp_62_ram[856] = 0;
    exp_62_ram[857] = 0;
    exp_62_ram[858] = 0;
    exp_62_ram[859] = 0;
    exp_62_ram[860] = 1;
    exp_62_ram[861] = 0;
    exp_62_ram[862] = 253;
    exp_62_ram[863] = 2;
    exp_62_ram[864] = 2;
    exp_62_ram[865] = 3;
    exp_62_ram[866] = 252;
    exp_62_ram[867] = 252;
    exp_62_ram[868] = 254;
    exp_62_ram[869] = 2;
    exp_62_ram[870] = 254;
    exp_62_ram[871] = 0;
    exp_62_ram[872] = 254;
    exp_62_ram[873] = 253;
    exp_62_ram[874] = 0;
    exp_62_ram[875] = 0;
    exp_62_ram[876] = 253;
    exp_62_ram[877] = 0;
    exp_62_ram[878] = 240;
    exp_62_ram[879] = 253;
    exp_62_ram[880] = 254;
    exp_62_ram[881] = 0;
    exp_62_ram[882] = 0;
    exp_62_ram[883] = 252;
    exp_62_ram[884] = 254;
    exp_62_ram[885] = 0;
    exp_62_ram[886] = 2;
    exp_62_ram[887] = 2;
    exp_62_ram[888] = 3;
    exp_62_ram[889] = 0;
    exp_62_ram[890] = 254;
    exp_62_ram[891] = 0;
    exp_62_ram[892] = 0;
    exp_62_ram[893] = 2;
    exp_62_ram[894] = 254;
    exp_62_ram[895] = 0;
    exp_62_ram[896] = 238;
    exp_62_ram[897] = 0;
    exp_62_ram[898] = 254;
    exp_62_ram[899] = 246;
    exp_62_ram[900] = 0;
    exp_62_ram[901] = 238;
    exp_62_ram[902] = 0;
    exp_62_ram[903] = 0;
    exp_62_ram[904] = 234;
    exp_62_ram[905] = 0;
    exp_62_ram[906] = 0;
    exp_62_ram[907] = 1;
    exp_62_ram[908] = 1;
    exp_62_ram[909] = 2;
    exp_62_ram[910] = 0;
    exp_62_ram[911] = 254;
    exp_62_ram[912] = 0;
    exp_62_ram[913] = 2;
    exp_62_ram[914] = 254;
    exp_62_ram[915] = 254;
    exp_62_ram[916] = 4;
    exp_62_ram[917] = 0;
    exp_62_ram[918] = 254;
    exp_62_ram[919] = 5;
    exp_62_ram[920] = 0;
    exp_62_ram[921] = 254;
    exp_62_ram[922] = 6;
    exp_62_ram[923] = 0;
    exp_62_ram[924] = 254;
    exp_62_ram[925] = 7;
    exp_62_ram[926] = 0;
    exp_62_ram[927] = 0;
    exp_62_ram[928] = 0;
    exp_62_ram[929] = 0;
    exp_62_ram[930] = 0;
    exp_62_ram[931] = 1;
    exp_62_ram[932] = 2;
    exp_62_ram[933] = 0;
    exp_62_ram[934] = 254;
    exp_62_ram[935] = 0;
    exp_62_ram[936] = 2;
    exp_62_ram[937] = 254;
    exp_62_ram[938] = 254;
    exp_62_ram[939] = 6;
    exp_62_ram[940] = 0;
    exp_62_ram[941] = 254;
    exp_62_ram[942] = 7;
    exp_62_ram[943] = 0;
    exp_62_ram[944] = 0;
    exp_62_ram[945] = 0;
    exp_62_ram[946] = 0;
    exp_62_ram[947] = 0;
    exp_62_ram[948] = 1;
    exp_62_ram[949] = 2;
    exp_62_ram[950] = 0;
    exp_62_ram[951] = 254;
    exp_62_ram[952] = 0;
    exp_62_ram[953] = 0;
    exp_62_ram[954] = 2;
    exp_62_ram[955] = 254;
    exp_62_ram[956] = 254;
    exp_62_ram[957] = 250;
    exp_62_ram[958] = 0;
    exp_62_ram[959] = 0;
    exp_62_ram[960] = 254;
    exp_62_ram[961] = 254;
    exp_62_ram[962] = 0;
    exp_62_ram[963] = 254;
    exp_62_ram[964] = 0;
    exp_62_ram[965] = 1;
    exp_62_ram[966] = 1;
    exp_62_ram[967] = 2;
    exp_62_ram[968] = 0;
    exp_62_ram[969] = 246;
    exp_62_ram[970] = 8;
    exp_62_ram[971] = 8;
    exp_62_ram[972] = 8;
    exp_62_ram[973] = 10;
    exp_62_ram[974] = 0;
    exp_62_ram[975] = 1;
    exp_62_ram[976] = 252;
    exp_62_ram[977] = 0;
    exp_62_ram[978] = 252;
    exp_62_ram[979] = 1;
    exp_62_ram[980] = 252;
    exp_62_ram[981] = 0;
    exp_62_ram[982] = 250;
    exp_62_ram[983] = 250;
    exp_62_ram[984] = 250;
    exp_62_ram[985] = 252;
    exp_62_ram[986] = 251;
    exp_62_ram[987] = 251;
    exp_62_ram[988] = 251;
    exp_62_ram[989] = 252;
    exp_62_ram[990] = 252;
    exp_62_ram[991] = 252;
    exp_62_ram[992] = 252;
    exp_62_ram[993] = 253;
    exp_62_ram[994] = 253;
    exp_62_ram[995] = 246;
    exp_62_ram[996] = 247;
    exp_62_ram[997] = 247;
    exp_62_ram[998] = 246;
    exp_62_ram[999] = 246;
    exp_62_ram[1000] = 246;
    exp_62_ram[1001] = 246;
    exp_62_ram[1002] = 246;
    exp_62_ram[1003] = 248;
    exp_62_ram[1004] = 246;
    exp_62_ram[1005] = 0;
    exp_62_ram[1006] = 82;
    exp_62_ram[1007] = 254;
    exp_62_ram[1008] = 254;
    exp_62_ram[1009] = 251;
    exp_62_ram[1010] = 254;
    exp_62_ram[1011] = 254;
    exp_62_ram[1012] = 0;
    exp_62_ram[1013] = 14;
    exp_62_ram[1014] = 252;
    exp_62_ram[1015] = 252;
    exp_62_ram[1016] = 64;
    exp_62_ram[1017] = 252;
    exp_62_ram[1018] = 251;
    exp_62_ram[1019] = 251;
    exp_62_ram[1020] = 251;
    exp_62_ram[1021] = 252;
    exp_62_ram[1022] = 252;
    exp_62_ram[1023] = 252;
    exp_62_ram[1024] = 252;
    exp_62_ram[1025] = 253;
    exp_62_ram[1026] = 253;
    exp_62_ram[1027] = 246;
    exp_62_ram[1028] = 247;
    exp_62_ram[1029] = 247;
    exp_62_ram[1030] = 246;
    exp_62_ram[1031] = 246;
    exp_62_ram[1032] = 246;
    exp_62_ram[1033] = 246;
    exp_62_ram[1034] = 246;
    exp_62_ram[1035] = 248;
    exp_62_ram[1036] = 246;
    exp_62_ram[1037] = 0;
    exp_62_ram[1038] = 74;
    exp_62_ram[1039] = 254;
    exp_62_ram[1040] = 254;
    exp_62_ram[1041] = 1;
    exp_62_ram[1042] = 250;
    exp_62_ram[1043] = 0;
    exp_62_ram[1044] = 250;
    exp_62_ram[1045] = 1;
    exp_62_ram[1046] = 248;
    exp_62_ram[1047] = 0;
    exp_62_ram[1048] = 248;
    exp_62_ram[1049] = 248;
    exp_62_ram[1050] = 248;
    exp_62_ram[1051] = 252;
    exp_62_ram[1052] = 249;
    exp_62_ram[1053] = 249;
    exp_62_ram[1054] = 249;
    exp_62_ram[1055] = 249;
    exp_62_ram[1056] = 250;
    exp_62_ram[1057] = 250;
    exp_62_ram[1058] = 250;
    exp_62_ram[1059] = 250;
    exp_62_ram[1060] = 251;
    exp_62_ram[1061] = 246;
    exp_62_ram[1062] = 247;
    exp_62_ram[1063] = 247;
    exp_62_ram[1064] = 246;
    exp_62_ram[1065] = 246;
    exp_62_ram[1066] = 246;
    exp_62_ram[1067] = 246;
    exp_62_ram[1068] = 246;
    exp_62_ram[1069] = 248;
    exp_62_ram[1070] = 246;
    exp_62_ram[1071] = 0;
    exp_62_ram[1072] = 65;
    exp_62_ram[1073] = 254;
    exp_62_ram[1074] = 254;
    exp_62_ram[1075] = 249;
    exp_62_ram[1076] = 254;
    exp_62_ram[1077] = 254;
    exp_62_ram[1078] = 0;
    exp_62_ram[1079] = 125;
    exp_62_ram[1080] = 249;
    exp_62_ram[1081] = 250;
    exp_62_ram[1082] = 64;
    exp_62_ram[1083] = 248;
    exp_62_ram[1084] = 249;
    exp_62_ram[1085] = 249;
    exp_62_ram[1086] = 249;
    exp_62_ram[1087] = 249;
    exp_62_ram[1088] = 250;
    exp_62_ram[1089] = 250;
    exp_62_ram[1090] = 250;
    exp_62_ram[1091] = 250;
    exp_62_ram[1092] = 251;
    exp_62_ram[1093] = 246;
    exp_62_ram[1094] = 247;
    exp_62_ram[1095] = 247;
    exp_62_ram[1096] = 246;
    exp_62_ram[1097] = 246;
    exp_62_ram[1098] = 246;
    exp_62_ram[1099] = 246;
    exp_62_ram[1100] = 246;
    exp_62_ram[1101] = 248;
    exp_62_ram[1102] = 246;
    exp_62_ram[1103] = 0;
    exp_62_ram[1104] = 57;
    exp_62_ram[1105] = 254;
    exp_62_ram[1106] = 254;
    exp_62_ram[1107] = 0;
    exp_62_ram[1108] = 0;
    exp_62_ram[1109] = 0;
    exp_62_ram[1110] = 0;
    exp_62_ram[1111] = 1;
    exp_62_ram[1112] = 1;
    exp_62_ram[1113] = 1;
    exp_62_ram[1114] = 1;
    exp_62_ram[1115] = 2;
    exp_62_ram[1116] = 246;
    exp_62_ram[1117] = 247;
    exp_62_ram[1118] = 247;
    exp_62_ram[1119] = 246;
    exp_62_ram[1120] = 246;
    exp_62_ram[1121] = 246;
    exp_62_ram[1122] = 246;
    exp_62_ram[1123] = 246;
    exp_62_ram[1124] = 248;
    exp_62_ram[1125] = 246;
    exp_62_ram[1126] = 0;
    exp_62_ram[1127] = 52;
    exp_62_ram[1128] = 252;
    exp_62_ram[1129] = 252;
    exp_62_ram[1130] = 254;
    exp_62_ram[1131] = 253;
    exp_62_ram[1132] = 4;
    exp_62_ram[1133] = 254;
    exp_62_ram[1134] = 253;
    exp_62_ram[1135] = 0;
    exp_62_ram[1136] = 254;
    exp_62_ram[1137] = 253;
    exp_62_ram[1138] = 2;
    exp_62_ram[1139] = 254;
    exp_62_ram[1140] = 253;
    exp_62_ram[1141] = 0;
    exp_62_ram[1142] = 254;
    exp_62_ram[1143] = 253;
    exp_62_ram[1144] = 0;
    exp_62_ram[1145] = 254;
    exp_62_ram[1146] = 253;
    exp_62_ram[1147] = 0;
    exp_62_ram[1148] = 0;
    exp_62_ram[1149] = 0;
    exp_62_ram[1150] = 0;
    exp_62_ram[1151] = 0;
    exp_62_ram[1152] = 9;
    exp_62_ram[1153] = 9;
    exp_62_ram[1154] = 9;
    exp_62_ram[1155] = 10;
    exp_62_ram[1156] = 0;
    exp_62_ram[1157] = 248;
    exp_62_ram[1158] = 6;
    exp_62_ram[1159] = 6;
    exp_62_ram[1160] = 8;
    exp_62_ram[1161] = 250;
    exp_62_ram[1162] = 250;
    exp_62_ram[1163] = 252;
    exp_62_ram[1164] = 251;
    exp_62_ram[1165] = 251;
    exp_62_ram[1166] = 0;
    exp_62_ram[1167] = 103;
    exp_62_ram[1168] = 252;
    exp_62_ram[1169] = 253;
    exp_62_ram[1170] = 253;
    exp_62_ram[1171] = 253;
    exp_62_ram[1172] = 253;
    exp_62_ram[1173] = 254;
    exp_62_ram[1174] = 254;
    exp_62_ram[1175] = 254;
    exp_62_ram[1176] = 254;
    exp_62_ram[1177] = 248;
    exp_62_ram[1178] = 249;
    exp_62_ram[1179] = 249;
    exp_62_ram[1180] = 248;
    exp_62_ram[1181] = 248;
    exp_62_ram[1182] = 248;
    exp_62_ram[1183] = 248;
    exp_62_ram[1184] = 248;
    exp_62_ram[1185] = 250;
    exp_62_ram[1186] = 248;
    exp_62_ram[1187] = 0;
    exp_62_ram[1188] = 201;
    exp_62_ram[1189] = 0;
    exp_62_ram[1190] = 0;
    exp_62_ram[1191] = 7;
    exp_62_ram[1192] = 7;
    exp_62_ram[1193] = 8;
    exp_62_ram[1194] = 0;
    exp_62_ram[1195] = 254;
    exp_62_ram[1196] = 0;
    exp_62_ram[1197] = 2;
    exp_62_ram[1198] = 1;
    exp_62_ram[1199] = 254;
    exp_62_ram[1200] = 1;
    exp_62_ram[1201] = 0;
    exp_62_ram[1202] = 254;
    exp_62_ram[1203] = 254;
    exp_62_ram[1204] = 0;
    exp_62_ram[1205] = 254;
    exp_62_ram[1206] = 254;
    exp_62_ram[1207] = 254;
    exp_62_ram[1208] = 0;
    exp_62_ram[1209] = 254;
    exp_62_ram[1210] = 254;
    exp_62_ram[1211] = 254;
    exp_62_ram[1212] = 0;
    exp_62_ram[1213] = 0;
    exp_62_ram[1214] = 0;
    exp_62_ram[1215] = 254;
    exp_62_ram[1216] = 0;
    exp_62_ram[1217] = 254;
    exp_62_ram[1218] = 254;
    exp_62_ram[1219] = 0;
    exp_62_ram[1220] = 254;
    exp_62_ram[1221] = 254;
    exp_62_ram[1222] = 254;
    exp_62_ram[1223] = 0;
    exp_62_ram[1224] = 0;
    exp_62_ram[1225] = 1;
    exp_62_ram[1226] = 2;
    exp_62_ram[1227] = 0;
    exp_62_ram[1228] = 254;
    exp_62_ram[1229] = 0;
    exp_62_ram[1230] = 0;
    exp_62_ram[1231] = 2;
    exp_62_ram[1232] = 254;
    exp_62_ram[1233] = 254;
    exp_62_ram[1234] = 254;
    exp_62_ram[1235] = 254;
    exp_62_ram[1236] = 254;
    exp_62_ram[1237] = 254;
    exp_62_ram[1238] = 254;
    exp_62_ram[1239] = 254;
    exp_62_ram[1240] = 64;
    exp_62_ram[1241] = 0;
    exp_62_ram[1242] = 1;
    exp_62_ram[1243] = 64;
    exp_62_ram[1244] = 65;
    exp_62_ram[1245] = 0;
    exp_62_ram[1246] = 0;
    exp_62_ram[1247] = 0;
    exp_62_ram[1248] = 0;
    exp_62_ram[1249] = 0;
    exp_62_ram[1250] = 169;
    exp_62_ram[1251] = 0;
    exp_62_ram[1252] = 0;
    exp_62_ram[1253] = 0;
    exp_62_ram[1254] = 0;
    exp_62_ram[1255] = 1;
    exp_62_ram[1256] = 1;
    exp_62_ram[1257] = 2;
    exp_62_ram[1258] = 0;
    exp_62_ram[1259] = 254;
    exp_62_ram[1260] = 0;
    exp_62_ram[1261] = 2;
    exp_62_ram[1262] = 254;
    exp_62_ram[1263] = 254;
    exp_62_ram[1264] = 0;
    exp_62_ram[1265] = 2;
    exp_62_ram[1266] = 254;
    exp_62_ram[1267] = 6;
    exp_62_ram[1268] = 2;
    exp_62_ram[1269] = 0;
    exp_62_ram[1270] = 254;
    exp_62_ram[1271] = 25;
    exp_62_ram[1272] = 2;
    exp_62_ram[1273] = 0;
    exp_62_ram[1274] = 0;
    exp_62_ram[1275] = 0;
    exp_62_ram[1276] = 0;
    exp_62_ram[1277] = 0;
    exp_62_ram[1278] = 1;
    exp_62_ram[1279] = 2;
    exp_62_ram[1280] = 0;
    exp_62_ram[1281] = 254;
    exp_62_ram[1282] = 0;
    exp_62_ram[1283] = 0;
    exp_62_ram[1284] = 2;
    exp_62_ram[1285] = 254;
    exp_62_ram[1286] = 254;
    exp_62_ram[1287] = 249;
    exp_62_ram[1288] = 0;
    exp_62_ram[1289] = 0;
    exp_62_ram[1290] = 22;
    exp_62_ram[1291] = 0;
    exp_62_ram[1292] = 22;
    exp_62_ram[1293] = 0;
    exp_62_ram[1294] = 1;
    exp_62_ram[1295] = 1;
    exp_62_ram[1296] = 2;
    exp_62_ram[1297] = 0;
    exp_62_ram[1298] = 254;
    exp_62_ram[1299] = 0;
    exp_62_ram[1300] = 0;
    exp_62_ram[1301] = 2;
    exp_62_ram[1302] = 254;
    exp_62_ram[1303] = 254;
    exp_62_ram[1304] = 254;
    exp_62_ram[1305] = 0;
    exp_62_ram[1306] = 2;
    exp_62_ram[1307] = 254;
    exp_62_ram[1308] = 0;
    exp_62_ram[1309] = 0;
    exp_62_ram[1310] = 254;
    exp_62_ram[1311] = 0;
    exp_62_ram[1312] = 0;
    exp_62_ram[1313] = 254;
    exp_62_ram[1314] = 0;
    exp_62_ram[1315] = 0;
    exp_62_ram[1316] = 1;
    exp_62_ram[1317] = 3;
    exp_62_ram[1318] = 254;
    exp_62_ram[1319] = 0;
    exp_62_ram[1320] = 2;
    exp_62_ram[1321] = 254;
    exp_62_ram[1322] = 240;
    exp_62_ram[1323] = 0;
    exp_62_ram[1324] = 0;
    exp_62_ram[1325] = 1;
    exp_62_ram[1326] = 1;
    exp_62_ram[1327] = 1;
    exp_62_ram[1328] = 0;
    exp_62_ram[1329] = 1;
    exp_62_ram[1330] = 0;
    exp_62_ram[1331] = 1;
    exp_62_ram[1332] = 1;
    exp_62_ram[1333] = 2;
    exp_62_ram[1334] = 0;
    exp_62_ram[1335] = 249;
    exp_62_ram[1336] = 6;
    exp_62_ram[1337] = 6;
    exp_62_ram[1338] = 6;
    exp_62_ram[1339] = 7;
    exp_62_ram[1340] = 5;
    exp_62_ram[1341] = 5;
    exp_62_ram[1342] = 5;
    exp_62_ram[1343] = 5;
    exp_62_ram[1344] = 5;
    exp_62_ram[1345] = 5;
    exp_62_ram[1346] = 5;
    exp_62_ram[1347] = 5;
    exp_62_ram[1348] = 3;
    exp_62_ram[1349] = 7;
    exp_62_ram[1350] = 0;
    exp_62_ram[1351] = 0;
    exp_62_ram[1352] = 0;
    exp_62_ram[1353] = 250;
    exp_62_ram[1354] = 251;
    exp_62_ram[1355] = 123;
    exp_62_ram[1356] = 250;
    exp_62_ram[1357] = 1;
    exp_62_ram[1358] = 250;
    exp_62_ram[1359] = 250;
    exp_62_ram[1360] = 118;
    exp_62_ram[1361] = 251;
    exp_62_ram[1362] = 6;
    exp_62_ram[1363] = 251;
    exp_62_ram[1364] = 235;
    exp_62_ram[1365] = 0;
    exp_62_ram[1366] = 0;
    exp_62_ram[1367] = 24;
    exp_62_ram[1368] = 2;
    exp_62_ram[1369] = 248;
    exp_62_ram[1370] = 248;
    exp_62_ram[1371] = 251;
    exp_62_ram[1372] = 251;
    exp_62_ram[1373] = 249;
    exp_62_ram[1374] = 249;
    exp_62_ram[1375] = 0;
    exp_62_ram[1376] = 0;
    exp_62_ram[1377] = 0;
    exp_62_ram[1378] = 0;
    exp_62_ram[1379] = 0;
    exp_62_ram[1380] = 0;
    exp_62_ram[1381] = 0;
    exp_62_ram[1382] = 0;
    exp_62_ram[1383] = 250;
    exp_62_ram[1384] = 250;
    exp_62_ram[1385] = 251;
    exp_62_ram[1386] = 0;
    exp_62_ram[1387] = 250;
    exp_62_ram[1388] = 248;
    exp_62_ram[1389] = 0;
    exp_62_ram[1390] = 250;
    exp_62_ram[1391] = 1;
    exp_62_ram[1392] = 0;
    exp_62_ram[1393] = 251;
    exp_62_ram[1394] = 6;
    exp_62_ram[1395] = 251;
    exp_62_ram[1396] = 251;
    exp_62_ram[1397] = 231;
    exp_62_ram[1398] = 0;
    exp_62_ram[1399] = 0;
    exp_62_ram[1400] = 24;
    exp_62_ram[1401] = 2;
    exp_62_ram[1402] = 0;
    exp_62_ram[1403] = 0;
    exp_62_ram[1404] = 251;
    exp_62_ram[1405] = 251;
    exp_62_ram[1406] = 1;
    exp_62_ram[1407] = 0;
    exp_62_ram[1408] = 0;
    exp_62_ram[1409] = 1;
    exp_62_ram[1410] = 0;
    exp_62_ram[1411] = 0;
    exp_62_ram[1412] = 250;
    exp_62_ram[1413] = 250;
    exp_62_ram[1414] = 251;
    exp_62_ram[1415] = 0;
    exp_62_ram[1416] = 250;
    exp_62_ram[1417] = 249;
    exp_62_ram[1418] = 0;
    exp_62_ram[1419] = 0;
    exp_62_ram[1420] = 255;
    exp_62_ram[1421] = 0;
    exp_62_ram[1422] = 24;
    exp_62_ram[1423] = 2;
    exp_62_ram[1424] = 0;
    exp_62_ram[1425] = 65;
    exp_62_ram[1426] = 0;
    exp_62_ram[1427] = 251;
    exp_62_ram[1428] = 251;
    exp_62_ram[1429] = 1;
    exp_62_ram[1430] = 0;
    exp_62_ram[1431] = 0;
    exp_62_ram[1432] = 1;
    exp_62_ram[1433] = 0;
    exp_62_ram[1434] = 0;
    exp_62_ram[1435] = 250;
    exp_62_ram[1436] = 250;
    exp_62_ram[1437] = 0;
    exp_62_ram[1438] = 0;
    exp_62_ram[1439] = 225;
    exp_62_ram[1440] = 2;
    exp_62_ram[1441] = 0;
    exp_62_ram[1442] = 65;
    exp_62_ram[1443] = 0;
    exp_62_ram[1444] = 251;
    exp_62_ram[1445] = 251;
    exp_62_ram[1446] = 1;
    exp_62_ram[1447] = 0;
    exp_62_ram[1448] = 0;
    exp_62_ram[1449] = 1;
    exp_62_ram[1450] = 0;
    exp_62_ram[1451] = 0;
    exp_62_ram[1452] = 250;
    exp_62_ram[1453] = 250;
    exp_62_ram[1454] = 0;
    exp_62_ram[1455] = 0;
    exp_62_ram[1456] = 0;
    exp_62_ram[1457] = 64;
    exp_62_ram[1458] = 0;
    exp_62_ram[1459] = 0;
    exp_62_ram[1460] = 65;
    exp_62_ram[1461] = 0;
    exp_62_ram[1462] = 251;
    exp_62_ram[1463] = 251;
    exp_62_ram[1464] = 1;
    exp_62_ram[1465] = 0;
    exp_62_ram[1466] = 0;
    exp_62_ram[1467] = 1;
    exp_62_ram[1468] = 0;
    exp_62_ram[1469] = 0;
    exp_62_ram[1470] = 250;
    exp_62_ram[1471] = 250;
    exp_62_ram[1472] = 0;
    exp_62_ram[1473] = 0;
    exp_62_ram[1474] = 65;
    exp_62_ram[1475] = 0;
    exp_62_ram[1476] = 251;
    exp_62_ram[1477] = 251;
    exp_62_ram[1478] = 1;
    exp_62_ram[1479] = 0;
    exp_62_ram[1480] = 0;
    exp_62_ram[1481] = 1;
    exp_62_ram[1482] = 0;
    exp_62_ram[1483] = 0;
    exp_62_ram[1484] = 250;
    exp_62_ram[1485] = 250;
    exp_62_ram[1486] = 251;
    exp_62_ram[1487] = 251;
    exp_62_ram[1488] = 0;
    exp_62_ram[1489] = 0;
    exp_62_ram[1490] = 6;
    exp_62_ram[1491] = 6;
    exp_62_ram[1492] = 6;
    exp_62_ram[1493] = 6;
    exp_62_ram[1494] = 5;
    exp_62_ram[1495] = 5;
    exp_62_ram[1496] = 5;
    exp_62_ram[1497] = 5;
    exp_62_ram[1498] = 4;
    exp_62_ram[1499] = 4;
    exp_62_ram[1500] = 4;
    exp_62_ram[1501] = 4;
    exp_62_ram[1502] = 3;
    exp_62_ram[1503] = 7;
    exp_62_ram[1504] = 0;
    exp_62_ram[1505] = 246;
    exp_62_ram[1506] = 8;
    exp_62_ram[1507] = 8;
    exp_62_ram[1508] = 8;
    exp_62_ram[1509] = 9;
    exp_62_ram[1510] = 9;
    exp_62_ram[1511] = 10;
    exp_62_ram[1512] = 248;
    exp_62_ram[1513] = 249;
    exp_62_ram[1514] = 0;
    exp_62_ram[1515] = 0;
    exp_62_ram[1516] = 0;
    exp_62_ram[1517] = 0;
    exp_62_ram[1518] = 1;
    exp_62_ram[1519] = 1;
    exp_62_ram[1520] = 1;
    exp_62_ram[1521] = 1;
    exp_62_ram[1522] = 2;
    exp_62_ram[1523] = 250;
    exp_62_ram[1524] = 251;
    exp_62_ram[1525] = 251;
    exp_62_ram[1526] = 250;
    exp_62_ram[1527] = 250;
    exp_62_ram[1528] = 252;
    exp_62_ram[1529] = 252;
    exp_62_ram[1530] = 252;
    exp_62_ram[1531] = 252;
    exp_62_ram[1532] = 250;
    exp_62_ram[1533] = 251;
    exp_62_ram[1534] = 251;
    exp_62_ram[1535] = 251;
    exp_62_ram[1536] = 251;
    exp_62_ram[1537] = 252;
    exp_62_ram[1538] = 252;
    exp_62_ram[1539] = 252;
    exp_62_ram[1540] = 252;
    exp_62_ram[1541] = 246;
    exp_62_ram[1542] = 247;
    exp_62_ram[1543] = 247;
    exp_62_ram[1544] = 246;
    exp_62_ram[1545] = 246;
    exp_62_ram[1546] = 246;
    exp_62_ram[1547] = 246;
    exp_62_ram[1548] = 246;
    exp_62_ram[1549] = 248;
    exp_62_ram[1550] = 246;
    exp_62_ram[1551] = 0;
    exp_62_ram[1552] = 201;
    exp_62_ram[1553] = 252;
    exp_62_ram[1554] = 252;
    exp_62_ram[1555] = 252;
    exp_62_ram[1556] = 2;
    exp_62_ram[1557] = 253;
    exp_62_ram[1558] = 253;
    exp_62_ram[1559] = 255;
    exp_62_ram[1560] = 31;
    exp_62_ram[1561] = 255;
    exp_62_ram[1562] = 0;
    exp_62_ram[1563] = 0;
    exp_62_ram[1564] = 0;
    exp_62_ram[1565] = 0;
    exp_62_ram[1566] = 0;
    exp_62_ram[1567] = 0;
    exp_62_ram[1568] = 252;
    exp_62_ram[1569] = 252;
    exp_62_ram[1570] = 11;
    exp_62_ram[1571] = 252;
    exp_62_ram[1572] = 10;
    exp_62_ram[1573] = 250;
    exp_62_ram[1574] = 251;
    exp_62_ram[1575] = 251;
    exp_62_ram[1576] = 251;
    exp_62_ram[1577] = 251;
    exp_62_ram[1578] = 252;
    exp_62_ram[1579] = 252;
    exp_62_ram[1580] = 252;
    exp_62_ram[1581] = 252;
    exp_62_ram[1582] = 246;
    exp_62_ram[1583] = 247;
    exp_62_ram[1584] = 247;
    exp_62_ram[1585] = 246;
    exp_62_ram[1586] = 246;
    exp_62_ram[1587] = 246;
    exp_62_ram[1588] = 246;
    exp_62_ram[1589] = 246;
    exp_62_ram[1590] = 248;
    exp_62_ram[1591] = 246;
    exp_62_ram[1592] = 0;
    exp_62_ram[1593] = 228;
    exp_62_ram[1594] = 0;
    exp_62_ram[1595] = 0;
    exp_62_ram[1596] = 0;
    exp_62_ram[1597] = 225;
    exp_62_ram[1598] = 0;
    exp_62_ram[1599] = 0;
    exp_62_ram[1600] = 0;
    exp_62_ram[1601] = 0;
    exp_62_ram[1602] = 253;
    exp_62_ram[1603] = 253;
    exp_62_ram[1604] = 64;
    exp_62_ram[1605] = 0;
    exp_62_ram[1606] = 1;
    exp_62_ram[1607] = 64;
    exp_62_ram[1608] = 65;
    exp_62_ram[1609] = 0;
    exp_62_ram[1610] = 252;
    exp_62_ram[1611] = 252;
    exp_62_ram[1612] = 1;
    exp_62_ram[1613] = 253;
    exp_62_ram[1614] = 253;
    exp_62_ram[1615] = 252;
    exp_62_ram[1616] = 252;
    exp_62_ram[1617] = 0;
    exp_62_ram[1618] = 254;
    exp_62_ram[1619] = 0;
    exp_62_ram[1620] = 65;
    exp_62_ram[1621] = 0;
    exp_62_ram[1622] = 253;
    exp_62_ram[1623] = 253;
    exp_62_ram[1624] = 65;
    exp_62_ram[1625] = 0;
    exp_62_ram[1626] = 0;
    exp_62_ram[1627] = 65;
    exp_62_ram[1628] = 64;
    exp_62_ram[1629] = 0;
    exp_62_ram[1630] = 252;
    exp_62_ram[1631] = 252;
    exp_62_ram[1632] = 249;
    exp_62_ram[1633] = 246;
    exp_62_ram[1634] = 253;
    exp_62_ram[1635] = 253;
    exp_62_ram[1636] = 0;
    exp_62_ram[1637] = 114;
    exp_62_ram[1638] = 246;
    exp_62_ram[1639] = 246;
    exp_62_ram[1640] = 246;
    exp_62_ram[1641] = 246;
    exp_62_ram[1642] = 247;
    exp_62_ram[1643] = 247;
    exp_62_ram[1644] = 247;
    exp_62_ram[1645] = 247;
    exp_62_ram[1646] = 248;
    exp_62_ram[1647] = 0;
    exp_62_ram[1648] = 1;
    exp_62_ram[1649] = 1;
    exp_62_ram[1650] = 0;
    exp_62_ram[1651] = 0;
    exp_62_ram[1652] = 0;
    exp_62_ram[1653] = 0;
    exp_62_ram[1654] = 0;
    exp_62_ram[1655] = 2;
    exp_62_ram[1656] = 252;
    exp_62_ram[1657] = 0;
    exp_62_ram[1658] = 249;
    exp_62_ram[1659] = 0;
    exp_62_ram[1660] = 2;
    exp_62_ram[1661] = 7;
    exp_62_ram[1662] = 252;
    exp_62_ram[1663] = 6;
    exp_62_ram[1664] = 250;
    exp_62_ram[1665] = 251;
    exp_62_ram[1666] = 251;
    exp_62_ram[1667] = 251;
    exp_62_ram[1668] = 251;
    exp_62_ram[1669] = 252;
    exp_62_ram[1670] = 252;
    exp_62_ram[1671] = 252;
    exp_62_ram[1672] = 252;
    exp_62_ram[1673] = 246;
    exp_62_ram[1674] = 247;
    exp_62_ram[1675] = 247;
    exp_62_ram[1676] = 246;
    exp_62_ram[1677] = 246;
    exp_62_ram[1678] = 246;
    exp_62_ram[1679] = 246;
    exp_62_ram[1680] = 246;
    exp_62_ram[1681] = 248;
    exp_62_ram[1682] = 246;
    exp_62_ram[1683] = 0;
    exp_62_ram[1684] = 205;
    exp_62_ram[1685] = 0;
    exp_62_ram[1686] = 249;
    exp_62_ram[1687] = 2;
    exp_62_ram[1688] = 0;
    exp_62_ram[1689] = 249;
    exp_62_ram[1690] = 2;
    exp_62_ram[1691] = 253;
    exp_62_ram[1692] = 253;
    exp_62_ram[1693] = 0;
    exp_62_ram[1694] = 0;
    exp_62_ram[1695] = 9;
    exp_62_ram[1696] = 9;
    exp_62_ram[1697] = 9;
    exp_62_ram[1698] = 9;
    exp_62_ram[1699] = 8;
    exp_62_ram[1700] = 10;
    exp_62_ram[1701] = 0;
    exp_62_ram[1702] = 252;
    exp_62_ram[1703] = 2;
    exp_62_ram[1704] = 2;
    exp_62_ram[1705] = 3;
    exp_62_ram[1706] = 3;
    exp_62_ram[1707] = 3;
    exp_62_ram[1708] = 3;
    exp_62_ram[1709] = 3;
    exp_62_ram[1710] = 3;
    exp_62_ram[1711] = 4;
    exp_62_ram[1712] = 252;
    exp_62_ram[1713] = 254;
    exp_62_ram[1714] = 0;
    exp_62_ram[1715] = 0;
    exp_62_ram[1716] = 0;
    exp_62_ram[1717] = 237;
    exp_62_ram[1718] = 0;
    exp_62_ram[1719] = 0;
    exp_62_ram[1720] = 0;
    exp_62_ram[1721] = 0;
    exp_62_ram[1722] = 0;
    exp_62_ram[1723] = 0;
    exp_62_ram[1724] = 217;
    exp_62_ram[1725] = 0;
    exp_62_ram[1726] = 0;
    exp_62_ram[1727] = 252;
    exp_62_ram[1728] = 0;
    exp_62_ram[1729] = 254;
    exp_62_ram[1730] = 254;
    exp_62_ram[1731] = 253;
    exp_62_ram[1732] = 0;
    exp_62_ram[1733] = 252;
    exp_62_ram[1734] = 252;
    exp_62_ram[1735] = 0;
    exp_62_ram[1736] = 253;
    exp_62_ram[1737] = 0;
    exp_62_ram[1738] = 0;
    exp_62_ram[1739] = 252;
    exp_62_ram[1740] = 1;
    exp_62_ram[1741] = 1;
    exp_62_ram[1742] = 253;
    exp_62_ram[1743] = 0;
    exp_62_ram[1744] = 0;
    exp_62_ram[1745] = 0;
    exp_62_ram[1746] = 0;
    exp_62_ram[1747] = 0;
    exp_62_ram[1748] = 0;
    exp_62_ram[1749] = 3;
    exp_62_ram[1750] = 3;
    exp_62_ram[1751] = 3;
    exp_62_ram[1752] = 3;
    exp_62_ram[1753] = 2;
    exp_62_ram[1754] = 2;
    exp_62_ram[1755] = 2;
    exp_62_ram[1756] = 2;
    exp_62_ram[1757] = 4;
    exp_62_ram[1758] = 0;
    exp_62_ram[1759] = 253;
    exp_62_ram[1760] = 2;
    exp_62_ram[1761] = 2;
    exp_62_ram[1762] = 3;
    exp_62_ram[1763] = 3;
    exp_62_ram[1764] = 3;
    exp_62_ram[1765] = 252;
    exp_62_ram[1766] = 252;
    exp_62_ram[1767] = 241;
    exp_62_ram[1768] = 0;
    exp_62_ram[1769] = 0;
    exp_62_ram[1770] = 0;
    exp_62_ram[1771] = 237;
    exp_62_ram[1772] = 0;
    exp_62_ram[1773] = 0;
    exp_62_ram[1774] = 0;
    exp_62_ram[1775] = 0;
    exp_62_ram[1776] = 0;
    exp_62_ram[1777] = 0;
    exp_62_ram[1778] = 204;
    exp_62_ram[1779] = 0;
    exp_62_ram[1780] = 0;
    exp_62_ram[1781] = 254;
    exp_62_ram[1782] = 254;
    exp_62_ram[1783] = 253;
    exp_62_ram[1784] = 253;
    exp_62_ram[1785] = 254;
    exp_62_ram[1786] = 254;
    exp_62_ram[1787] = 64;
    exp_62_ram[1788] = 0;
    exp_62_ram[1789] = 1;
    exp_62_ram[1790] = 64;
    exp_62_ram[1791] = 65;
    exp_62_ram[1792] = 0;
    exp_62_ram[1793] = 0;
    exp_62_ram[1794] = 0;
    exp_62_ram[1795] = 0;
    exp_62_ram[1796] = 254;
    exp_62_ram[1797] = 254;
    exp_62_ram[1798] = 0;
    exp_62_ram[1799] = 2;
    exp_62_ram[1800] = 2;
    exp_62_ram[1801] = 2;
    exp_62_ram[1802] = 2;
    exp_62_ram[1803] = 3;
    exp_62_ram[1804] = 0;
    exp_62_ram[1805] = 249;
    exp_62_ram[1806] = 6;
    exp_62_ram[1807] = 6;
    exp_62_ram[1808] = 7;
    exp_62_ram[1809] = 248;
    exp_62_ram[1810] = 0;
    exp_62_ram[1811] = 138;
    exp_62_ram[1812] = 0;
    exp_62_ram[1813] = 0;
    exp_62_ram[1814] = 0;
    exp_62_ram[1815] = 0;
    exp_62_ram[1816] = 1;
    exp_62_ram[1817] = 252;
    exp_62_ram[1818] = 252;
    exp_62_ram[1819] = 252;
    exp_62_ram[1820] = 254;
    exp_62_ram[1821] = 254;
    exp_62_ram[1822] = 1;
    exp_62_ram[1823] = 254;
    exp_62_ram[1824] = 0;
    exp_62_ram[1825] = 140;
    exp_62_ram[1826] = 0;
    exp_62_ram[1827] = 0;
    exp_62_ram[1828] = 0;
    exp_62_ram[1829] = 0;
    exp_62_ram[1830] = 1;
    exp_62_ram[1831] = 1;
    exp_62_ram[1832] = 1;
    exp_62_ram[1833] = 1;
    exp_62_ram[1834] = 2;
    exp_62_ram[1835] = 251;
    exp_62_ram[1836] = 250;
    exp_62_ram[1837] = 251;
    exp_62_ram[1838] = 251;
    exp_62_ram[1839] = 250;
    exp_62_ram[1840] = 252;
    exp_62_ram[1841] = 252;
    exp_62_ram[1842] = 252;
    exp_62_ram[1843] = 252;
    exp_62_ram[1844] = 2;
    exp_62_ram[1845] = 252;
    exp_62_ram[1846] = 254;
    exp_62_ram[1847] = 4;
    exp_62_ram[1848] = 249;
    exp_62_ram[1849] = 1;
    exp_62_ram[1850] = 0;
    exp_62_ram[1851] = 0;
    exp_62_ram[1852] = 0;
    exp_62_ram[1853] = 254;
    exp_62_ram[1854] = 0;
    exp_62_ram[1855] = 255;
    exp_62_ram[1856] = 0;
    exp_62_ram[1857] = 254;
    exp_62_ram[1858] = 0;
    exp_62_ram[1859] = 255;
    exp_62_ram[1860] = 254;
    exp_62_ram[1861] = 0;
    exp_62_ram[1862] = 0;
    exp_62_ram[1863] = 254;
    exp_62_ram[1864] = 0;
    exp_62_ram[1865] = 254;
    exp_62_ram[1866] = 254;
    exp_62_ram[1867] = 0;
    exp_62_ram[1868] = 250;
    exp_62_ram[1869] = 0;
    exp_62_ram[1870] = 255;
    exp_62_ram[1871] = 2;
    exp_62_ram[1872] = 0;
    exp_62_ram[1873] = 254;
    exp_62_ram[1874] = 5;
    exp_62_ram[1875] = 249;
    exp_62_ram[1876] = 1;
    exp_62_ram[1877] = 0;
    exp_62_ram[1878] = 0;
    exp_62_ram[1879] = 0;
    exp_62_ram[1880] = 254;
    exp_62_ram[1881] = 0;
    exp_62_ram[1882] = 254;
    exp_62_ram[1883] = 0;
    exp_62_ram[1884] = 255;
    exp_62_ram[1885] = 0;
    exp_62_ram[1886] = 251;
    exp_62_ram[1887] = 0;
    exp_62_ram[1888] = 255;
    exp_62_ram[1889] = 0;
    exp_62_ram[1890] = 0;
    exp_62_ram[1891] = 254;
    exp_62_ram[1892] = 0;
    exp_62_ram[1893] = 254;
    exp_62_ram[1894] = 254;
    exp_62_ram[1895] = 0;
    exp_62_ram[1896] = 250;
    exp_62_ram[1897] = 0;
    exp_62_ram[1898] = 255;
    exp_62_ram[1899] = 2;
    exp_62_ram[1900] = 0;
    exp_62_ram[1901] = 249;
    exp_62_ram[1902] = 0;
    exp_62_ram[1903] = 0;
    exp_62_ram[1904] = 0;
    exp_62_ram[1905] = 13;
    exp_62_ram[1906] = 0;
    exp_62_ram[1907] = 0;
    exp_62_ram[1908] = 250;
    exp_62_ram[1909] = 250;
    exp_62_ram[1910] = 250;
    exp_62_ram[1911] = 15;
    exp_62_ram[1912] = 3;
    exp_62_ram[1913] = 15;
    exp_62_ram[1914] = 0;
    exp_62_ram[1915] = 255;
    exp_62_ram[1916] = 0;
    exp_62_ram[1917] = 250;
    exp_62_ram[1918] = 15;
    exp_62_ram[1919] = 3;
    exp_62_ram[1920] = 15;
    exp_62_ram[1921] = 0;
    exp_62_ram[1922] = 255;
    exp_62_ram[1923] = 0;
    exp_62_ram[1924] = 0;
    exp_62_ram[1925] = 255;
    exp_62_ram[1926] = 2;
    exp_62_ram[1927] = 0;
    exp_62_ram[1928] = 249;
    exp_62_ram[1929] = 0;
    exp_62_ram[1930] = 0;
    exp_62_ram[1931] = 0;
    exp_62_ram[1932] = 6;
    exp_62_ram[1933] = 0;
    exp_62_ram[1934] = 0;
    exp_62_ram[1935] = 250;
    exp_62_ram[1936] = 250;
    exp_62_ram[1937] = 250;
    exp_62_ram[1938] = 15;
    exp_62_ram[1939] = 3;
    exp_62_ram[1940] = 15;
    exp_62_ram[1941] = 0;
    exp_62_ram[1942] = 255;
    exp_62_ram[1943] = 0;
    exp_62_ram[1944] = 250;
    exp_62_ram[1945] = 15;
    exp_62_ram[1946] = 3;
    exp_62_ram[1947] = 15;
    exp_62_ram[1948] = 0;
    exp_62_ram[1949] = 255;
    exp_62_ram[1950] = 0;
    exp_62_ram[1951] = 0;
    exp_62_ram[1952] = 255;
    exp_62_ram[1953] = 3;
    exp_62_ram[1954] = 0;
    exp_62_ram[1955] = 249;
    exp_62_ram[1956] = 0;
    exp_62_ram[1957] = 0;
    exp_62_ram[1958] = 0;
    exp_62_ram[1959] = 0;
    exp_62_ram[1960] = 0;
    exp_62_ram[1961] = 0;
    exp_62_ram[1962] = 250;
    exp_62_ram[1963] = 250;
    exp_62_ram[1964] = 250;
    exp_62_ram[1965] = 15;
    exp_62_ram[1966] = 3;
    exp_62_ram[1967] = 15;
    exp_62_ram[1968] = 0;
    exp_62_ram[1969] = 255;
    exp_62_ram[1970] = 0;
    exp_62_ram[1971] = 250;
    exp_62_ram[1972] = 15;
    exp_62_ram[1973] = 3;
    exp_62_ram[1974] = 15;
    exp_62_ram[1975] = 0;
    exp_62_ram[1976] = 255;
    exp_62_ram[1977] = 0;
    exp_62_ram[1978] = 0;
    exp_62_ram[1979] = 255;
    exp_62_ram[1980] = 3;
    exp_62_ram[1981] = 0;
    exp_62_ram[1982] = 249;
    exp_62_ram[1983] = 0;
    exp_62_ram[1984] = 0;
    exp_62_ram[1985] = 0;
    exp_62_ram[1986] = 121;
    exp_62_ram[1987] = 0;
    exp_62_ram[1988] = 0;
    exp_62_ram[1989] = 250;
    exp_62_ram[1990] = 250;
    exp_62_ram[1991] = 250;
    exp_62_ram[1992] = 15;
    exp_62_ram[1993] = 3;
    exp_62_ram[1994] = 15;
    exp_62_ram[1995] = 0;
    exp_62_ram[1996] = 255;
    exp_62_ram[1997] = 0;
    exp_62_ram[1998] = 250;
    exp_62_ram[1999] = 15;
    exp_62_ram[2000] = 3;
    exp_62_ram[2001] = 15;
    exp_62_ram[2002] = 0;
    exp_62_ram[2003] = 255;
    exp_62_ram[2004] = 0;
    exp_62_ram[2005] = 0;
    exp_62_ram[2006] = 255;
    exp_62_ram[2007] = 2;
    exp_62_ram[2008] = 0;
    exp_62_ram[2009] = 249;
    exp_62_ram[2010] = 1;
    exp_62_ram[2011] = 118;
    exp_62_ram[2012] = 62;
    exp_62_ram[2013] = 0;
    exp_62_ram[2014] = 114;
    exp_62_ram[2015] = 0;
    exp_62_ram[2016] = 0;
    exp_62_ram[2017] = 250;
    exp_62_ram[2018] = 250;
    exp_62_ram[2019] = 250;
    exp_62_ram[2020] = 15;
    exp_62_ram[2021] = 3;
    exp_62_ram[2022] = 15;
    exp_62_ram[2023] = 0;
    exp_62_ram[2024] = 255;
    exp_62_ram[2025] = 0;
    exp_62_ram[2026] = 250;
    exp_62_ram[2027] = 6;
    exp_62_ram[2028] = 0;
    exp_62_ram[2029] = 110;
    exp_62_ram[2030] = 0;
    exp_62_ram[2031] = 0;
    exp_62_ram[2032] = 250;
    exp_62_ram[2033] = 250;
    exp_62_ram[2034] = 250;
    exp_62_ram[2035] = 15;
    exp_62_ram[2036] = 3;
    exp_62_ram[2037] = 15;
    exp_62_ram[2038] = 0;
    exp_62_ram[2039] = 255;
    exp_62_ram[2040] = 0;
    exp_62_ram[2041] = 250;
    exp_62_ram[2042] = 0;
    exp_62_ram[2043] = 0;
    exp_62_ram[2044] = 106;
    exp_62_ram[2045] = 0;
    exp_62_ram[2046] = 0;
    exp_62_ram[2047] = 250;
    exp_62_ram[2048] = 250;
    exp_62_ram[2049] = 250;
    exp_62_ram[2050] = 15;
    exp_62_ram[2051] = 3;
    exp_62_ram[2052] = 15;
    exp_62_ram[2053] = 0;
    exp_62_ram[2054] = 255;
    exp_62_ram[2055] = 0;
    exp_62_ram[2056] = 250;
    exp_62_ram[2057] = 15;
    exp_62_ram[2058] = 3;
    exp_62_ram[2059] = 15;
    exp_62_ram[2060] = 0;
    exp_62_ram[2061] = 255;
    exp_62_ram[2062] = 0;
    exp_62_ram[2063] = 0;
    exp_62_ram[2064] = 255;
    exp_62_ram[2065] = 0;
    exp_62_ram[2066] = 0;
    exp_62_ram[2067] = 0;
    exp_62_ram[2068] = 255;
    exp_62_ram[2069] = 0;
    exp_62_ram[2070] = 0;
    exp_62_ram[2071] = 255;
    exp_62_ram[2072] = 0;
    exp_62_ram[2073] = 6;
    exp_62_ram[2074] = 6;
    exp_62_ram[2075] = 7;
    exp_62_ram[2076] = 0;
    exp_62_ram[2077] = 254;
    exp_62_ram[2078] = 0;
    exp_62_ram[2079] = 0;
    exp_62_ram[2080] = 2;
    exp_62_ram[2081] = 254;
    exp_62_ram[2082] = 254;
    exp_62_ram[2083] = 55;
    exp_62_ram[2084] = 0;
    exp_62_ram[2085] = 0;
    exp_62_ram[2086] = 185;
    exp_62_ram[2087] = 0;
    exp_62_ram[2088] = 0;
    exp_62_ram[2089] = 1;
    exp_62_ram[2090] = 1;
    exp_62_ram[2091] = 2;
    exp_62_ram[2092] = 0;
    exp_62_ram[2093] = 248;
    exp_62_ram[2094] = 6;
    exp_62_ram[2095] = 6;
    exp_62_ram[2096] = 7;
    exp_62_ram[2097] = 7;
    exp_62_ram[2098] = 7;
    exp_62_ram[2099] = 7;
    exp_62_ram[2100] = 7;
    exp_62_ram[2101] = 7;
    exp_62_ram[2102] = 5;
    exp_62_ram[2103] = 5;
    exp_62_ram[2104] = 8;
    exp_62_ram[2105] = 248;
    exp_62_ram[2106] = 248;
    exp_62_ram[2107] = 248;
    exp_62_ram[2108] = 123;
    exp_62_ram[2109] = 250;
    exp_62_ram[2110] = 0;
    exp_62_ram[2111] = 250;
    exp_62_ram[2112] = 251;
    exp_62_ram[2113] = 0;
    exp_62_ram[2114] = 175;
    exp_62_ram[2115] = 252;
    exp_62_ram[2116] = 252;
    exp_62_ram[2117] = 0;
    exp_62_ram[2118] = 24;
    exp_62_ram[2119] = 2;
    exp_62_ram[2120] = 252;
    exp_62_ram[2121] = 252;
    exp_62_ram[2122] = 0;
    exp_62_ram[2123] = 0;
    exp_62_ram[2124] = 248;
    exp_62_ram[2125] = 0;
    exp_62_ram[2126] = 6;
    exp_62_ram[2127] = 248;
    exp_62_ram[2128] = 0;
    exp_62_ram[2129] = 0;
    exp_62_ram[2130] = 248;
    exp_62_ram[2131] = 0;
    exp_62_ram[2132] = 4;
    exp_62_ram[2133] = 251;
    exp_62_ram[2134] = 0;
    exp_62_ram[2135] = 250;
    exp_62_ram[2136] = 251;
    exp_62_ram[2137] = 0;
    exp_62_ram[2138] = 252;
    exp_62_ram[2139] = 0;
    exp_62_ram[2140] = 250;
    exp_62_ram[2141] = 252;
    exp_62_ram[2142] = 0;
    exp_62_ram[2143] = 0;
    exp_62_ram[2144] = 248;
    exp_62_ram[2145] = 248;
    exp_62_ram[2146] = 65;
    exp_62_ram[2147] = 0;
    exp_62_ram[2148] = 0;
    exp_62_ram[2149] = 65;
    exp_62_ram[2150] = 64;
    exp_62_ram[2151] = 0;
    exp_62_ram[2152] = 248;
    exp_62_ram[2153] = 248;
    exp_62_ram[2154] = 245;
    exp_62_ram[2155] = 0;
    exp_62_ram[2156] = 250;
    exp_62_ram[2157] = 252;
    exp_62_ram[2158] = 251;
    exp_62_ram[2159] = 0;
    exp_62_ram[2160] = 251;
    exp_62_ram[2161] = 0;
    exp_62_ram[2162] = 0;
    exp_62_ram[2163] = 167;
    exp_62_ram[2164] = 252;
    exp_62_ram[2165] = 252;
    exp_62_ram[2166] = 0;
    exp_62_ram[2167] = 24;
    exp_62_ram[2168] = 2;
    exp_62_ram[2169] = 252;
    exp_62_ram[2170] = 252;
    exp_62_ram[2171] = 0;
    exp_62_ram[2172] = 0;
    exp_62_ram[2173] = 248;
    exp_62_ram[2174] = 0;
    exp_62_ram[2175] = 8;
    exp_62_ram[2176] = 248;
    exp_62_ram[2177] = 0;
    exp_62_ram[2178] = 0;
    exp_62_ram[2179] = 248;
    exp_62_ram[2180] = 0;
    exp_62_ram[2181] = 6;
    exp_62_ram[2182] = 251;
    exp_62_ram[2183] = 0;
    exp_62_ram[2184] = 250;
    exp_62_ram[2185] = 251;
    exp_62_ram[2186] = 0;
    exp_62_ram[2187] = 252;
    exp_62_ram[2188] = 0;
    exp_62_ram[2189] = 250;
    exp_62_ram[2190] = 252;
    exp_62_ram[2191] = 0;
    exp_62_ram[2192] = 252;
    exp_62_ram[2193] = 0;
    exp_62_ram[2194] = 252;
    exp_62_ram[2195] = 252;
    exp_62_ram[2196] = 0;
    exp_62_ram[2197] = 0;
    exp_62_ram[2198] = 248;
    exp_62_ram[2199] = 248;
    exp_62_ram[2200] = 65;
    exp_62_ram[2201] = 0;
    exp_62_ram[2202] = 0;
    exp_62_ram[2203] = 65;
    exp_62_ram[2204] = 64;
    exp_62_ram[2205] = 0;
    exp_62_ram[2206] = 248;
    exp_62_ram[2207] = 248;
    exp_62_ram[2208] = 243;
    exp_62_ram[2209] = 0;
    exp_62_ram[2210] = 251;
    exp_62_ram[2211] = 137;
    exp_62_ram[2212] = 250;
    exp_62_ram[2213] = 248;
    exp_62_ram[2214] = 0;
    exp_62_ram[2215] = 24;
    exp_62_ram[2216] = 0;
    exp_62_ram[2217] = 63;
    exp_62_ram[2218] = 0;
    exp_62_ram[2219] = 0;
    exp_62_ram[2220] = 248;
    exp_62_ram[2221] = 250;
    exp_62_ram[2222] = 249;
    exp_62_ram[2223] = 0;
    exp_62_ram[2224] = 250;
    exp_62_ram[2225] = 251;
    exp_62_ram[2226] = 249;
    exp_62_ram[2227] = 0;
    exp_62_ram[2228] = 250;
    exp_62_ram[2229] = 251;
    exp_62_ram[2230] = 0;
    exp_62_ram[2231] = 2;
    exp_62_ram[2232] = 250;
    exp_62_ram[2233] = 252;
    exp_62_ram[2234] = 249;
    exp_62_ram[2235] = 0;
    exp_62_ram[2236] = 252;
    exp_62_ram[2237] = 250;
    exp_62_ram[2238] = 248;
    exp_62_ram[2239] = 65;
    exp_62_ram[2240] = 248;
    exp_62_ram[2241] = 248;
    exp_62_ram[2242] = 0;
    exp_62_ram[2243] = 225;
    exp_62_ram[2244] = 0;
    exp_62_ram[2245] = 56;
    exp_62_ram[2246] = 0;
    exp_62_ram[2247] = 0;
    exp_62_ram[2248] = 248;
    exp_62_ram[2249] = 250;
    exp_62_ram[2250] = 249;
    exp_62_ram[2251] = 250;
    exp_62_ram[2252] = 250;
    exp_62_ram[2253] = 248;
    exp_62_ram[2254] = 65;
    exp_62_ram[2255] = 248;
    exp_62_ram[2256] = 248;
    exp_62_ram[2257] = 3;
    exp_62_ram[2258] = 0;
    exp_62_ram[2259] = 53;
    exp_62_ram[2260] = 0;
    exp_62_ram[2261] = 0;
    exp_62_ram[2262] = 248;
    exp_62_ram[2263] = 250;
    exp_62_ram[2264] = 249;
    exp_62_ram[2265] = 250;
    exp_62_ram[2266] = 250;
    exp_62_ram[2267] = 248;
    exp_62_ram[2268] = 65;
    exp_62_ram[2269] = 248;
    exp_62_ram[2270] = 248;
    exp_62_ram[2271] = 250;
    exp_62_ram[2272] = 248;
    exp_62_ram[2273] = 250;
    exp_62_ram[2274] = 250;
    exp_62_ram[2275] = 250;
    exp_62_ram[2276] = 251;
    exp_62_ram[2277] = 251;
    exp_62_ram[2278] = 251;
    exp_62_ram[2279] = 251;
    exp_62_ram[2280] = 252;
    exp_62_ram[2281] = 252;
    exp_62_ram[2282] = 1;
    exp_62_ram[2283] = 0;
    exp_62_ram[2284] = 1;
    exp_62_ram[2285] = 1;
    exp_62_ram[2286] = 0;
    exp_62_ram[2287] = 0;
    exp_62_ram[2288] = 0;
    exp_62_ram[2289] = 0;
    exp_62_ram[2290] = 2;
    exp_62_ram[2291] = 248;
    exp_62_ram[2292] = 7;
    exp_62_ram[2293] = 7;
    exp_62_ram[2294] = 7;
    exp_62_ram[2295] = 7;
    exp_62_ram[2296] = 6;
    exp_62_ram[2297] = 6;
    exp_62_ram[2298] = 6;
    exp_62_ram[2299] = 6;
    exp_62_ram[2300] = 5;
    exp_62_ram[2301] = 5;
    exp_62_ram[2302] = 8;
    exp_62_ram[2303] = 0;
    exp_62_ram[2304] = 246;
    exp_62_ram[2305] = 8;
    exp_62_ram[2306] = 8;
    exp_62_ram[2307] = 8;
    exp_62_ram[2308] = 9;
    exp_62_ram[2309] = 9;
    exp_62_ram[2310] = 10;
    exp_62_ram[2311] = 248;
    exp_62_ram[2312] = 0;
    exp_62_ram[2313] = 0;
    exp_62_ram[2314] = 252;
    exp_62_ram[2315] = 253;
    exp_62_ram[2316] = 249;
    exp_62_ram[2317] = 0;
    exp_62_ram[2318] = 0;
    exp_62_ram[2319] = 252;
    exp_62_ram[2320] = 252;
    exp_62_ram[2321] = 253;
    exp_62_ram[2322] = 253;
    exp_62_ram[2323] = 220;
    exp_62_ram[2324] = 0;
    exp_62_ram[2325] = 0;
    exp_62_ram[2326] = 0;
    exp_62_ram[2327] = 225;
    exp_62_ram[2328] = 0;
    exp_62_ram[2329] = 252;
    exp_62_ram[2330] = 252;
    exp_62_ram[2331] = 0;
    exp_62_ram[2332] = 254;
    exp_62_ram[2333] = 0;
    exp_62_ram[2334] = 65;
    exp_62_ram[2335] = 0;
    exp_62_ram[2336] = 253;
    exp_62_ram[2337] = 253;
    exp_62_ram[2338] = 0;
    exp_62_ram[2339] = 0;
    exp_62_ram[2340] = 1;
    exp_62_ram[2341] = 0;
    exp_62_ram[2342] = 0;
    exp_62_ram[2343] = 0;
    exp_62_ram[2344] = 0;
    exp_62_ram[2345] = 0;
    exp_62_ram[2346] = 253;
    exp_62_ram[2347] = 253;
    exp_62_ram[2348] = 0;
    exp_62_ram[2349] = 0;
    exp_62_ram[2350] = 0;
    exp_62_ram[2351] = 0;
    exp_62_ram[2352] = 0;
    exp_62_ram[2353] = 0;
    exp_62_ram[2354] = 252;
    exp_62_ram[2355] = 252;
    exp_62_ram[2356] = 0;
    exp_62_ram[2357] = 0;
    exp_62_ram[2358] = 246;
    exp_62_ram[2359] = 252;
    exp_62_ram[2360] = 252;
    exp_62_ram[2361] = 0;
    exp_62_ram[2362] = 188;
    exp_62_ram[2363] = 246;
    exp_62_ram[2364] = 246;
    exp_62_ram[2365] = 246;
    exp_62_ram[2366] = 246;
    exp_62_ram[2367] = 247;
    exp_62_ram[2368] = 247;
    exp_62_ram[2369] = 247;
    exp_62_ram[2370] = 247;
    exp_62_ram[2371] = 248;
    exp_62_ram[2372] = 0;
    exp_62_ram[2373] = 1;
    exp_62_ram[2374] = 1;
    exp_62_ram[2375] = 0;
    exp_62_ram[2376] = 0;
    exp_62_ram[2377] = 0;
    exp_62_ram[2378] = 0;
    exp_62_ram[2379] = 0;
    exp_62_ram[2380] = 2;
    exp_62_ram[2381] = 253;
    exp_62_ram[2382] = 253;
    exp_62_ram[2383] = 205;
    exp_62_ram[2384] = 0;
    exp_62_ram[2385] = 0;
    exp_62_ram[2386] = 0;
    exp_62_ram[2387] = 2;
    exp_62_ram[2388] = 0;
    exp_62_ram[2389] = 0;
    exp_62_ram[2390] = 0;
    exp_62_ram[2391] = 9;
    exp_62_ram[2392] = 9;
    exp_62_ram[2393] = 9;
    exp_62_ram[2394] = 9;
    exp_62_ram[2395] = 8;
    exp_62_ram[2396] = 10;
    exp_62_ram[2397] = 0;
    exp_62_ram[2398] = 253;
    exp_62_ram[2399] = 2;
    exp_62_ram[2400] = 2;
    exp_62_ram[2401] = 3;
    exp_62_ram[2402] = 252;
    exp_62_ram[2403] = 254;
    exp_62_ram[2404] = 253;
    exp_62_ram[2405] = 240;
    exp_62_ram[2406] = 0;
    exp_62_ram[2407] = 254;
    exp_62_ram[2408] = 254;
    exp_62_ram[2409] = 253;
    exp_62_ram[2410] = 0;
    exp_62_ram[2411] = 2;
    exp_62_ram[2412] = 254;
    exp_62_ram[2413] = 0;
    exp_62_ram[2414] = 0;
    exp_62_ram[2415] = 0;
    exp_62_ram[2416] = 0;
    exp_62_ram[2417] = 254;
    exp_62_ram[2418] = 254;
    exp_62_ram[2419] = 254;
    exp_62_ram[2420] = 0;
    exp_62_ram[2421] = 253;
    exp_62_ram[2422] = 254;
    exp_62_ram[2423] = 251;
    exp_62_ram[2424] = 0;
    exp_62_ram[2425] = 254;
    exp_62_ram[2426] = 0;
    exp_62_ram[2427] = 2;
    exp_62_ram[2428] = 2;
    exp_62_ram[2429] = 3;
    exp_62_ram[2430] = 0;
    exp_62_ram[2431] = 255;
    exp_62_ram[2432] = 0;
    exp_62_ram[2433] = 0;
    exp_62_ram[2434] = 1;
    exp_62_ram[2435] = 0;
    exp_62_ram[2436] = 237;
    exp_62_ram[2437] = 0;
    exp_62_ram[2438] = 246;
    exp_62_ram[2439] = 0;
    exp_62_ram[2440] = 0;
    exp_62_ram[2441] = 0;
    exp_62_ram[2442] = 0;
    exp_62_ram[2443] = 1;
    exp_62_ram[2444] = 0;
    exp_62_ram[2445] = 253;
    exp_62_ram[2446] = 2;
    exp_62_ram[2447] = 2;
    exp_62_ram[2448] = 3;
    exp_62_ram[2449] = 252;
    exp_62_ram[2450] = 252;
    exp_62_ram[2451] = 252;
    exp_62_ram[2452] = 59;
    exp_62_ram[2453] = 160;
    exp_62_ram[2454] = 254;
    exp_62_ram[2455] = 0;
    exp_62_ram[2456] = 254;
    exp_62_ram[2457] = 254;
    exp_62_ram[2458] = 9;
    exp_62_ram[2459] = 253;
    exp_62_ram[2460] = 254;
    exp_62_ram[2461] = 2;
    exp_62_ram[2462] = 254;
    exp_62_ram[2463] = 254;
    exp_62_ram[2464] = 0;
    exp_62_ram[2465] = 254;
    exp_62_ram[2466] = 0;
    exp_62_ram[2467] = 254;
    exp_62_ram[2468] = 0;
    exp_62_ram[2469] = 2;
    exp_62_ram[2470] = 254;
    exp_62_ram[2471] = 3;
    exp_62_ram[2472] = 253;
    exp_62_ram[2473] = 0;
    exp_62_ram[2474] = 225;
    exp_62_ram[2475] = 0;
    exp_62_ram[2476] = 254;
    exp_62_ram[2477] = 2;
    exp_62_ram[2478] = 254;
    exp_62_ram[2479] = 253;
    exp_62_ram[2480] = 0;
    exp_62_ram[2481] = 254;
    exp_62_ram[2482] = 3;
    exp_62_ram[2483] = 253;
    exp_62_ram[2484] = 0;
    exp_62_ram[2485] = 223;
    exp_62_ram[2486] = 253;
    exp_62_ram[2487] = 254;
    exp_62_ram[2488] = 2;
    exp_62_ram[2489] = 252;
    exp_62_ram[2490] = 254;
    exp_62_ram[2491] = 0;
    exp_62_ram[2492] = 2;
    exp_62_ram[2493] = 254;
    exp_62_ram[2494] = 254;
    exp_62_ram[2495] = 255;
    exp_62_ram[2496] = 254;
    exp_62_ram[2497] = 254;
    exp_62_ram[2498] = 246;
    exp_62_ram[2499] = 0;
    exp_62_ram[2500] = 0;
    exp_62_ram[2501] = 2;
    exp_62_ram[2502] = 2;
    exp_62_ram[2503] = 3;
    exp_62_ram[2504] = 0;
    exp_62_ram[2505] = 254;
    exp_62_ram[2506] = 0;
    exp_62_ram[2507] = 0;
    exp_62_ram[2508] = 2;
    exp_62_ram[2509] = 254;
    exp_62_ram[2510] = 254;
    exp_62_ram[2511] = 254;
    exp_62_ram[2512] = 254;
    exp_62_ram[2513] = 0;
    exp_62_ram[2514] = 238;
    exp_62_ram[2515] = 0;
    exp_62_ram[2516] = 0;
    exp_62_ram[2517] = 0;
    exp_62_ram[2518] = 237;
    exp_62_ram[2519] = 0;
    exp_62_ram[2520] = 1;
    exp_62_ram[2521] = 1;
    exp_62_ram[2522] = 2;
    exp_62_ram[2523] = 0;
    exp_62_ram[2524] = 253;
    exp_62_ram[2525] = 2;
    exp_62_ram[2526] = 2;
    exp_62_ram[2527] = 3;
    exp_62_ram[2528] = 3;
    exp_62_ram[2529] = 3;
    exp_62_ram[2530] = 252;
    exp_62_ram[2531] = 178;
    exp_62_ram[2532] = 254;
    exp_62_ram[2533] = 254;
    exp_62_ram[2534] = 0;
    exp_62_ram[2535] = 177;
    exp_62_ram[2536] = 0;
    exp_62_ram[2537] = 0;
    exp_62_ram[2538] = 254;
    exp_62_ram[2539] = 254;
    exp_62_ram[2540] = 64;
    exp_62_ram[2541] = 0;
    exp_62_ram[2542] = 1;
    exp_62_ram[2543] = 64;
    exp_62_ram[2544] = 65;
    exp_62_ram[2545] = 0;
    exp_62_ram[2546] = 253;
    exp_62_ram[2547] = 0;
    exp_62_ram[2548] = 0;
    exp_62_ram[2549] = 0;
    exp_62_ram[2550] = 0;
    exp_62_ram[2551] = 252;
    exp_62_ram[2552] = 0;
    exp_62_ram[2553] = 0;
    exp_62_ram[2554] = 0;
    exp_62_ram[2555] = 0;
    exp_62_ram[2556] = 0;
    exp_62_ram[2557] = 250;
    exp_62_ram[2558] = 0;
    exp_62_ram[2559] = 0;
    exp_62_ram[2560] = 2;
    exp_62_ram[2561] = 2;
    exp_62_ram[2562] = 2;
    exp_62_ram[2563] = 2;
    exp_62_ram[2564] = 3;
    exp_62_ram[2565] = 0;
    exp_62_ram[2566] = 255;
    exp_62_ram[2567] = 0;
    exp_62_ram[2568] = 0;
    exp_62_ram[2569] = 1;
    exp_62_ram[2570] = 0;
    exp_62_ram[2571] = 142;
    exp_62_ram[2572] = 219;
    exp_62_ram[2573] = 0;
    exp_62_ram[2574] = 0;
    exp_62_ram[2575] = 0;
    exp_62_ram[2576] = 1;
    exp_62_ram[2577] = 0;
    exp_62_ram[2578] = 254;
    exp_62_ram[2579] = 0;
    exp_62_ram[2580] = 0;
    exp_62_ram[2581] = 2;
    exp_62_ram[2582] = 0;
    exp_62_ram[2583] = 143;
    exp_62_ram[2584] = 216;
    exp_62_ram[2585] = 0;
    exp_62_ram[2586] = 254;
    exp_62_ram[2587] = 254;
    exp_62_ram[2588] = 11;
    exp_62_ram[2589] = 0;
    exp_62_ram[2590] = 254;
    exp_62_ram[2591] = 234;
    exp_62_ram[2592] = 0;
    exp_62_ram[2593] = 199;
    exp_62_ram[2594] = 3;
    exp_62_ram[2595] = 254;
    exp_62_ram[2596] = 0;
    exp_62_ram[2597] = 254;
    exp_62_ram[2598] = 0;
    exp_62_ram[2599] = 238;
    exp_62_ram[2600] = 0;
    exp_62_ram[2601] = 254;
    exp_62_ram[2602] = 193;
    exp_62_ram[2603] = 0;
    exp_62_ram[2604] = 237;
    exp_62_ram[2605] = 0;
    exp_62_ram[2606] = 2;
    exp_62_ram[2607] = 0;
    exp_62_ram[2608] = 235;
    exp_62_ram[2609] = 254;
    exp_62_ram[2610] = 7;
    exp_62_ram[2611] = 252;
    exp_62_ram[2612] = 3;
    exp_62_ram[2613] = 254;
    exp_62_ram[2614] = 64;
    exp_62_ram[2615] = 254;
    exp_62_ram[2616] = 0;
    exp_62_ram[2617] = 238;
    exp_62_ram[2618] = 0;
    exp_62_ram[2619] = 254;
    exp_62_ram[2620] = 189;
    exp_62_ram[2621] = 0;
    exp_62_ram[2622] = 237;
    exp_62_ram[2623] = 0;
    exp_62_ram[2624] = 2;
    exp_62_ram[2625] = 0;
    exp_62_ram[2626] = 230;
    exp_62_ram[2627] = 254;
    exp_62_ram[2628] = 0;
    exp_62_ram[2629] = 252;
    exp_62_ram[2630] = 254;
    exp_62_ram[2631] = 0;
    exp_62_ram[2632] = 254;
    exp_62_ram[2633] = 254;
    exp_62_ram[2634] = 0;
    exp_62_ram[2635] = 244;
    exp_62_ram[2636] = 0;
    exp_62_ram[2637] = 238;
    exp_62_ram[2638] = 0;
    exp_62_ram[2639] = 0;
    exp_62_ram[2640] = 184;
    exp_62_ram[2641] = 0;
    exp_62_ram[2642] = 1;
    exp_62_ram[2643] = 1;
    exp_62_ram[2644] = 2;
    exp_62_ram[2645] = 0;
    exp_62_ram[2646] = 254;
    exp_62_ram[2647] = 0;
    exp_62_ram[2648] = 0;
    exp_62_ram[2649] = 2;
    exp_62_ram[2650] = 0;
    exp_62_ram[2651] = 145;
    exp_62_ram[2652] = 199;
    exp_62_ram[2653] = 254;
    exp_62_ram[2654] = 11;
    exp_62_ram[2655] = 0;
    exp_62_ram[2656] = 254;
    exp_62_ram[2657] = 218;
    exp_62_ram[2658] = 0;
    exp_62_ram[2659] = 183;
    exp_62_ram[2660] = 254;
    exp_62_ram[2661] = 3;
    exp_62_ram[2662] = 0;
    exp_62_ram[2663] = 238;
    exp_62_ram[2664] = 0;
    exp_62_ram[2665] = 254;
    exp_62_ram[2666] = 177;
    exp_62_ram[2667] = 0;
    exp_62_ram[2668] = 237;
    exp_62_ram[2669] = 62;
    exp_62_ram[2670] = 2;
    exp_62_ram[2671] = 0;
    exp_62_ram[2672] = 219;
    exp_62_ram[2673] = 254;
    exp_62_ram[2674] = 0;
    exp_62_ram[2675] = 254;
    exp_62_ram[2676] = 254;
    exp_62_ram[2677] = 63;
    exp_62_ram[2678] = 252;
    exp_62_ram[2679] = 63;
    exp_62_ram[2680] = 254;
    exp_62_ram[2681] = 3;
    exp_62_ram[2682] = 0;
    exp_62_ram[2683] = 238;
    exp_62_ram[2684] = 0;
    exp_62_ram[2685] = 254;
    exp_62_ram[2686] = 172;
    exp_62_ram[2687] = 0;
    exp_62_ram[2688] = 237;
    exp_62_ram[2689] = 62;
    exp_62_ram[2690] = 2;
    exp_62_ram[2691] = 0;
    exp_62_ram[2692] = 214;
    exp_62_ram[2693] = 254;
    exp_62_ram[2694] = 255;
    exp_62_ram[2695] = 254;
    exp_62_ram[2696] = 254;
    exp_62_ram[2697] = 252;
    exp_62_ram[2698] = 254;
    exp_62_ram[2699] = 0;
    exp_62_ram[2700] = 254;
    exp_62_ram[2701] = 254;
    exp_62_ram[2702] = 0;
    exp_62_ram[2703] = 244;
    exp_62_ram[2704] = 0;
    exp_62_ram[2705] = 238;
    exp_62_ram[2706] = 0;
    exp_62_ram[2707] = 0;
    exp_62_ram[2708] = 167;
    exp_62_ram[2709] = 0;
    exp_62_ram[2710] = 1;
    exp_62_ram[2711] = 1;
    exp_62_ram[2712] = 2;
    exp_62_ram[2713] = 0;
    exp_62_ram[2714] = 249;
    exp_62_ram[2715] = 6;
    exp_62_ram[2716] = 6;
    exp_62_ram[2717] = 7;
    exp_62_ram[2718] = 7;
    exp_62_ram[2719] = 5;
    exp_62_ram[2720] = 5;
    exp_62_ram[2721] = 5;
    exp_62_ram[2722] = 5;
    exp_62_ram[2723] = 5;
    exp_62_ram[2724] = 5;
    exp_62_ram[2725] = 5;
    exp_62_ram[2726] = 5;
    exp_62_ram[2727] = 7;
    exp_62_ram[2728] = 0;
    exp_62_ram[2729] = 250;
    exp_62_ram[2730] = 0;
    exp_62_ram[2731] = 0;
    exp_62_ram[2732] = 250;
    exp_62_ram[2733] = 250;
    exp_62_ram[2734] = 255;
    exp_62_ram[2735] = 252;
    exp_62_ram[2736] = 252;
    exp_62_ram[2737] = 252;
    exp_62_ram[2738] = 6;
    exp_62_ram[2739] = 251;
    exp_62_ram[2740] = 18;
    exp_62_ram[2741] = 103;
    exp_62_ram[2742] = 2;
    exp_62_ram[2743] = 250;
    exp_62_ram[2744] = 251;
    exp_62_ram[2745] = 18;
    exp_62_ram[2746] = 103;
    exp_62_ram[2747] = 2;
    exp_62_ram[2748] = 250;
    exp_62_ram[2749] = 251;
    exp_62_ram[2750] = 18;
    exp_62_ram[2751] = 103;
    exp_62_ram[2752] = 2;
    exp_62_ram[2753] = 250;
    exp_62_ram[2754] = 251;
    exp_62_ram[2755] = 18;
    exp_62_ram[2756] = 103;
    exp_62_ram[2757] = 2;
    exp_62_ram[2758] = 250;
    exp_62_ram[2759] = 252;
    exp_62_ram[2760] = 0;
    exp_62_ram[2761] = 252;
    exp_62_ram[2762] = 248;
    exp_62_ram[2763] = 0;
    exp_62_ram[2764] = 0;
    exp_62_ram[2765] = 252;
    exp_62_ram[2766] = 252;
    exp_62_ram[2767] = 64;
    exp_62_ram[2768] = 0;
    exp_62_ram[2769] = 1;
    exp_62_ram[2770] = 64;
    exp_62_ram[2771] = 65;
    exp_62_ram[2772] = 0;
    exp_62_ram[2773] = 0;
    exp_62_ram[2774] = 237;
    exp_62_ram[2775] = 250;
    exp_62_ram[2776] = 250;
    exp_62_ram[2777] = 250;
    exp_62_ram[2778] = 250;
    exp_62_ram[2779] = 0;
    exp_62_ram[2780] = 0;
    exp_62_ram[2781] = 244;
    exp_62_ram[2782] = 0;
    exp_62_ram[2783] = 0;
    exp_62_ram[2784] = 0;
    exp_62_ram[2785] = 0;
    exp_62_ram[2786] = 0;
    exp_62_ram[2787] = 244;
    exp_62_ram[2788] = 252;
    exp_62_ram[2789] = 0;
    exp_62_ram[2790] = 0;
    exp_62_ram[2791] = 184;
    exp_62_ram[2792] = 0;
    exp_62_ram[2793] = 146;
    exp_62_ram[2794] = 164;
    exp_62_ram[2795] = 240;
    exp_62_ram[2796] = 252;
    exp_62_ram[2797] = 252;
    exp_62_ram[2798] = 252;
    exp_62_ram[2799] = 18;
    exp_62_ram[2800] = 251;
    exp_62_ram[2801] = 251;
    exp_62_ram[2802] = 18;
    exp_62_ram[2803] = 103;
    exp_62_ram[2804] = 2;
    exp_62_ram[2805] = 0;
    exp_62_ram[2806] = 2;
    exp_62_ram[2807] = 0;
    exp_62_ram[2808] = 18;
    exp_62_ram[2809] = 103;
    exp_62_ram[2810] = 2;
    exp_62_ram[2811] = 2;
    exp_62_ram[2812] = 0;
    exp_62_ram[2813] = 1;
    exp_62_ram[2814] = 0;
    exp_62_ram[2815] = 251;
    exp_62_ram[2816] = 251;
    exp_62_ram[2817] = 251;
    exp_62_ram[2818] = 251;
    exp_62_ram[2819] = 18;
    exp_62_ram[2820] = 103;
    exp_62_ram[2821] = 2;
    exp_62_ram[2822] = 0;
    exp_62_ram[2823] = 2;
    exp_62_ram[2824] = 0;
    exp_62_ram[2825] = 18;
    exp_62_ram[2826] = 103;
    exp_62_ram[2827] = 2;
    exp_62_ram[2828] = 2;
    exp_62_ram[2829] = 0;
    exp_62_ram[2830] = 1;
    exp_62_ram[2831] = 0;
    exp_62_ram[2832] = 251;
    exp_62_ram[2833] = 251;
    exp_62_ram[2834] = 251;
    exp_62_ram[2835] = 251;
    exp_62_ram[2836] = 18;
    exp_62_ram[2837] = 103;
    exp_62_ram[2838] = 2;
    exp_62_ram[2839] = 0;
    exp_62_ram[2840] = 2;
    exp_62_ram[2841] = 0;
    exp_62_ram[2842] = 18;
    exp_62_ram[2843] = 103;
    exp_62_ram[2844] = 2;
    exp_62_ram[2845] = 2;
    exp_62_ram[2846] = 0;
    exp_62_ram[2847] = 1;
    exp_62_ram[2848] = 0;
    exp_62_ram[2849] = 251;
    exp_62_ram[2850] = 251;
    exp_62_ram[2851] = 251;
    exp_62_ram[2852] = 251;
    exp_62_ram[2853] = 18;
    exp_62_ram[2854] = 103;
    exp_62_ram[2855] = 2;
    exp_62_ram[2856] = 0;
    exp_62_ram[2857] = 2;
    exp_62_ram[2858] = 0;
    exp_62_ram[2859] = 18;
    exp_62_ram[2860] = 103;
    exp_62_ram[2861] = 2;
    exp_62_ram[2862] = 2;
    exp_62_ram[2863] = 0;
    exp_62_ram[2864] = 1;
    exp_62_ram[2865] = 0;
    exp_62_ram[2866] = 251;
    exp_62_ram[2867] = 251;
    exp_62_ram[2868] = 252;
    exp_62_ram[2869] = 0;
    exp_62_ram[2870] = 252;
    exp_62_ram[2871] = 221;
    exp_62_ram[2872] = 0;
    exp_62_ram[2873] = 0;
    exp_62_ram[2874] = 252;
    exp_62_ram[2875] = 252;
    exp_62_ram[2876] = 64;
    exp_62_ram[2877] = 0;
    exp_62_ram[2878] = 1;
    exp_62_ram[2879] = 64;
    exp_62_ram[2880] = 65;
    exp_62_ram[2881] = 0;
    exp_62_ram[2882] = 0;
    exp_62_ram[2883] = 237;
    exp_62_ram[2884] = 250;
    exp_62_ram[2885] = 250;
    exp_62_ram[2886] = 250;
    exp_62_ram[2887] = 250;
    exp_62_ram[2888] = 0;
    exp_62_ram[2889] = 0;
    exp_62_ram[2890] = 232;
    exp_62_ram[2891] = 0;
    exp_62_ram[2892] = 0;
    exp_62_ram[2893] = 0;
    exp_62_ram[2894] = 0;
    exp_62_ram[2895] = 0;
    exp_62_ram[2896] = 232;
    exp_62_ram[2897] = 252;
    exp_62_ram[2898] = 0;
    exp_62_ram[2899] = 0;
    exp_62_ram[2900] = 157;
    exp_62_ram[2901] = 0;
    exp_62_ram[2902] = 149;
    exp_62_ram[2903] = 136;
    exp_62_ram[2904] = 212;
    exp_62_ram[2905] = 252;
    exp_62_ram[2906] = 252;
    exp_62_ram[2907] = 252;
    exp_62_ram[2908] = 6;
    exp_62_ram[2909] = 251;
    exp_62_ram[2910] = 18;
    exp_62_ram[2911] = 103;
    exp_62_ram[2912] = 2;
    exp_62_ram[2913] = 250;
    exp_62_ram[2914] = 251;
    exp_62_ram[2915] = 18;
    exp_62_ram[2916] = 103;
    exp_62_ram[2917] = 2;
    exp_62_ram[2918] = 250;
    exp_62_ram[2919] = 251;
    exp_62_ram[2920] = 18;
    exp_62_ram[2921] = 103;
    exp_62_ram[2922] = 2;
    exp_62_ram[2923] = 250;
    exp_62_ram[2924] = 251;
    exp_62_ram[2925] = 18;
    exp_62_ram[2926] = 103;
    exp_62_ram[2927] = 2;
    exp_62_ram[2928] = 250;
    exp_62_ram[2929] = 252;
    exp_62_ram[2930] = 0;
    exp_62_ram[2931] = 252;
    exp_62_ram[2932] = 205;
    exp_62_ram[2933] = 0;
    exp_62_ram[2934] = 0;
    exp_62_ram[2935] = 252;
    exp_62_ram[2936] = 252;
    exp_62_ram[2937] = 64;
    exp_62_ram[2938] = 0;
    exp_62_ram[2939] = 1;
    exp_62_ram[2940] = 64;
    exp_62_ram[2941] = 65;
    exp_62_ram[2942] = 0;
    exp_62_ram[2943] = 0;
    exp_62_ram[2944] = 237;
    exp_62_ram[2945] = 248;
    exp_62_ram[2946] = 248;
    exp_62_ram[2947] = 249;
    exp_62_ram[2948] = 249;
    exp_62_ram[2949] = 0;
    exp_62_ram[2950] = 0;
    exp_62_ram[2951] = 244;
    exp_62_ram[2952] = 0;
    exp_62_ram[2953] = 0;
    exp_62_ram[2954] = 0;
    exp_62_ram[2955] = 0;
    exp_62_ram[2956] = 0;
    exp_62_ram[2957] = 244;
    exp_62_ram[2958] = 252;
    exp_62_ram[2959] = 0;
    exp_62_ram[2960] = 0;
    exp_62_ram[2961] = 142;
    exp_62_ram[2962] = 0;
    exp_62_ram[2963] = 151;
    exp_62_ram[2964] = 249;
    exp_62_ram[2965] = 197;
    exp_62_ram[2966] = 252;
    exp_62_ram[2967] = 252;
    exp_62_ram[2968] = 252;
    exp_62_ram[2969] = 13;
    exp_62_ram[2970] = 251;
    exp_62_ram[2971] = 251;
    exp_62_ram[2972] = 18;
    exp_62_ram[2973] = 103;
    exp_62_ram[2974] = 0;
    exp_62_ram[2975] = 0;
    exp_62_ram[2976] = 0;
    exp_62_ram[2977] = 160;
    exp_62_ram[2978] = 0;
    exp_62_ram[2979] = 0;
    exp_62_ram[2980] = 250;
    exp_62_ram[2981] = 250;
    exp_62_ram[2982] = 251;
    exp_62_ram[2983] = 251;
    exp_62_ram[2984] = 18;
    exp_62_ram[2985] = 103;
    exp_62_ram[2986] = 0;
    exp_62_ram[2987] = 0;
    exp_62_ram[2988] = 0;
    exp_62_ram[2989] = 157;
    exp_62_ram[2990] = 0;
    exp_62_ram[2991] = 0;
    exp_62_ram[2992] = 250;
    exp_62_ram[2993] = 250;
    exp_62_ram[2994] = 251;
    exp_62_ram[2995] = 251;
    exp_62_ram[2996] = 18;
    exp_62_ram[2997] = 103;
    exp_62_ram[2998] = 0;
    exp_62_ram[2999] = 0;
    exp_62_ram[3000] = 0;
    exp_62_ram[3001] = 154;
    exp_62_ram[3002] = 0;
    exp_62_ram[3003] = 0;
    exp_62_ram[3004] = 250;
    exp_62_ram[3005] = 250;
    exp_62_ram[3006] = 251;
    exp_62_ram[3007] = 251;
    exp_62_ram[3008] = 18;
    exp_62_ram[3009] = 103;
    exp_62_ram[3010] = 0;
    exp_62_ram[3011] = 0;
    exp_62_ram[3012] = 0;
    exp_62_ram[3013] = 151;
    exp_62_ram[3014] = 0;
    exp_62_ram[3015] = 0;
    exp_62_ram[3016] = 250;
    exp_62_ram[3017] = 250;
    exp_62_ram[3018] = 252;
    exp_62_ram[3019] = 0;
    exp_62_ram[3020] = 252;
    exp_62_ram[3021] = 183;
    exp_62_ram[3022] = 0;
    exp_62_ram[3023] = 0;
    exp_62_ram[3024] = 252;
    exp_62_ram[3025] = 252;
    exp_62_ram[3026] = 64;
    exp_62_ram[3027] = 0;
    exp_62_ram[3028] = 1;
    exp_62_ram[3029] = 64;
    exp_62_ram[3030] = 65;
    exp_62_ram[3031] = 0;
    exp_62_ram[3032] = 0;
    exp_62_ram[3033] = 237;
    exp_62_ram[3034] = 0;
    exp_62_ram[3035] = 0;
    exp_62_ram[3036] = 0;
    exp_62_ram[3037] = 0;
    exp_62_ram[3038] = 238;
    exp_62_ram[3039] = 0;
    exp_62_ram[3040] = 0;
    exp_62_ram[3041] = 0;
    exp_62_ram[3042] = 0;
    exp_62_ram[3043] = 0;
    exp_62_ram[3044] = 236;
    exp_62_ram[3045] = 252;
    exp_62_ram[3046] = 0;
    exp_62_ram[3047] = 0;
    exp_62_ram[3048] = 248;
    exp_62_ram[3049] = 0;
    exp_62_ram[3050] = 154;
    exp_62_ram[3051] = 227;
    exp_62_ram[3052] = 0;
    exp_62_ram[3053] = 6;
    exp_62_ram[3054] = 6;
    exp_62_ram[3055] = 6;
    exp_62_ram[3056] = 6;
    exp_62_ram[3057] = 5;
    exp_62_ram[3058] = 5;
    exp_62_ram[3059] = 5;
    exp_62_ram[3060] = 5;
    exp_62_ram[3061] = 4;
    exp_62_ram[3062] = 4;
    exp_62_ram[3063] = 4;
    exp_62_ram[3064] = 4;
    exp_62_ram[3065] = 7;
    exp_62_ram[3066] = 0;
    exp_62_ram[3067] = 250;
    exp_62_ram[3068] = 4;
    exp_62_ram[3069] = 4;
    exp_62_ram[3070] = 5;
    exp_62_ram[3071] = 5;
    exp_62_ram[3072] = 5;
    exp_62_ram[3073] = 5;
    exp_62_ram[3074] = 6;
    exp_62_ram[3075] = 0;
    exp_62_ram[3076] = 156;
    exp_62_ram[3077] = 221;
    exp_62_ram[3078] = 222;
    exp_62_ram[3079] = 0;
    exp_62_ram[3080] = 137;
    exp_62_ram[3081] = 252;
    exp_62_ram[3082] = 0;
    exp_62_ram[3083] = 156;
    exp_62_ram[3084] = 219;
    exp_62_ram[3085] = 220;
    exp_62_ram[3086] = 0;
    exp_62_ram[3087] = 255;
    exp_62_ram[3088] = 252;
    exp_62_ram[3089] = 0;
    exp_62_ram[3090] = 157;
    exp_62_ram[3091] = 217;
    exp_62_ram[3092] = 218;
    exp_62_ram[3093] = 0;
    exp_62_ram[3094] = 250;
    exp_62_ram[3095] = 0;
    exp_62_ram[3096] = 157;
    exp_62_ram[3097] = 216;
    exp_62_ram[3098] = 217;
    exp_62_ram[3099] = 0;
    exp_62_ram[3100] = 250;
    exp_62_ram[3101] = 0;
    exp_62_ram[3102] = 158;
    exp_62_ram[3103] = 214;
    exp_62_ram[3104] = 215;
    exp_62_ram[3105] = 0;
    exp_62_ram[3106] = 250;
    exp_62_ram[3107] = 3;
    exp_62_ram[3108] = 250;
    exp_62_ram[3109] = 0;
    exp_62_ram[3110] = 252;
    exp_62_ram[3111] = 251;
    exp_62_ram[3112] = 0;
    exp_62_ram[3113] = 238;
    exp_62_ram[3114] = 0;
    exp_62_ram[3115] = 0;
    exp_62_ram[3116] = 250;
    exp_62_ram[3117] = 250;
    exp_62_ram[3118] = 250;
    exp_62_ram[3119] = 250;
    exp_62_ram[3120] = 0;
    exp_62_ram[3121] = 0;
    exp_62_ram[3122] = 171;
    exp_62_ram[3123] = 158;
    exp_62_ram[3124] = 252;
    exp_62_ram[3125] = 252;
    exp_62_ram[3126] = 252;
    exp_62_ram[3127] = 13;
    exp_62_ram[3128] = 0;
    exp_62_ram[3129] = 156;
    exp_62_ram[3130] = 0;
    exp_62_ram[3131] = 0;
    exp_62_ram[3132] = 253;
    exp_62_ram[3133] = 253;
    exp_62_ram[3134] = 0;
    exp_62_ram[3135] = 0;
    exp_62_ram[3136] = 163;
    exp_62_ram[3137] = 0;
    exp_62_ram[3138] = 0;
    exp_62_ram[3139] = 0;
    exp_62_ram[3140] = 237;
    exp_62_ram[3141] = 0;
    exp_62_ram[3142] = 200;
    exp_62_ram[3143] = 0;
    exp_62_ram[3144] = 0;
    exp_62_ram[3145] = 0;
    exp_62_ram[3146] = 0;
    exp_62_ram[3147] = 0;
    exp_62_ram[3148] = 0;
    exp_62_ram[3149] = 184;
    exp_62_ram[3150] = 0;
    exp_62_ram[3151] = 250;
    exp_62_ram[3152] = 0;
    exp_62_ram[3153] = 237;
    exp_62_ram[3154] = 0;
    exp_62_ram[3155] = 0;
    exp_62_ram[3156] = 253;
    exp_62_ram[3157] = 253;
    exp_62_ram[3158] = 1;
    exp_62_ram[3159] = 0;
    exp_62_ram[3160] = 0;
    exp_62_ram[3161] = 1;
    exp_62_ram[3162] = 0;
    exp_62_ram[3163] = 0;
    exp_62_ram[3164] = 252;
    exp_62_ram[3165] = 252;
    exp_62_ram[3166] = 0;
    exp_62_ram[3167] = 145;
    exp_62_ram[3168] = 0;
    exp_62_ram[3169] = 0;
    exp_62_ram[3170] = 250;
    exp_62_ram[3171] = 250;
    exp_62_ram[3172] = 250;
    exp_62_ram[3173] = 0;
    exp_62_ram[3174] = 237;
    exp_62_ram[3175] = 0;
    exp_62_ram[3176] = 0;
    exp_62_ram[3177] = 196;
    exp_62_ram[3178] = 253;
    exp_62_ram[3179] = 0;
    exp_62_ram[3180] = 252;
    exp_62_ram[3181] = 253;
    exp_62_ram[3182] = 6;
    exp_62_ram[3183] = 242;
    exp_62_ram[3184] = 0;
    exp_62_ram[3185] = 0;
    exp_62_ram[3186] = 5;
    exp_62_ram[3187] = 5;
    exp_62_ram[3188] = 5;
    exp_62_ram[3189] = 5;
    exp_62_ram[3190] = 4;
    exp_62_ram[3191] = 4;
    exp_62_ram[3192] = 6;
    exp_62_ram[3193] = 0;
    exp_62_ram[3194] = 254;
    exp_62_ram[3195] = 0;
    exp_62_ram[3196] = 0;
    exp_62_ram[3197] = 2;
    exp_62_ram[3198] = 0;
    exp_62_ram[3199] = 158;
    exp_62_ram[3200] = 190;
    exp_62_ram[3201] = 0;
    exp_62_ram[3202] = 159;
    exp_62_ram[3203] = 189;
    exp_62_ram[3204] = 0;
    exp_62_ram[3205] = 160;
    exp_62_ram[3206] = 189;
    exp_62_ram[3207] = 0;
    exp_62_ram[3208] = 161;
    exp_62_ram[3209] = 188;
    exp_62_ram[3210] = 0;
    exp_62_ram[3211] = 163;
    exp_62_ram[3212] = 187;
    exp_62_ram[3213] = 0;
    exp_62_ram[3214] = 164;
    exp_62_ram[3215] = 186;
    exp_62_ram[3216] = 0;
    exp_62_ram[3217] = 165;
    exp_62_ram[3218] = 186;
    exp_62_ram[3219] = 175;
    exp_62_ram[3220] = 0;
    exp_62_ram[3221] = 254;
    exp_62_ram[3222] = 254;
    exp_62_ram[3223] = 249;
    exp_62_ram[3224] = 0;
    exp_62_ram[3225] = 248;
    exp_62_ram[3226] = 0;
    exp_62_ram[3227] = 0;
    exp_62_ram[3228] = 238;
    exp_62_ram[3229] = 0;
    exp_62_ram[3230] = 0;
    exp_62_ram[3231] = 0;
    exp_62_ram[3232] = 217;
    exp_62_ram[3233] = 2;
    exp_62_ram[3234] = 220;
    exp_62_ram[3235] = 2;
    exp_62_ram[3236] = 253;
    exp_62_ram[3237] = 1;
    exp_62_ram[3238] = 213;
    exp_62_ram[3239] = 1;
    exp_62_ram[3240] = 13;
    exp_62_ram[3241] = 0;
    exp_62_ram[3242] = 235;
    exp_62_ram[3243] = 0;
    exp_62_ram[3244] = 244;
    exp_62_ram[3245] = 254;
    exp_62_ram[3246] = 0;
    exp_62_ram[3247] = 2;
    exp_62_ram[3248] = 0;
    exp_62_ram[3249] = 254;
    exp_62_ram[3250] = 254;
    exp_62_ram[3251] = 1;
    exp_62_ram[3252] = 1;
    exp_62_ram[3253] = 2;
    exp_62_ram[3254] = 15;
    exp_62_ram[3255] = 0;
    exp_62_ram[3256] = 1;
    exp_62_ram[3257] = 2;
    exp_62_ram[3258] = 0;
    exp_62_ram[3259] = 252;
    exp_62_ram[3260] = 2;
    exp_62_ram[3261] = 2;
    exp_62_ram[3262] = 2;
    exp_62_ram[3263] = 4;
    exp_62_ram[3264] = 252;
    exp_62_ram[3265] = 252;
    exp_62_ram[3266] = 252;
    exp_62_ram[3267] = 252;
    exp_62_ram[3268] = 252;
    exp_62_ram[3269] = 0;
    exp_62_ram[3270] = 0;
    exp_62_ram[3271] = 252;
    exp_62_ram[3272] = 0;
    exp_62_ram[3273] = 252;
    exp_62_ram[3274] = 0;
    exp_62_ram[3275] = 252;
    exp_62_ram[3276] = 0;
    exp_62_ram[3277] = 251;
    exp_62_ram[3278] = 15;
    exp_62_ram[3279] = 253;
    exp_62_ram[3280] = 10;
    exp_62_ram[3281] = 0;
    exp_62_ram[3282] = 251;
    exp_62_ram[3283] = 15;
    exp_62_ram[3284] = 253;
    exp_62_ram[3285] = 10;
    exp_62_ram[3286] = 0;
    exp_62_ram[3287] = 251;
    exp_62_ram[3288] = 15;
    exp_62_ram[3289] = 253;
    exp_62_ram[3290] = 10;
    exp_62_ram[3291] = 253;
    exp_62_ram[3292] = 1;
    exp_62_ram[3293] = 0;
    exp_62_ram[3294] = 251;
    exp_62_ram[3295] = 15;
    exp_62_ram[3296] = 253;
    exp_62_ram[3297] = 10;
    exp_62_ram[3298] = 253;
    exp_62_ram[3299] = 1;
    exp_62_ram[3300] = 0;
    exp_62_ram[3301] = 251;
    exp_62_ram[3302] = 15;
    exp_62_ram[3303] = 253;
    exp_62_ram[3304] = 10;
    exp_62_ram[3305] = 252;
    exp_62_ram[3306] = 251;
    exp_62_ram[3307] = 15;
    exp_62_ram[3308] = 253;
    exp_62_ram[3309] = 10;
    exp_62_ram[3310] = 252;
    exp_62_ram[3311] = 251;
    exp_62_ram[3312] = 15;
    exp_62_ram[3313] = 253;
    exp_62_ram[3314] = 10;
    exp_62_ram[3315] = 252;
    exp_62_ram[3316] = 251;
    exp_62_ram[3317] = 15;
    exp_62_ram[3318] = 253;
    exp_62_ram[3319] = 10;
    exp_62_ram[3320] = 254;
    exp_62_ram[3321] = 21;
    exp_62_ram[3322] = 254;
    exp_62_ram[3323] = 253;
    exp_62_ram[3324] = 0;
    exp_62_ram[3325] = 0;
    exp_62_ram[3326] = 251;
    exp_62_ram[3327] = 254;
    exp_62_ram[3328] = 254;
    exp_62_ram[3329] = 253;
    exp_62_ram[3330] = 0;
    exp_62_ram[3331] = 0;
    exp_62_ram[3332] = 251;
    exp_62_ram[3333] = 254;
    exp_62_ram[3334] = 254;
    exp_62_ram[3335] = 253;
    exp_62_ram[3336] = 0;
    exp_62_ram[3337] = 0;
    exp_62_ram[3338] = 251;
    exp_62_ram[3339] = 254;
    exp_62_ram[3340] = 254;
    exp_62_ram[3341] = 252;
    exp_62_ram[3342] = 0;
    exp_62_ram[3343] = 0;
    exp_62_ram[3344] = 251;
    exp_62_ram[3345] = 254;
    exp_62_ram[3346] = 254;
    exp_62_ram[3347] = 0;
    exp_62_ram[3348] = 230;
    exp_62_ram[3349] = 0;
    exp_62_ram[3350] = 0;
    exp_62_ram[3351] = 253;
    exp_62_ram[3352] = 0;
    exp_62_ram[3353] = 254;
    exp_62_ram[3354] = 0;
    exp_62_ram[3355] = 254;
    exp_62_ram[3356] = 0;
    exp_62_ram[3357] = 228;
    exp_62_ram[3358] = 0;
    exp_62_ram[3359] = 0;
    exp_62_ram[3360] = 253;
    exp_62_ram[3361] = 0;
    exp_62_ram[3362] = 254;
    exp_62_ram[3363] = 4;
    exp_62_ram[3364] = 254;
    exp_62_ram[3365] = 0;
    exp_62_ram[3366] = 225;
    exp_62_ram[3367] = 0;
    exp_62_ram[3368] = 0;
    exp_62_ram[3369] = 253;
    exp_62_ram[3370] = 0;
    exp_62_ram[3371] = 254;
    exp_62_ram[3372] = 2;
    exp_62_ram[3373] = 254;
    exp_62_ram[3374] = 253;
    exp_62_ram[3375] = 0;
    exp_62_ram[3376] = 254;
    exp_62_ram[3377] = 0;
    exp_62_ram[3378] = 254;
    exp_62_ram[3379] = 254;
    exp_62_ram[3380] = 0;
    exp_62_ram[3381] = 222;
    exp_62_ram[3382] = 0;
    exp_62_ram[3383] = 0;
    exp_62_ram[3384] = 253;
    exp_62_ram[3385] = 0;
    exp_62_ram[3386] = 6;
    exp_62_ram[3387] = 254;
    exp_62_ram[3388] = 254;
    exp_62_ram[3389] = 0;
    exp_62_ram[3390] = 219;
    exp_62_ram[3391] = 0;
    exp_62_ram[3392] = 0;
    exp_62_ram[3393] = 253;
    exp_62_ram[3394] = 0;
    exp_62_ram[3395] = 8;
    exp_62_ram[3396] = 254;
    exp_62_ram[3397] = 254;
    exp_62_ram[3398] = 0;
    exp_62_ram[3399] = 217;
    exp_62_ram[3400] = 0;
    exp_62_ram[3401] = 0;
    exp_62_ram[3402] = 253;
    exp_62_ram[3403] = 0;
    exp_62_ram[3404] = 8;
    exp_62_ram[3405] = 254;
    exp_62_ram[3406] = 0;
    exp_62_ram[3407] = 254;
    exp_62_ram[3408] = 254;
    exp_62_ram[3409] = 1;
    exp_62_ram[3410] = 234;
    exp_62_ram[3411] = 0;
    exp_62_ram[3412] = 0;
    exp_62_ram[3413] = 3;
    exp_62_ram[3414] = 3;
    exp_62_ram[3415] = 3;
    exp_62_ram[3416] = 4;
    exp_62_ram[3417] = 0;
    exp_62_ram[3418] = 253;
    exp_62_ram[3419] = 2;
    exp_62_ram[3420] = 2;
    exp_62_ram[3421] = 3;
    exp_62_ram[3422] = 252;
    exp_62_ram[3423] = 0;
    exp_62_ram[3424] = 252;
    exp_62_ram[3425] = 253;
    exp_62_ram[3426] = 11;
    exp_62_ram[3427] = 253;
    exp_62_ram[3428] = 11;
    exp_62_ram[3429] = 2;
    exp_62_ram[3430] = 253;
    exp_62_ram[3431] = 11;
    exp_62_ram[3432] = 0;
    exp_62_ram[3433] = 15;
    exp_62_ram[3434] = 0;
    exp_62_ram[3435] = 208;
    exp_62_ram[3436] = 0;
    exp_62_ram[3437] = 0;
    exp_62_ram[3438] = 253;
    exp_62_ram[3439] = 10;
    exp_62_ram[3440] = 253;
    exp_62_ram[3441] = 11;
    exp_62_ram[3442] = 253;
    exp_62_ram[3443] = 11;
    exp_62_ram[3444] = 2;
    exp_62_ram[3445] = 253;
    exp_62_ram[3446] = 11;
    exp_62_ram[3447] = 0;
    exp_62_ram[3448] = 15;
    exp_62_ram[3449] = 0;
    exp_62_ram[3450] = 204;
    exp_62_ram[3451] = 0;
    exp_62_ram[3452] = 0;
    exp_62_ram[3453] = 253;
    exp_62_ram[3454] = 10;
    exp_62_ram[3455] = 253;
    exp_62_ram[3456] = 11;
    exp_62_ram[3457] = 0;
    exp_62_ram[3458] = 15;
    exp_62_ram[3459] = 0;
    exp_62_ram[3460] = 202;
    exp_62_ram[3461] = 0;
    exp_62_ram[3462] = 0;
    exp_62_ram[3463] = 253;
    exp_62_ram[3464] = 10;
    exp_62_ram[3465] = 253;
    exp_62_ram[3466] = 251;
    exp_62_ram[3467] = 254;
    exp_62_ram[3468] = 253;
    exp_62_ram[3469] = 11;
    exp_62_ram[3470] = 254;
    exp_62_ram[3471] = 0;
    exp_62_ram[3472] = 15;
    exp_62_ram[3473] = 253;
    exp_62_ram[3474] = 11;
    exp_62_ram[3475] = 64;
    exp_62_ram[3476] = 15;
    exp_62_ram[3477] = 0;
    exp_62_ram[3478] = 197;
    exp_62_ram[3479] = 0;
    exp_62_ram[3480] = 0;
    exp_62_ram[3481] = 253;
    exp_62_ram[3482] = 0;
    exp_62_ram[3483] = 3;
    exp_62_ram[3484] = 253;
    exp_62_ram[3485] = 11;
    exp_62_ram[3486] = 64;
    exp_62_ram[3487] = 15;
    exp_62_ram[3488] = 253;
    exp_62_ram[3489] = 11;
    exp_62_ram[3490] = 0;
    exp_62_ram[3491] = 15;
    exp_62_ram[3492] = 0;
    exp_62_ram[3493] = 194;
    exp_62_ram[3494] = 0;
    exp_62_ram[3495] = 254;
    exp_62_ram[3496] = 253;
    exp_62_ram[3497] = 11;
    exp_62_ram[3498] = 254;
    exp_62_ram[3499] = 0;
    exp_62_ram[3500] = 15;
    exp_62_ram[3501] = 253;
    exp_62_ram[3502] = 11;
    exp_62_ram[3503] = 64;
    exp_62_ram[3504] = 15;
    exp_62_ram[3505] = 0;
    exp_62_ram[3506] = 190;
    exp_62_ram[3507] = 0;
    exp_62_ram[3508] = 0;
    exp_62_ram[3509] = 253;
    exp_62_ram[3510] = 0;
    exp_62_ram[3511] = 4;
    exp_62_ram[3512] = 253;
    exp_62_ram[3513] = 11;
    exp_62_ram[3514] = 64;
    exp_62_ram[3515] = 15;
    exp_62_ram[3516] = 253;
    exp_62_ram[3517] = 11;
    exp_62_ram[3518] = 0;
    exp_62_ram[3519] = 15;
    exp_62_ram[3520] = 0;
    exp_62_ram[3521] = 187;
    exp_62_ram[3522] = 0;
    exp_62_ram[3523] = 254;
    exp_62_ram[3524] = 253;
    exp_62_ram[3525] = 11;
    exp_62_ram[3526] = 254;
    exp_62_ram[3527] = 0;
    exp_62_ram[3528] = 15;
    exp_62_ram[3529] = 253;
    exp_62_ram[3530] = 11;
    exp_62_ram[3531] = 64;
    exp_62_ram[3532] = 15;
    exp_62_ram[3533] = 0;
    exp_62_ram[3534] = 183;
    exp_62_ram[3535] = 0;
    exp_62_ram[3536] = 0;
    exp_62_ram[3537] = 253;
    exp_62_ram[3538] = 0;
    exp_62_ram[3539] = 1;
    exp_62_ram[3540] = 253;
    exp_62_ram[3541] = 11;
    exp_62_ram[3542] = 64;
    exp_62_ram[3543] = 15;
    exp_62_ram[3544] = 253;
    exp_62_ram[3545] = 11;
    exp_62_ram[3546] = 0;
    exp_62_ram[3547] = 15;
    exp_62_ram[3548] = 0;
    exp_62_ram[3549] = 180;
    exp_62_ram[3550] = 0;
    exp_62_ram[3551] = 254;
    exp_62_ram[3552] = 254;
    exp_62_ram[3553] = 253;
    exp_62_ram[3554] = 0;
    exp_62_ram[3555] = 0;
    exp_62_ram[3556] = 254;
    exp_62_ram[3557] = 253;
    exp_62_ram[3558] = 11;
    exp_62_ram[3559] = 254;
    exp_62_ram[3560] = 0;
    exp_62_ram[3561] = 15;
    exp_62_ram[3562] = 253;
    exp_62_ram[3563] = 11;
    exp_62_ram[3564] = 64;
    exp_62_ram[3565] = 15;
    exp_62_ram[3566] = 0;
    exp_62_ram[3567] = 175;
    exp_62_ram[3568] = 0;
    exp_62_ram[3569] = 0;
    exp_62_ram[3570] = 253;
    exp_62_ram[3571] = 0;
    exp_62_ram[3572] = 6;
    exp_62_ram[3573] = 253;
    exp_62_ram[3574] = 11;
    exp_62_ram[3575] = 64;
    exp_62_ram[3576] = 15;
    exp_62_ram[3577] = 253;
    exp_62_ram[3578] = 11;
    exp_62_ram[3579] = 0;
    exp_62_ram[3580] = 15;
    exp_62_ram[3581] = 0;
    exp_62_ram[3582] = 171;
    exp_62_ram[3583] = 0;
    exp_62_ram[3584] = 254;
    exp_62_ram[3585] = 253;
    exp_62_ram[3586] = 11;
    exp_62_ram[3587] = 254;
    exp_62_ram[3588] = 0;
    exp_62_ram[3589] = 15;
    exp_62_ram[3590] = 253;
    exp_62_ram[3591] = 11;
    exp_62_ram[3592] = 64;
    exp_62_ram[3593] = 15;
    exp_62_ram[3594] = 0;
    exp_62_ram[3595] = 168;
    exp_62_ram[3596] = 0;
    exp_62_ram[3597] = 0;
    exp_62_ram[3598] = 253;
    exp_62_ram[3599] = 0;
    exp_62_ram[3600] = 9;
    exp_62_ram[3601] = 253;
    exp_62_ram[3602] = 11;
    exp_62_ram[3603] = 64;
    exp_62_ram[3604] = 15;
    exp_62_ram[3605] = 253;
    exp_62_ram[3606] = 11;
    exp_62_ram[3607] = 0;
    exp_62_ram[3608] = 15;
    exp_62_ram[3609] = 0;
    exp_62_ram[3610] = 164;
    exp_62_ram[3611] = 0;
    exp_62_ram[3612] = 254;
    exp_62_ram[3613] = 253;
    exp_62_ram[3614] = 11;
    exp_62_ram[3615] = 254;
    exp_62_ram[3616] = 0;
    exp_62_ram[3617] = 15;
    exp_62_ram[3618] = 253;
    exp_62_ram[3619] = 11;
    exp_62_ram[3620] = 64;
    exp_62_ram[3621] = 15;
    exp_62_ram[3622] = 0;
    exp_62_ram[3623] = 161;
    exp_62_ram[3624] = 0;
    exp_62_ram[3625] = 0;
    exp_62_ram[3626] = 253;
    exp_62_ram[3627] = 0;
    exp_62_ram[3628] = 8;
    exp_62_ram[3629] = 253;
    exp_62_ram[3630] = 11;
    exp_62_ram[3631] = 64;
    exp_62_ram[3632] = 15;
    exp_62_ram[3633] = 253;
    exp_62_ram[3634] = 11;
    exp_62_ram[3635] = 0;
    exp_62_ram[3636] = 15;
    exp_62_ram[3637] = 0;
    exp_62_ram[3638] = 157;
    exp_62_ram[3639] = 0;
    exp_62_ram[3640] = 254;
    exp_62_ram[3641] = 254;
    exp_62_ram[3642] = 4;
    exp_62_ram[3643] = 15;
    exp_62_ram[3644] = 0;
    exp_62_ram[3645] = 2;
    exp_62_ram[3646] = 2;
    exp_62_ram[3647] = 3;
    exp_62_ram[3648] = 0;
    exp_62_ram[3649] = 254;
    exp_62_ram[3650] = 0;
    exp_62_ram[3651] = 0;
    exp_62_ram[3652] = 2;
    exp_62_ram[3653] = 194;
    exp_62_ram[3654] = 0;
    exp_62_ram[3655] = 254;
    exp_62_ram[3656] = 254;
    exp_62_ram[3657] = 3;
    exp_62_ram[3658] = 0;
    exp_62_ram[3659] = 0;
    exp_62_ram[3660] = 240;
    exp_62_ram[3661] = 6;
    exp_62_ram[3662] = 254;
    exp_62_ram[3663] = 3;
    exp_62_ram[3664] = 0;
    exp_62_ram[3665] = 0;
    exp_62_ram[3666] = 242;
    exp_62_ram[3667] = 4;
    exp_62_ram[3668] = 254;
    exp_62_ram[3669] = 3;
    exp_62_ram[3670] = 0;
    exp_62_ram[3671] = 0;
    exp_62_ram[3672] = 243;
    exp_62_ram[3673] = 3;
    exp_62_ram[3674] = 254;
    exp_62_ram[3675] = 3;
    exp_62_ram[3676] = 0;
    exp_62_ram[3677] = 0;
    exp_62_ram[3678] = 245;
    exp_62_ram[3679] = 1;
    exp_62_ram[3680] = 254;
    exp_62_ram[3681] = 3;
    exp_62_ram[3682] = 248;
    exp_62_ram[3683] = 0;
    exp_62_ram[3684] = 247;
    exp_62_ram[3685] = 0;
    exp_62_ram[3686] = 1;
    exp_62_ram[3687] = 1;
    exp_62_ram[3688] = 2;
    exp_62_ram[3689] = 0;
    exp_62_ram[3690] = 254;
    exp_62_ram[3691] = 0;
    exp_62_ram[3692] = 0;
    exp_62_ram[3693] = 2;
    exp_62_ram[3694] = 184;
    exp_62_ram[3695] = 0;
    exp_62_ram[3696] = 254;
    exp_62_ram[3697] = 254;
    exp_62_ram[3698] = 0;
    exp_62_ram[3699] = 209;
    exp_62_ram[3700] = 0;
    exp_62_ram[3701] = 4;
    exp_62_ram[3702] = 0;
    exp_62_ram[3703] = 0;
    exp_62_ram[3704] = 249;
    exp_62_ram[3705] = 4;
    exp_62_ram[3706] = 254;
    exp_62_ram[3707] = 0;
    exp_62_ram[3708] = 206;
    exp_62_ram[3709] = 0;
    exp_62_ram[3710] = 4;
    exp_62_ram[3711] = 0;
    exp_62_ram[3712] = 0;
    exp_62_ram[3713] = 250;
    exp_62_ram[3714] = 2;
    exp_62_ram[3715] = 254;
    exp_62_ram[3716] = 0;
    exp_62_ram[3717] = 204;
    exp_62_ram[3718] = 0;
    exp_62_ram[3719] = 4;
    exp_62_ram[3720] = 248;
    exp_62_ram[3721] = 0;
    exp_62_ram[3722] = 252;
    exp_62_ram[3723] = 0;
    exp_62_ram[3724] = 1;
    exp_62_ram[3725] = 1;
    exp_62_ram[3726] = 2;
    exp_62_ram[3727] = 0;
    exp_62_ram[3728] = 254;
    exp_62_ram[3729] = 0;
    exp_62_ram[3730] = 0;
    exp_62_ram[3731] = 2;
    exp_62_ram[3732] = 175;
    exp_62_ram[3733] = 0;
    exp_62_ram[3734] = 254;
    exp_62_ram[3735] = 254;
    exp_62_ram[3736] = 0;
    exp_62_ram[3737] = 189;
    exp_62_ram[3738] = 0;
    exp_62_ram[3739] = 254;
    exp_62_ram[3740] = 254;
    exp_62_ram[3741] = 0;
    exp_62_ram[3742] = 198;
    exp_62_ram[3743] = 0;
    exp_62_ram[3744] = 15;
    exp_62_ram[3745] = 0;
    exp_62_ram[3746] = 1;
    exp_62_ram[3747] = 1;
    exp_62_ram[3748] = 2;
    exp_62_ram[3749] = 0;
    exp_62_ram[3750] = 254;
    exp_62_ram[3751] = 0;
    exp_62_ram[3752] = 0;
    exp_62_ram[3753] = 2;
    exp_62_ram[3754] = 0;
    exp_62_ram[3755] = 15;
    exp_62_ram[3756] = 0;
    exp_62_ram[3757] = 15;
    exp_62_ram[3758] = 0;
    exp_62_ram[3759] = 15;
    exp_62_ram[3760] = 0;
    exp_62_ram[3761] = 15;
    exp_62_ram[3762] = 0;
    exp_62_ram[3763] = 16;
    exp_62_ram[3764] = 0;
    exp_62_ram[3765] = 16;
    exp_62_ram[3766] = 0;
    exp_62_ram[3767] = 16;
    exp_62_ram[3768] = 0;
    exp_62_ram[3769] = 16;
    exp_62_ram[3770] = 0;
    exp_62_ram[3771] = 16;
    exp_62_ram[3772] = 0;
    exp_62_ram[3773] = 16;
    exp_62_ram[3774] = 0;
    exp_62_ram[3775] = 0;
    exp_62_ram[3776] = 0;
    exp_62_ram[3777] = 0;
    exp_62_ram[3778] = 0;
    exp_62_ram[3779] = 0;
    exp_62_ram[3780] = 0;
    exp_62_ram[3781] = 3;
    exp_62_ram[3782] = 253;
    exp_62_ram[3783] = 0;
    exp_62_ram[3784] = 166;
    exp_62_ram[3785] = 172;
    exp_62_ram[3786] = 0;
    exp_62_ram[3787] = 16;
    exp_62_ram[3788] = 0;
    exp_62_ram[3789] = 156;
    exp_62_ram[3790] = 0;
    exp_62_ram[3791] = 16;
    exp_62_ram[3792] = 0;
    exp_62_ram[3793] = 155;
    exp_62_ram[3794] = 0;
    exp_62_ram[3795] = 16;
    exp_62_ram[3796] = 0;
    exp_62_ram[3797] = 154;
    exp_62_ram[3798] = 0;
    exp_62_ram[3799] = 167;
    exp_62_ram[3800] = 168;
    exp_62_ram[3801] = 0;
    exp_62_ram[3802] = 1;
    exp_62_ram[3803] = 1;
    exp_62_ram[3804] = 2;
    exp_62_ram[3805] = 0;
    exp_62_ram[3806] = 254;
    exp_62_ram[3807] = 0;
    exp_62_ram[3808] = 0;
    exp_62_ram[3809] = 2;
    exp_62_ram[3810] = 0;
    exp_62_ram[3811] = 0;
    exp_62_ram[3812] = 240;
    exp_62_ram[3813] = 14;
    exp_62_ram[3814] = 0;
    exp_62_ram[3815] = 0;
    exp_62_ram[3816] = 242;
    exp_62_ram[3817] = 14;
    exp_62_ram[3818] = 0;
    exp_62_ram[3819] = 0;
    exp_62_ram[3820] = 243;
    exp_62_ram[3821] = 14;
    exp_62_ram[3822] = 0;
    exp_62_ram[3823] = 0;
    exp_62_ram[3824] = 250;
    exp_62_ram[3825] = 14;
    exp_62_ram[3826] = 0;
    exp_62_ram[3827] = 4;
    exp_62_ram[3828] = 16;
    exp_62_ram[3829] = 0;
    exp_62_ram[3830] = 4;
    exp_62_ram[3831] = 16;
    exp_62_ram[3832] = 0;
    exp_62_ram[3833] = 4;
    exp_62_ram[3834] = 16;
    exp_62_ram[3835] = 0;
    exp_62_ram[3836] = 4;
    exp_62_ram[3837] = 16;
    exp_62_ram[3838] = 0;
    exp_62_ram[3839] = 4;
    exp_62_ram[3840] = 16;
    exp_62_ram[3841] = 0;
    exp_62_ram[3842] = 4;
    exp_62_ram[3843] = 16;
    exp_62_ram[3844] = 232;
    exp_62_ram[3845] = 0;
    exp_62_ram[3846] = 167;
    exp_62_ram[3847] = 156;
    exp_62_ram[3848] = 0;
    exp_62_ram[3849] = 168;
    exp_62_ram[3850] = 156;
    exp_62_ram[3851] = 0;
    exp_62_ram[3852] = 170;
    exp_62_ram[3853] = 155;
    exp_62_ram[3854] = 0;
    exp_62_ram[3855] = 174;
    exp_62_ram[3856] = 154;
    exp_62_ram[3857] = 0;
    exp_62_ram[3858] = 176;
    exp_62_ram[3859] = 153;
    exp_62_ram[3860] = 0;
    exp_62_ram[3861] = 180;
    exp_62_ram[3862] = 153;
    exp_62_ram[3863] = 0;
    exp_62_ram[3864] = 184;
    exp_62_ram[3865] = 152;
    exp_62_ram[3866] = 254;
    exp_62_ram[3867] = 141;
    exp_62_ram[3868] = 0;
    exp_62_ram[3869] = 254;
    exp_62_ram[3870] = 254;
    exp_62_ram[3871] = 0;
    exp_62_ram[3872] = 155;
    exp_62_ram[3873] = 0;
    exp_62_ram[3874] = 10;
    exp_62_ram[3875] = 254;
    exp_62_ram[3876] = 4;
    exp_62_ram[3877] = 0;
    exp_62_ram[3878] = 3;
    exp_62_ram[3879] = 11;
    exp_62_ram[3880] = 4;
    exp_62_ram[3881] = 0;
    exp_62_ram[3882] = 133;
    exp_62_ram[3883] = 0;
    exp_62_ram[3884] = 3;
    exp_62_ram[3885] = 11;
    exp_62_ram[3886] = 4;
    exp_62_ram[3887] = 0;
    exp_62_ram[3888] = 132;
    exp_62_ram[3889] = 0;
    exp_62_ram[3890] = 3;
    exp_62_ram[3891] = 11;
    exp_62_ram[3892] = 4;
    exp_62_ram[3893] = 0;
    exp_62_ram[3894] = 130;
    exp_62_ram[3895] = 0;
    exp_62_ram[3896] = 184;
    exp_62_ram[3897] = 144;
    exp_62_ram[3898] = 254;
    exp_62_ram[3899] = 0;
    exp_62_ram[3900] = 158;
    exp_62_ram[3901] = 0;
    exp_62_ram[3902] = 15;
    exp_62_ram[3903] = 0;
    exp_62_ram[3904] = 0;
    exp_62_ram[3905] = 3;
    exp_62_ram[3906] = 134;
    exp_62_ram[3907] = 0;
    exp_62_ram[3908] = 0;
    exp_62_ram[3909] = 254;
    exp_62_ram[3910] = 254;
    exp_62_ram[3911] = 4;
    exp_62_ram[3912] = 0;
    exp_62_ram[3913] = 254;
    exp_62_ram[3914] = 0;
    exp_62_ram[3915] = 253;
    exp_62_ram[3916] = 243;
    exp_62_ram[3917] = 254;
    exp_62_ram[3918] = 0;
    exp_62_ram[3919] = 254;
    exp_62_ram[3920] = 242;
    exp_62_ram[3921] = 254;
    exp_62_ram[3922] = 253;
    exp_62_ram[3923] = 0;
    exp_62_ram[3924] = 240;
    exp_62_ram[3925] = 254;
    exp_62_ram[3926] = 3;
    exp_62_ram[3927] = 4;
    exp_62_ram[3928] = 0;
    exp_62_ram[3929] = 185;
    exp_62_ram[3930] = 136;
    exp_62_ram[3931] = 185;
    exp_62_ram[3932] = 0;
    exp_62_ram[3933] = 0;
    exp_62_ram[3934] = 14;
    exp_62_ram[3935] = 184;
    exp_62_ram[3936] = 0;
    exp_62_ram[3937] = 0;
    exp_62_ram[3938] = 14;
    exp_62_ram[3939] = 183;
    exp_62_ram[3940] = 0;
    exp_62_ram[3941] = 0;
    exp_62_ram[3942] = 14;
    exp_62_ram[3943] = 207;
    exp_62_ram[3944] = 254;
    exp_62_ram[3945] = 236;
    exp_62_ram[3946] = 254;
    exp_62_ram[3947] = 3;
    exp_62_ram[3948] = 2;
    exp_62_ram[3949] = 0;
    exp_62_ram[3950] = 185;
    exp_62_ram[3951] = 130;
    exp_62_ram[3952] = 190;
    exp_62_ram[3953] = 0;
    exp_62_ram[3954] = 0;
    exp_62_ram[3955] = 14;
    exp_62_ram[3956] = 204;
    exp_62_ram[3957] = 254;
    exp_62_ram[3958] = 233;
    exp_62_ram[3959] = 254;
    exp_62_ram[3960] = 3;
    exp_62_ram[3961] = 4;
    exp_62_ram[3962] = 0;
    exp_62_ram[3963] = 185;
    exp_62_ram[3964] = 255;
    exp_62_ram[3965] = 196;
    exp_62_ram[3966] = 0;
    exp_62_ram[3967] = 0;
    exp_62_ram[3968] = 0;
    exp_62_ram[3969] = 16;
    exp_62_ram[3970] = 195;
    exp_62_ram[3971] = 0;
    exp_62_ram[3972] = 0;
    exp_62_ram[3973] = 0;
    exp_62_ram[3974] = 16;
    exp_62_ram[3975] = 194;
    exp_62_ram[3976] = 0;
    exp_62_ram[3977] = 0;
    exp_62_ram[3978] = 0;
    exp_62_ram[3979] = 16;
    exp_62_ram[3980] = 198;
    exp_62_ram[3981] = 254;
    exp_62_ram[3982] = 227;
    exp_62_ram[3983] = 254;
    exp_62_ram[3984] = 3;
    exp_62_ram[3985] = 226;
    exp_62_ram[3986] = 0;
    exp_62_ram[3987] = 185;
    exp_62_ram[3988] = 249;
    exp_62_ram[3989] = 190;
    exp_62_ram[3990] = 0;
    exp_62_ram[3991] = 0;
    exp_62_ram[3992] = 0;
    exp_62_ram[3993] = 16;
    exp_62_ram[3994] = 189;
    exp_62_ram[3995] = 0;
    exp_62_ram[3996] = 0;
    exp_62_ram[3997] = 0;
    exp_62_ram[3998] = 16;
    exp_62_ram[3999] = 188;
    exp_62_ram[4000] = 0;
    exp_62_ram[4001] = 0;
    exp_62_ram[4002] = 0;
    exp_62_ram[4003] = 16;
    exp_62_ram[4004] = 192;
    exp_62_ram[4005] = 254;
    exp_62_ram[4006] = 221;
    exp_62_ram[4007] = 0;
    exp_62_ram[4008] = 0;
    exp_62_ram[4009] = 2;
    exp_62_ram[4010] = 255;
    exp_62_ram[4011] = 2;
    exp_62_ram[4012] = 0;
    exp_62_ram[4013] = 0;
    exp_62_ram[4014] = 0;
    exp_62_ram[4015] = 64;
    exp_62_ram[4016] = 1;
    exp_62_ram[4017] = 0;
    exp_62_ram[4018] = 254;
    exp_62_ram[4019] = 255;
    exp_62_ram[4020] = 0;
    exp_62_ram[4021] = 254;
    exp_62_ram[4022] = 2;
    exp_62_ram[4023] = 2;
    exp_62_ram[4024] = 3;
    exp_62_ram[4025] = 4;
    exp_62_ram[4026] = 5;
    exp_62_ram[4027] = 0;
    exp_62_ram[4028] = 0;
    exp_62_ram[4029] = 0;
    exp_62_ram[4030] = 0;
    exp_62_ram[4031] = 0;
    exp_62_ram[4032] = 0;
    exp_62_ram[4033] = 70;
    exp_62_ram[4034] = 81;
    exp_62_ram[4035] = 84;
    exp_62_ram[4036] = 72;
    exp_62_ram[4037] = 80;
    exp_62_ram[4038] = 82;
    exp_62_ram[4039] = 0;
    exp_62_ram[4040] = 75;
    exp_62_ram[4041] = 85;
    exp_62_ram[4042] = 72;
    exp_62_ram[4043] = 67;
    exp_62_ram[4044] = 78;
    exp_62_ram[4045] = 86;
    exp_62_ram[4046] = 0;
    exp_62_ram[4047] = 72;
    exp_62_ram[4048] = 80;
    exp_62_ram[4049] = 86;
    exp_62_ram[4050] = 69;
    exp_62_ram[4051] = 65;
    exp_62_ram[4052] = 83;
    exp_62_ram[4053] = 0;
    exp_62_ram[4054] = 86;
    exp_62_ram[4055] = 65;
    exp_62_ram[4056] = 73;
    exp_62_ram[4057] = 76;
    exp_62_ram[4058] = 71;
    exp_62_ram[4059] = 77;
    exp_62_ram[4060] = 0;
    exp_62_ram[4061] = 82;
    exp_62_ram[4062] = 89;
    exp_62_ram[4063] = 68;
    exp_62_ram[4064] = 88;
    exp_62_ram[4065] = 74;
    exp_62_ram[4066] = 69;
    exp_62_ram[4067] = 0;
    exp_62_ram[4068] = 90;
    exp_62_ram[4069] = 88;
    exp_62_ram[4070] = 70;
    exp_62_ram[4071] = 85;
    exp_62_ram[4072] = 83;
    exp_62_ram[4073] = 72;
    exp_62_ram[4074] = 0;
    exp_62_ram[4075] = 72;
    exp_62_ram[4076] = 68;
    exp_62_ram[4077] = 71;
    exp_62_ram[4078] = 73;
    exp_62_ram[4079] = 90;
    exp_62_ram[4080] = 74;
    exp_62_ram[4081] = 0;
    exp_62_ram[4082] = 74;
    exp_62_ram[4083] = 89;
    exp_62_ram[4084] = 90;
    exp_62_ram[4085] = 67;
    exp_62_ram[4086] = 81;
    exp_62_ram[4087] = 77;
    exp_62_ram[4088] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_60) begin
      exp_62_ram[exp_56] <= exp_58;
    end
  end
  assign exp_62 = exp_62_ram[exp_57];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_88) begin
        exp_62_ram[exp_84] <= exp_86;
    end
  end
  assign exp_90 = exp_62_ram[exp_85];
  assign exp_61 = exp_129;
  assign exp_129 = 1;
  assign exp_57 = exp_128;
  assign exp_128 = exp_18[31:2];
  assign exp_18 = exp_9;
  assign exp_60 = exp_124;
  assign exp_124 = exp_122 & exp_123;
  assign exp_122 = exp_22 & exp_23;
  assign exp_123 = exp_24[3:3];
  assign exp_24 = exp_13;
  assign exp_13 = exp_536;

      reg [3:0] exp_536_reg = 0;
      always@(posedge clk) begin
        if (exp_529) begin
          exp_536_reg <= exp_527;
        end
      end
      assign exp_536 = exp_536_reg;
      assign exp_527 = exp_818;

  reg [3:0] exp_818_reg;
  always@(*) begin
    case (exp_670)
      0:exp_818_reg <= exp_805;
      1:exp_818_reg <= exp_810;
      2:exp_818_reg <= exp_811;
      3:exp_818_reg <= exp_812;
      4:exp_818_reg <= exp_813;
      5:exp_818_reg <= exp_814;
      6:exp_818_reg <= exp_815;
      7:exp_818_reg <= exp_816;
      default:exp_818_reg <= exp_817;
    endcase
  end
  assign exp_818 = exp_818_reg;
  assign exp_817 = 0;
  assign exp_805 = exp_801 << exp_804;
  assign exp_801 = 1;
  assign exp_804 = exp_803 + exp_802;
  assign exp_803 = 0;
  assign exp_802 = exp_738[1:0];
  assign exp_810 = exp_806 << exp_809;
  assign exp_806 = 3;
  assign exp_809 = exp_808 + exp_807;
  assign exp_808 = 0;
  assign exp_807 = exp_738[1:1];
  assign exp_811 = 15;
  assign exp_812 = 0;
  assign exp_813 = 0;
  assign exp_814 = 0;
  assign exp_815 = 0;
  assign exp_816 = 0;
  assign exp_56 = exp_120;
  assign exp_120 = exp_18[31:2];
  assign exp_58 = exp_121;
  assign exp_121 = exp_19[31:24];
  assign exp_19 = exp_10;
  assign exp_10 = exp_533;

      reg [31:0] exp_533_reg = 0;
      always@(posedge clk) begin
        if (exp_529) begin
          exp_533_reg <= exp_522;
        end
      end
      assign exp_533 = exp_533_reg;
      assign exp_522 = exp_800;

  reg [31:0] exp_800_reg;
  always@(*) begin
    case (exp_670)
      0:exp_800_reg <= exp_787;
      1:exp_800_reg <= exp_791;
      2:exp_800_reg <= exp_793;
      3:exp_800_reg <= exp_794;
      4:exp_800_reg <= exp_795;
      5:exp_800_reg <= exp_796;
      6:exp_800_reg <= exp_797;
      7:exp_800_reg <= exp_798;
      default:exp_800_reg <= exp_799;
    endcase
  end
  assign exp_800 = exp_800_reg;
  assign exp_799 = 0;

  reg [31:0] exp_787_reg;
  always@(*) begin
    case (exp_741)
      0:exp_787_reg <= exp_773;
      1:exp_787_reg <= exp_781;
      2:exp_787_reg <= exp_783;
      3:exp_787_reg <= exp_785;
      default:exp_787_reg <= exp_786;
    endcase
  end
  assign exp_787 = exp_787_reg;
  assign exp_786 = 0;
  assign exp_773 = exp_772;
  assign exp_772 = exp_771 + exp_770;
  assign exp_771 = 0;
  assign exp_770 = exp_660[7:0];

      reg [31:0] exp_660_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_660_reg <= exp_603;
        end
      end
      assign exp_660 = exp_660_reg;
      assign exp_781 = exp_773 << exp_780;
  assign exp_780 = 8;
  assign exp_783 = exp_773 << exp_782;
  assign exp_782 = 16;
  assign exp_785 = exp_773 << exp_784;
  assign exp_784 = 24;

  reg [31:0] exp_791_reg;
  always@(*) begin
    case (exp_744)
      0:exp_791_reg <= exp_777;
      1:exp_791_reg <= exp_789;
      default:exp_791_reg <= exp_790;
    endcase
  end
  assign exp_791 = exp_791_reg;
  assign exp_744 = exp_743 + exp_742;
  assign exp_743 = 0;
  assign exp_742 = exp_738[1:1];
  assign exp_790 = 0;
  assign exp_777 = exp_776;
  assign exp_776 = exp_775 + exp_774;
  assign exp_775 = 0;
  assign exp_774 = exp_660[15:0];
  assign exp_789 = exp_777 << exp_788;
  assign exp_788 = 16;
  assign exp_793 = exp_792 + exp_779;
  assign exp_792 = 0;
  assign exp_779 = exp_778 + exp_660;
  assign exp_778 = 0;
  assign exp_794 = 0;
  assign exp_795 = 0;
  assign exp_796 = 0;
  assign exp_797 = 0;
  assign exp_798 = 0;

  //Create RAM
  reg [7:0] exp_55_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_55_ram[0] = 0;
    exp_55_ram[1] = 0;
    exp_55_ram[2] = 0;
    exp_55_ram[3] = 0;
    exp_55_ram[4] = 0;
    exp_55_ram[5] = 0;
    exp_55_ram[6] = 0;
    exp_55_ram[7] = 0;
    exp_55_ram[8] = 0;
    exp_55_ram[9] = 0;
    exp_55_ram[10] = 0;
    exp_55_ram[11] = 0;
    exp_55_ram[12] = 0;
    exp_55_ram[13] = 0;
    exp_55_ram[14] = 0;
    exp_55_ram[15] = 0;
    exp_55_ram[16] = 0;
    exp_55_ram[17] = 0;
    exp_55_ram[18] = 0;
    exp_55_ram[19] = 0;
    exp_55_ram[20] = 0;
    exp_55_ram[21] = 0;
    exp_55_ram[22] = 0;
    exp_55_ram[23] = 0;
    exp_55_ram[24] = 0;
    exp_55_ram[25] = 0;
    exp_55_ram[26] = 0;
    exp_55_ram[27] = 0;
    exp_55_ram[28] = 0;
    exp_55_ram[29] = 0;
    exp_55_ram[30] = 0;
    exp_55_ram[31] = 0;
    exp_55_ram[32] = 1;
    exp_55_ram[33] = 64;
    exp_55_ram[34] = 0;
    exp_55_ram[35] = 5;
    exp_55_ram[36] = 5;
    exp_55_ram[37] = 6;
    exp_55_ram[38] = 6;
    exp_55_ram[39] = 8;
    exp_55_ram[40] = 6;
    exp_55_ram[41] = 0;
    exp_55_ram[42] = 70;
    exp_55_ram[43] = 197;
    exp_55_ram[44] = 1;
    exp_55_ram[45] = 230;
    exp_55_ram[46] = 240;
    exp_55_ram[47] = 199;
    exp_55_ram[48] = 55;
    exp_55_ram[49] = 230;
    exp_55_ram[50] = 166;
    exp_55_ram[51] = 6;
    exp_55_ram[52] = 0;
    exp_55_ram[53] = 230;
    exp_55_ram[54] = 229;
    exp_55_ram[55] = 229;
    exp_55_ram[56] = 215;
    exp_55_ram[57] = 232;
    exp_55_ram[58] = 214;
    exp_55_ram[59] = 183;
    exp_55_ram[60] = 216;
    exp_55_ram[61] = 8;
    exp_55_ram[62] = 21;
    exp_55_ram[63] = 8;
    exp_55_ram[64] = 6;
    exp_55_ram[65] = 3;
    exp_55_ram[66] = 21;
    exp_55_ram[67] = 6;
    exp_55_ram[68] = 214;
    exp_55_ram[69] = 7;
    exp_55_ram[70] = 247;
    exp_55_ram[71] = 183;
    exp_55_ram[72] = 7;
    exp_55_ram[73] = 246;
    exp_55_ram[74] = 7;
    exp_55_ram[75] = 183;
    exp_55_ram[76] = 230;
    exp_55_ram[77] = 7;
    exp_55_ram[78] = 183;
    exp_55_ram[79] = 23;
    exp_55_ram[80] = 3;
    exp_55_ram[81] = 3;
    exp_55_ram[82] = 23;
    exp_55_ram[83] = 7;
    exp_55_ram[84] = 103;
    exp_55_ram[85] = 246;
    exp_55_ram[86] = 7;
    exp_55_ram[87] = 211;
    exp_55_ram[88] = 104;
    exp_55_ram[89] = 247;
    exp_55_ram[90] = 3;
    exp_55_ram[91] = 211;
    exp_55_ram[92] = 231;
    exp_55_ram[93] = 5;
    exp_55_ram[94] = 197;
    exp_55_ram[95] = 0;
    exp_55_ram[96] = 64;
    exp_55_ram[97] = 0;
    exp_55_ram[98] = 0;
    exp_55_ram[99] = 166;
    exp_55_ram[100] = 128;
    exp_55_ram[101] = 31;
    exp_55_ram[102] = 6;
    exp_55_ram[103] = 16;
    exp_55_ram[104] = 199;
    exp_55_ram[105] = 1;
    exp_55_ram[106] = 232;
    exp_55_ram[107] = 240;
    exp_55_ram[108] = 7;
    exp_55_ram[109] = 128;
    exp_55_ram[110] = 168;
    exp_55_ram[111] = 230;
    exp_55_ram[112] = 6;
    exp_55_ram[113] = 0;
    exp_55_ram[114] = 167;
    exp_55_ram[115] = 230;
    exp_55_ram[116] = 230;
    exp_55_ram[117] = 7;
    exp_55_ram[118] = 16;
    exp_55_ram[119] = 8;
    exp_55_ram[120] = 8;
    exp_55_ram[121] = 6;
    exp_55_ram[122] = 3;
    exp_55_ram[123] = 23;
    exp_55_ram[124] = 23;
    exp_55_ram[125] = 6;
    exp_55_ram[126] = 230;
    exp_55_ram[127] = 246;
    exp_55_ram[128] = 7;
    exp_55_ram[129] = 199;
    exp_55_ram[130] = 7;
    exp_55_ram[131] = 247;
    exp_55_ram[132] = 7;
    exp_55_ram[133] = 199;
    exp_55_ram[134] = 231;
    exp_55_ram[135] = 7;
    exp_55_ram[136] = 199;
    exp_55_ram[137] = 23;
    exp_55_ram[138] = 3;
    exp_55_ram[139] = 3;
    exp_55_ram[140] = 23;
    exp_55_ram[141] = 7;
    exp_55_ram[142] = 103;
    exp_55_ram[143] = 230;
    exp_55_ram[144] = 7;
    exp_55_ram[145] = 211;
    exp_55_ram[146] = 104;
    exp_55_ram[147] = 247;
    exp_55_ram[148] = 3;
    exp_55_ram[149] = 211;
    exp_55_ram[150] = 231;
    exp_55_ram[151] = 5;
    exp_55_ram[152] = 197;
    exp_55_ram[153] = 0;
    exp_55_ram[154] = 0;
    exp_55_ram[155] = 0;
    exp_55_ram[156] = 232;
    exp_55_ram[157] = 128;
    exp_55_ram[158] = 31;
    exp_55_ram[159] = 216;
    exp_55_ram[160] = 231;
    exp_55_ram[161] = 216;
    exp_55_ram[162] = 215;
    exp_55_ram[163] = 232;
    exp_55_ram[164] = 8;
    exp_55_ram[165] = 247;
    exp_55_ram[166] = 21;
    exp_55_ram[167] = 8;
    exp_55_ram[168] = 7;
    exp_55_ram[169] = 6;
    exp_55_ram[170] = 21;
    exp_55_ram[171] = 7;
    exp_55_ram[172] = 183;
    exp_55_ram[173] = 167;
    exp_55_ram[174] = 5;
    exp_55_ram[175] = 215;
    exp_55_ram[176] = 7;
    exp_55_ram[177] = 245;
    exp_55_ram[178] = 7;
    exp_55_ram[179] = 215;
    exp_55_ram[180] = 229;
    exp_55_ram[181] = 7;
    exp_55_ram[182] = 215;
    exp_55_ram[183] = 22;
    exp_55_ram[184] = 6;
    exp_55_ram[185] = 6;
    exp_55_ram[186] = 22;
    exp_55_ram[187] = 7;
    exp_55_ram[188] = 215;
    exp_55_ram[189] = 199;
    exp_55_ram[190] = 6;
    exp_55_ram[191] = 167;
    exp_55_ram[192] = 7;
    exp_55_ram[193] = 246;
    exp_55_ram[194] = 7;
    exp_55_ram[195] = 167;
    exp_55_ram[196] = 230;
    exp_55_ram[197] = 7;
    exp_55_ram[198] = 5;
    exp_55_ram[199] = 167;
    exp_55_ram[200] = 229;
    exp_55_ram[201] = 159;
    exp_55_ram[202] = 213;
    exp_55_ram[203] = 1;
    exp_55_ram[204] = 230;
    exp_55_ram[205] = 240;
    exp_55_ram[206] = 215;
    exp_55_ram[207] = 53;
    exp_55_ram[208] = 0;
    exp_55_ram[209] = 182;
    exp_55_ram[210] = 71;
    exp_55_ram[211] = 167;
    exp_55_ram[212] = 7;
    exp_55_ram[213] = 0;
    exp_55_ram[214] = 183;
    exp_55_ram[215] = 229;
    exp_55_ram[216] = 229;
    exp_55_ram[217] = 16;
    exp_55_ram[218] = 246;
    exp_55_ram[219] = 200;
    exp_55_ram[220] = 21;
    exp_55_ram[221] = 31;
    exp_55_ram[222] = 0;
    exp_55_ram[223] = 0;
    exp_55_ram[224] = 230;
    exp_55_ram[225] = 128;
    exp_55_ram[226] = 159;
    exp_55_ram[227] = 230;
    exp_55_ram[228] = 182;
    exp_55_ram[229] = 216;
    exp_55_ram[230] = 231;
    exp_55_ram[231] = 8;
    exp_55_ram[232] = 222;
    exp_55_ram[233] = 183;
    exp_55_ram[234] = 232;
    exp_55_ram[235] = 182;
    exp_55_ram[236] = 247;
    exp_55_ram[237] = 8;
    exp_55_ram[238] = 7;
    exp_55_ram[239] = 6;
    exp_55_ram[240] = 222;
    exp_55_ram[241] = 6;
    exp_55_ram[242] = 230;
    exp_55_ram[243] = 199;
    exp_55_ram[244] = 14;
    exp_55_ram[245] = 231;
    exp_55_ram[246] = 7;
    exp_55_ram[247] = 254;
    exp_55_ram[248] = 7;
    exp_55_ram[249] = 231;
    exp_55_ram[250] = 238;
    exp_55_ram[251] = 7;
    exp_55_ram[252] = 231;
    exp_55_ram[253] = 215;
    exp_55_ram[254] = 215;
    exp_55_ram[255] = 6;
    exp_55_ram[256] = 231;
    exp_55_ram[257] = 6;
    exp_55_ram[258] = 7;
    exp_55_ram[259] = 246;
    exp_55_ram[260] = 7;
    exp_55_ram[261] = 199;
    exp_55_ram[262] = 7;
    exp_55_ram[263] = 247;
    exp_55_ram[264] = 7;
    exp_55_ram[265] = 199;
    exp_55_ram[266] = 231;
    exp_55_ram[267] = 7;
    exp_55_ram[268] = 5;
    exp_55_ram[269] = 1;
    exp_55_ram[270] = 197;
    exp_55_ram[271] = 254;
    exp_55_ram[272] = 213;
    exp_55_ram[273] = 5;
    exp_55_ram[274] = 211;
    exp_55_ram[275] = 3;
    exp_55_ram[276] = 199;
    exp_55_ram[277] = 216;
    exp_55_ram[278] = 214;
    exp_55_ram[279] = 14;
    exp_55_ram[280] = 104;
    exp_55_ram[281] = 216;
    exp_55_ram[282] = 7;
    exp_55_ram[283] = 102;
    exp_55_ram[284] = 215;
    exp_55_ram[285] = 214;
    exp_55_ram[286] = 7;
    exp_55_ram[287] = 198;
    exp_55_ram[288] = 199;
    exp_55_ram[289] = 199;
    exp_55_ram[290] = 1;
    exp_55_ram[291] = 247;
    exp_55_ram[292] = 247;
    exp_55_ram[293] = 7;
    exp_55_ram[294] = 254;
    exp_55_ram[295] = 184;
    exp_55_ram[296] = 199;
    exp_55_ram[297] = 0;
    exp_55_ram[298] = 232;
    exp_55_ram[299] = 245;
    exp_55_ram[300] = 223;
    exp_55_ram[301] = 0;
    exp_55_ram[302] = 0;
    exp_55_ram[303] = 159;
    exp_55_ram[304] = 16;
    exp_55_ram[305] = 247;
    exp_55_ram[306] = 69;
    exp_55_ram[307] = 183;
    exp_55_ram[308] = 5;
    exp_55_ram[309] = 5;
    exp_55_ram[310] = 248;
    exp_55_ram[311] = 245;
    exp_55_ram[312] = 240;
    exp_55_ram[313] = 70;
    exp_55_ram[314] = 215;
    exp_55_ram[315] = 6;
    exp_55_ram[316] = 245;
    exp_55_ram[317] = 246;
    exp_55_ram[318] = 216;
    exp_55_ram[319] = 248;
    exp_55_ram[320] = 14;
    exp_55_ram[321] = 32;
    exp_55_ram[322] = 0;
    exp_55_ram[323] = 213;
    exp_55_ram[324] = 199;
    exp_55_ram[325] = 14;
    exp_55_ram[326] = 8;
    exp_55_ram[327] = 248;
    exp_55_ram[328] = 23;
    exp_55_ram[329] = 5;
    exp_55_ram[330] = 199;
    exp_55_ram[331] = 6;
    exp_55_ram[332] = 7;
    exp_55_ram[333] = 213;
    exp_55_ram[334] = 5;
    exp_55_ram[335] = 5;
    exp_55_ram[336] = 240;
    exp_55_ram[337] = 0;
    exp_55_ram[338] = 240;
    exp_55_ram[339] = 6;
    exp_55_ram[340] = 6;
    exp_55_ram[341] = 0;
    exp_55_ram[342] = 184;
    exp_55_ram[343] = 5;
    exp_55_ram[344] = 0;
    exp_55_ram[345] = 23;
    exp_55_ram[346] = 232;
    exp_55_ram[347] = 110;
    exp_55_ram[348] = 195;
    exp_55_ram[349] = 0;
    exp_55_ram[350] = 0;
    exp_55_ram[351] = 16;
    exp_55_ram[352] = 0;
    exp_55_ram[353] = 7;
    exp_55_ram[354] = 95;
    exp_55_ram[355] = 232;
    exp_55_ram[356] = 95;
    exp_55_ram[357] = 5;
    exp_55_ram[358] = 5;
    exp_55_ram[359] = 0;
    exp_55_ram[360] = 159;
    exp_55_ram[361] = 1;
    exp_55_ram[362] = 129;
    exp_55_ram[363] = 17;
    exp_55_ram[364] = 5;
    exp_55_ram[365] = 5;
    exp_55_ram[366] = 64;
    exp_55_ram[367] = 224;
    exp_55_ram[368] = 160;
    exp_55_ram[369] = 167;
    exp_55_ram[370] = 167;
    exp_55_ram[371] = 176;
    exp_55_ram[372] = 167;
    exp_55_ram[373] = 85;
    exp_55_ram[374] = 244;
    exp_55_ram[375] = 164;
    exp_55_ram[376] = 193;
    exp_55_ram[377] = 4;
    exp_55_ram[378] = 199;
    exp_55_ram[379] = 129;
    exp_55_ram[380] = 71;
    exp_55_ram[381] = 199;
    exp_55_ram[382] = 247;
    exp_55_ram[383] = 6;
    exp_55_ram[384] = 1;
    exp_55_ram[385] = 0;
    exp_55_ram[386] = 85;
    exp_55_ram[387] = 244;
    exp_55_ram[388] = 0;
    exp_55_ram[389] = 223;
    exp_55_ram[390] = 0;
    exp_55_ram[391] = 0;
    exp_55_ram[392] = 31;
    exp_55_ram[393] = 1;
    exp_55_ram[394] = 17;
    exp_55_ram[395] = 129;
    exp_55_ram[396] = 145;
    exp_55_ram[397] = 33;
    exp_55_ram[398] = 49;
    exp_55_ram[399] = 65;
    exp_55_ram[400] = 181;
    exp_55_ram[401] = 7;
    exp_55_ram[402] = 5;
    exp_55_ram[403] = 5;
    exp_55_ram[404] = 5;
    exp_55_ram[405] = 5;
    exp_55_ram[406] = 5;
    exp_55_ram[407] = 0;
    exp_55_ram[408] = 5;
    exp_55_ram[409] = 224;
    exp_55_ram[410] = 58;
    exp_55_ram[411] = 48;
    exp_55_ram[412] = 71;
    exp_55_ram[413] = 176;
    exp_55_ram[414] = 4;
    exp_55_ram[415] = 55;
    exp_55_ram[416] = 160;
    exp_55_ram[417] = 55;
    exp_55_ram[418] = 176;
    exp_55_ram[419] = 89;
    exp_55_ram[420] = 52;
    exp_55_ram[421] = 148;
    exp_55_ram[422] = 233;
    exp_55_ram[423] = 180;
    exp_55_ram[424] = 228;
    exp_55_ram[425] = 193;
    exp_55_ram[426] = 129;
    exp_55_ram[427] = 196;
    exp_55_ram[428] = 74;
    exp_55_ram[429] = 197;
    exp_55_ram[430] = 186;
    exp_55_ram[431] = 65;
    exp_55_ram[432] = 1;
    exp_55_ram[433] = 193;
    exp_55_ram[434] = 129;
    exp_55_ram[435] = 7;
    exp_55_ram[436] = 7;
    exp_55_ram[437] = 1;
    exp_55_ram[438] = 0;
    exp_55_ram[439] = 0;
    exp_55_ram[440] = 5;
    exp_55_ram[441] = 31;
    exp_55_ram[442] = 89;
    exp_55_ram[443] = 180;
    exp_55_ram[444] = 0;
    exp_55_ram[445] = 31;
    exp_55_ram[446] = 96;
    exp_55_ram[447] = 71;
    exp_55_ram[448] = 137;
    exp_55_ram[449] = 4;
    exp_55_ram[450] = 9;
    exp_55_ram[451] = 128;
    exp_55_ram[452] = 181;
    exp_55_ram[453] = 128;
    exp_55_ram[454] = 160;
    exp_55_ram[455] = 9;
    exp_55_ram[456] = 4;
    exp_55_ram[457] = 54;
    exp_55_ram[458] = 64;
    exp_55_ram[459] = 164;
    exp_55_ram[460] = 5;
    exp_55_ram[461] = 128;
    exp_55_ram[462] = 4;
    exp_55_ram[463] = 9;
    exp_55_ram[464] = 55;
    exp_55_ram[465] = 112;
    exp_55_ram[466] = 55;
    exp_55_ram[467] = 137;
    exp_55_ram[468] = 233;
    exp_55_ram[469] = 128;
    exp_55_ram[470] = 57;
    exp_55_ram[471] = 36;
    exp_55_ram[472] = 185;
    exp_55_ram[473] = 228;
    exp_55_ram[474] = 128;
    exp_55_ram[475] = 247;
    exp_55_ram[476] = 229;
    exp_55_ram[477] = 119;
    exp_55_ram[478] = 7;
    exp_55_ram[479] = 247;
    exp_55_ram[480] = 64;
    exp_55_ram[481] = 215;
    exp_55_ram[482] = 71;
    exp_55_ram[483] = 247;
    exp_55_ram[484] = 245;
    exp_55_ram[485] = 7;
    exp_55_ram[486] = 128;
    exp_55_ram[487] = 229;
    exp_55_ram[488] = 7;
    exp_55_ram[489] = 128;
    exp_55_ram[490] = 247;
    exp_55_ram[491] = 240;
    exp_55_ram[492] = 229;
    exp_55_ram[493] = 58;
    exp_55_ram[494] = 55;
    exp_55_ram[495] = 213;
    exp_55_ram[496] = 245;
    exp_55_ram[497] = 53;
    exp_55_ram[498] = 223;
    exp_55_ram[499] = 137;
    exp_55_ram[500] = 180;
    exp_55_ram[501] = 0;
    exp_55_ram[502] = 31;
    exp_55_ram[503] = 0;
    exp_55_ram[504] = 0;
    exp_55_ram[505] = 0;
    exp_55_ram[506] = 223;
    exp_55_ram[507] = 6;
    exp_55_ram[508] = 0;
    exp_55_ram[509] = 199;
    exp_55_ram[510] = 240;
    exp_55_ram[511] = 6;
    exp_55_ram[512] = 0;
    exp_55_ram[513] = 165;
    exp_55_ram[514] = 7;
    exp_55_ram[515] = 0;
    exp_55_ram[516] = 197;
    exp_55_ram[517] = 197;
    exp_55_ram[518] = 245;
    exp_55_ram[519] = 181;
    exp_55_ram[520] = 159;
    exp_55_ram[521] = 6;
    exp_55_ram[522] = 0;
    exp_55_ram[523] = 199;
    exp_55_ram[524] = 240;
    exp_55_ram[525] = 6;
    exp_55_ram[526] = 0;
    exp_55_ram[527] = 181;
    exp_55_ram[528] = 7;
    exp_55_ram[529] = 0;
    exp_55_ram[530] = 197;
    exp_55_ram[531] = 197;
    exp_55_ram[532] = 245;
    exp_55_ram[533] = 165;
    exp_55_ram[534] = 159;
    exp_55_ram[535] = 1;
    exp_55_ram[536] = 245;
    exp_55_ram[537] = 240;
    exp_55_ram[538] = 167;
    exp_55_ram[539] = 55;
    exp_55_ram[540] = 0;
    exp_55_ram[541] = 0;
    exp_55_ram[542] = 246;
    exp_55_ram[543] = 245;
    exp_55_ram[544] = 71;
    exp_55_ram[545] = 167;
    exp_55_ram[546] = 5;
    exp_55_ram[547] = 166;
    exp_55_ram[548] = 0;
    exp_55_ram[549] = 0;
    exp_55_ram[550] = 0;
    exp_55_ram[551] = 229;
    exp_55_ram[552] = 128;
    exp_55_ram[553] = 223;
    exp_55_ram[554] = 110;
    exp_55_ram[555] = 84;
    exp_55_ram[556] = 101;
    exp_55_ram[557] = 117;
    exp_55_ram[558] = 83;
    exp_55_ram[559] = 0;
    exp_55_ram[560] = 110;
    exp_55_ram[561] = 77;
    exp_55_ram[562] = 112;
    exp_55_ram[563] = 121;
    exp_55_ram[564] = 74;
    exp_55_ram[565] = 117;
    exp_55_ram[566] = 112;
    exp_55_ram[567] = 78;
    exp_55_ram[568] = 101;
    exp_55_ram[569] = 0;
    exp_55_ram[570] = 108;
    exp_55_ram[571] = 87;
    exp_55_ram[572] = 100;
    exp_55_ram[573] = 0;
    exp_55_ram[574] = 110;
    exp_55_ram[575] = 103;
    exp_55_ram[576] = 105;
    exp_55_ram[577] = 32;
    exp_55_ram[578] = 101;
    exp_55_ram[579] = 101;
    exp_55_ram[580] = 46;
    exp_55_ram[581] = 0;
    exp_55_ram[582] = 110;
    exp_55_ram[583] = 103;
    exp_55_ram[584] = 77;
    exp_55_ram[585] = 109;
    exp_55_ram[586] = 46;
    exp_55_ram[587] = 50;
    exp_55_ram[588] = 116;
    exp_55_ram[589] = 116;
    exp_55_ram[590] = 114;
    exp_55_ram[591] = 108;
    exp_55_ram[592] = 108;
    exp_55_ram[593] = 32;
    exp_55_ram[594] = 49;
    exp_55_ram[595] = 99;
    exp_55_ram[596] = 0;
    exp_55_ram[597] = 52;
    exp_55_ram[598] = 116;
    exp_55_ram[599] = 116;
    exp_55_ram[600] = 114;
    exp_55_ram[601] = 108;
    exp_55_ram[602] = 108;
    exp_55_ram[603] = 32;
    exp_55_ram[604] = 49;
    exp_55_ram[605] = 99;
    exp_55_ram[606] = 0;
    exp_55_ram[607] = 50;
    exp_55_ram[608] = 116;
    exp_55_ram[609] = 116;
    exp_55_ram[610] = 114;
    exp_55_ram[611] = 118;
    exp_55_ram[612] = 115;
    exp_55_ram[613] = 32;
    exp_55_ram[614] = 101;
    exp_55_ram[615] = 100;
    exp_55_ram[616] = 52;
    exp_55_ram[617] = 116;
    exp_55_ram[618] = 116;
    exp_55_ram[619] = 114;
    exp_55_ram[620] = 118;
    exp_55_ram[621] = 115;
    exp_55_ram[622] = 32;
    exp_55_ram[623] = 101;
    exp_55_ram[624] = 100;
    exp_55_ram[625] = 97;
    exp_55_ram[626] = 0;
    exp_55_ram[627] = 110;
    exp_55_ram[628] = 0;
    exp_55_ram[629] = 121;
    exp_55_ram[630] = 0;
    exp_55_ram[631] = 117;
    exp_55_ram[632] = 0;
    exp_55_ram[633] = 110;
    exp_55_ram[634] = 58;
    exp_55_ram[635] = 104;
    exp_55_ram[636] = 45;
    exp_55_ram[637] = 101;
    exp_55_ram[638] = 0;
    exp_55_ram[639] = 41;
    exp_55_ram[640] = 108;
    exp_55_ram[641] = 87;
    exp_55_ram[642] = 100;
    exp_55_ram[643] = 32;
    exp_55_ram[644] = 103;
    exp_55_ram[645] = 82;
    exp_55_ram[646] = 114;
    exp_55_ram[647] = 32;
    exp_55_ram[648] = 116;
    exp_55_ram[649] = 108;
    exp_55_ram[650] = 108;
    exp_55_ram[651] = 116;
    exp_55_ram[652] = 0;
    exp_55_ram[653] = 32;
    exp_55_ram[654] = 108;
    exp_55_ram[655] = 111;
    exp_55_ram[656] = 0;
    exp_55_ram[657] = 32;
    exp_55_ram[658] = 103;
    exp_55_ram[659] = 77;
    exp_55_ram[660] = 105;
    exp_55_ram[661] = 0;
    exp_55_ram[662] = 32;
    exp_55_ram[663] = 32;
    exp_55_ram[664] = 111;
    exp_55_ram[665] = 116;
    exp_55_ram[666] = 112;
    exp_55_ram[667] = 116;
    exp_55_ram[668] = 115;
    exp_55_ram[669] = 0;
    exp_55_ram[670] = 0;
    exp_55_ram[671] = 105;
    exp_55_ram[672] = 32;
    exp_55_ram[673] = 104;
    exp_55_ram[674] = 10;
    exp_55_ram[675] = 61;
    exp_55_ram[676] = 61;
    exp_55_ram[677] = 61;
    exp_55_ram[678] = 10;
    exp_55_ram[679] = 0;
    exp_55_ram[680] = 32;
    exp_55_ram[681] = 101;
    exp_55_ram[682] = 101;
    exp_55_ram[683] = 110;
    exp_55_ram[684] = 40;
    exp_55_ram[685] = 122;
    exp_55_ram[686] = 97;
    exp_55_ram[687] = 32;
    exp_55_ram[688] = 62;
    exp_55_ram[689] = 108;
    exp_55_ram[690] = 44;
    exp_55_ram[691] = 100;
    exp_55_ram[692] = 44;
    exp_55_ram[693] = 103;
    exp_55_ram[694] = 101;
    exp_55_ram[695] = 32;
    exp_55_ram[696] = 10;
    exp_55_ram[697] = 32;
    exp_55_ram[698] = 108;
    exp_55_ram[699] = 111;
    exp_55_ram[700] = 97;
    exp_55_ram[701] = 41;
    exp_55_ram[702] = 103;
    exp_55_ram[703] = 10;
    exp_55_ram[704] = 32;
    exp_55_ram[705] = 103;
    exp_55_ram[706] = 116;
    exp_55_ram[707] = 103;
    exp_55_ram[708] = 82;
    exp_55_ram[709] = 115;
    exp_55_ram[710] = 108;
    exp_55_ram[711] = 41;
    exp_55_ram[712] = 45;
    exp_55_ram[713] = 32;
    exp_55_ram[714] = 116;
    exp_55_ram[715] = 105;
    exp_55_ram[716] = 101;
    exp_55_ram[717] = 105;
    exp_55_ram[718] = 32;
    exp_55_ram[719] = 46;
    exp_55_ram[720] = 97;
    exp_55_ram[721] = 0;
    exp_55_ram[722] = 32;
    exp_55_ram[723] = 111;
    exp_55_ram[724] = 111;
    exp_55_ram[725] = 105;
    exp_55_ram[726] = 32;
    exp_55_ram[727] = 62;
    exp_55_ram[728] = 108;
    exp_55_ram[729] = 44;
    exp_55_ram[730] = 100;
    exp_55_ram[731] = 44;
    exp_55_ram[732] = 103;
    exp_55_ram[733] = 101;
    exp_55_ram[734] = 32;
    exp_55_ram[735] = 10;
    exp_55_ram[736] = 97;
    exp_55_ram[737] = 46;
    exp_55_ram[738] = 0;
    exp_55_ram[739] = 0;
    exp_55_ram[740] = 10;
    exp_55_ram[741] = 2;
    exp_55_ram[742] = 3;
    exp_55_ram[743] = 4;
    exp_55_ram[744] = 4;
    exp_55_ram[745] = 5;
    exp_55_ram[746] = 5;
    exp_55_ram[747] = 5;
    exp_55_ram[748] = 5;
    exp_55_ram[749] = 6;
    exp_55_ram[750] = 6;
    exp_55_ram[751] = 6;
    exp_55_ram[752] = 6;
    exp_55_ram[753] = 6;
    exp_55_ram[754] = 6;
    exp_55_ram[755] = 6;
    exp_55_ram[756] = 6;
    exp_55_ram[757] = 7;
    exp_55_ram[758] = 7;
    exp_55_ram[759] = 7;
    exp_55_ram[760] = 7;
    exp_55_ram[761] = 7;
    exp_55_ram[762] = 7;
    exp_55_ram[763] = 7;
    exp_55_ram[764] = 7;
    exp_55_ram[765] = 7;
    exp_55_ram[766] = 7;
    exp_55_ram[767] = 7;
    exp_55_ram[768] = 7;
    exp_55_ram[769] = 7;
    exp_55_ram[770] = 7;
    exp_55_ram[771] = 7;
    exp_55_ram[772] = 7;
    exp_55_ram[773] = 8;
    exp_55_ram[774] = 8;
    exp_55_ram[775] = 8;
    exp_55_ram[776] = 8;
    exp_55_ram[777] = 8;
    exp_55_ram[778] = 8;
    exp_55_ram[779] = 8;
    exp_55_ram[780] = 8;
    exp_55_ram[781] = 8;
    exp_55_ram[782] = 8;
    exp_55_ram[783] = 8;
    exp_55_ram[784] = 8;
    exp_55_ram[785] = 8;
    exp_55_ram[786] = 8;
    exp_55_ram[787] = 8;
    exp_55_ram[788] = 8;
    exp_55_ram[789] = 8;
    exp_55_ram[790] = 8;
    exp_55_ram[791] = 8;
    exp_55_ram[792] = 8;
    exp_55_ram[793] = 8;
    exp_55_ram[794] = 8;
    exp_55_ram[795] = 8;
    exp_55_ram[796] = 8;
    exp_55_ram[797] = 8;
    exp_55_ram[798] = 8;
    exp_55_ram[799] = 8;
    exp_55_ram[800] = 8;
    exp_55_ram[801] = 8;
    exp_55_ram[802] = 8;
    exp_55_ram[803] = 8;
    exp_55_ram[804] = 8;
    exp_55_ram[805] = 1;
    exp_55_ram[806] = 129;
    exp_55_ram[807] = 1;
    exp_55_ram[808] = 164;
    exp_55_ram[809] = 196;
    exp_55_ram[810] = 244;
    exp_55_ram[811] = 196;
    exp_55_ram[812] = 7;
    exp_55_ram[813] = 7;
    exp_55_ram[814] = 193;
    exp_55_ram[815] = 1;
    exp_55_ram[816] = 0;
    exp_55_ram[817] = 1;
    exp_55_ram[818] = 129;
    exp_55_ram[819] = 1;
    exp_55_ram[820] = 164;
    exp_55_ram[821] = 180;
    exp_55_ram[822] = 132;
    exp_55_ram[823] = 244;
    exp_55_ram[824] = 196;
    exp_55_ram[825] = 196;
    exp_55_ram[826] = 231;
    exp_55_ram[827] = 196;
    exp_55_ram[828] = 7;
    exp_55_ram[829] = 193;
    exp_55_ram[830] = 1;
    exp_55_ram[831] = 0;
    exp_55_ram[832] = 1;
    exp_55_ram[833] = 17;
    exp_55_ram[834] = 129;
    exp_55_ram[835] = 1;
    exp_55_ram[836] = 164;
    exp_55_ram[837] = 0;
    exp_55_ram[838] = 7;
    exp_55_ram[839] = 7;
    exp_55_ram[840] = 196;
    exp_55_ram[841] = 31;
    exp_55_ram[842] = 5;
    exp_55_ram[843] = 7;
    exp_55_ram[844] = 193;
    exp_55_ram[845] = 129;
    exp_55_ram[846] = 1;
    exp_55_ram[847] = 0;
    exp_55_ram[848] = 1;
    exp_55_ram[849] = 17;
    exp_55_ram[850] = 129;
    exp_55_ram[851] = 1;
    exp_55_ram[852] = 0;
    exp_55_ram[853] = 199;
    exp_55_ram[854] = 7;
    exp_55_ram[855] = 159;
    exp_55_ram[856] = 5;
    exp_55_ram[857] = 7;
    exp_55_ram[858] = 193;
    exp_55_ram[859] = 129;
    exp_55_ram[860] = 1;
    exp_55_ram[861] = 0;
    exp_55_ram[862] = 1;
    exp_55_ram[863] = 17;
    exp_55_ram[864] = 129;
    exp_55_ram[865] = 1;
    exp_55_ram[866] = 164;
    exp_55_ram[867] = 180;
    exp_55_ram[868] = 4;
    exp_55_ram[869] = 128;
    exp_55_ram[870] = 196;
    exp_55_ram[871] = 23;
    exp_55_ram[872] = 228;
    exp_55_ram[873] = 196;
    exp_55_ram[874] = 247;
    exp_55_ram[875] = 7;
    exp_55_ram[876] = 132;
    exp_55_ram[877] = 7;
    exp_55_ram[878] = 223;
    exp_55_ram[879] = 196;
    exp_55_ram[880] = 196;
    exp_55_ram[881] = 247;
    exp_55_ram[882] = 7;
    exp_55_ram[883] = 7;
    exp_55_ram[884] = 196;
    exp_55_ram[885] = 7;
    exp_55_ram[886] = 193;
    exp_55_ram[887] = 129;
    exp_55_ram[888] = 1;
    exp_55_ram[889] = 0;
    exp_55_ram[890] = 1;
    exp_55_ram[891] = 17;
    exp_55_ram[892] = 129;
    exp_55_ram[893] = 1;
    exp_55_ram[894] = 164;
    exp_55_ram[895] = 0;
    exp_55_ram[896] = 7;
    exp_55_ram[897] = 7;
    exp_55_ram[898] = 196;
    exp_55_ram[899] = 223;
    exp_55_ram[900] = 0;
    exp_55_ram[901] = 7;
    exp_55_ram[902] = 7;
    exp_55_ram[903] = 160;
    exp_55_ram[904] = 95;
    exp_55_ram[905] = 0;
    exp_55_ram[906] = 7;
    exp_55_ram[907] = 193;
    exp_55_ram[908] = 129;
    exp_55_ram[909] = 1;
    exp_55_ram[910] = 0;
    exp_55_ram[911] = 1;
    exp_55_ram[912] = 129;
    exp_55_ram[913] = 1;
    exp_55_ram[914] = 164;
    exp_55_ram[915] = 196;
    exp_55_ram[916] = 0;
    exp_55_ram[917] = 231;
    exp_55_ram[918] = 196;
    exp_55_ram[919] = 160;
    exp_55_ram[920] = 231;
    exp_55_ram[921] = 196;
    exp_55_ram[922] = 0;
    exp_55_ram[923] = 231;
    exp_55_ram[924] = 196;
    exp_55_ram[925] = 160;
    exp_55_ram[926] = 231;
    exp_55_ram[927] = 16;
    exp_55_ram[928] = 128;
    exp_55_ram[929] = 0;
    exp_55_ram[930] = 7;
    exp_55_ram[931] = 193;
    exp_55_ram[932] = 1;
    exp_55_ram[933] = 0;
    exp_55_ram[934] = 1;
    exp_55_ram[935] = 129;
    exp_55_ram[936] = 1;
    exp_55_ram[937] = 164;
    exp_55_ram[938] = 196;
    exp_55_ram[939] = 0;
    exp_55_ram[940] = 231;
    exp_55_ram[941] = 196;
    exp_55_ram[942] = 160;
    exp_55_ram[943] = 231;
    exp_55_ram[944] = 16;
    exp_55_ram[945] = 128;
    exp_55_ram[946] = 0;
    exp_55_ram[947] = 7;
    exp_55_ram[948] = 193;
    exp_55_ram[949] = 1;
    exp_55_ram[950] = 0;
    exp_55_ram[951] = 1;
    exp_55_ram[952] = 17;
    exp_55_ram[953] = 129;
    exp_55_ram[954] = 1;
    exp_55_ram[955] = 164;
    exp_55_ram[956] = 196;
    exp_55_ram[957] = 95;
    exp_55_ram[958] = 5;
    exp_55_ram[959] = 7;
    exp_55_ram[960] = 196;
    exp_55_ram[961] = 7;
    exp_55_ram[962] = 128;
    exp_55_ram[963] = 196;
    exp_55_ram[964] = 7;
    exp_55_ram[965] = 193;
    exp_55_ram[966] = 129;
    exp_55_ram[967] = 1;
    exp_55_ram[968] = 0;
    exp_55_ram[969] = 1;
    exp_55_ram[970] = 17;
    exp_55_ram[971] = 129;
    exp_55_ram[972] = 145;
    exp_55_ram[973] = 1;
    exp_55_ram[974] = 5;
    exp_55_ram[975] = 68;
    exp_55_ram[976] = 244;
    exp_55_ram[977] = 144;
    exp_55_ram[978] = 244;
    exp_55_ram[979] = 240;
    exp_55_ram[980] = 244;
    exp_55_ram[981] = 16;
    exp_55_ram[982] = 244;
    exp_55_ram[983] = 4;
    exp_55_ram[984] = 4;
    exp_55_ram[985] = 4;
    exp_55_ram[986] = 68;
    exp_55_ram[987] = 132;
    exp_55_ram[988] = 196;
    exp_55_ram[989] = 4;
    exp_55_ram[990] = 68;
    exp_55_ram[991] = 132;
    exp_55_ram[992] = 196;
    exp_55_ram[993] = 4;
    exp_55_ram[994] = 68;
    exp_55_ram[995] = 100;
    exp_55_ram[996] = 20;
    exp_55_ram[997] = 4;
    exp_55_ram[998] = 164;
    exp_55_ram[999] = 180;
    exp_55_ram[1000] = 196;
    exp_55_ram[1001] = 212;
    exp_55_ram[1002] = 228;
    exp_55_ram[1003] = 244;
    exp_55_ram[1004] = 4;
    exp_55_ram[1005] = 7;
    exp_55_ram[1006] = 64;
    exp_55_ram[1007] = 164;
    exp_55_ram[1008] = 180;
    exp_55_ram[1009] = 68;
    exp_55_ram[1010] = 132;
    exp_55_ram[1011] = 196;
    exp_55_ram[1012] = 7;
    exp_55_ram[1013] = 0;
    exp_55_ram[1014] = 4;
    exp_55_ram[1015] = 196;
    exp_55_ram[1016] = 247;
    exp_55_ram[1017] = 244;
    exp_55_ram[1018] = 68;
    exp_55_ram[1019] = 132;
    exp_55_ram[1020] = 196;
    exp_55_ram[1021] = 4;
    exp_55_ram[1022] = 68;
    exp_55_ram[1023] = 132;
    exp_55_ram[1024] = 196;
    exp_55_ram[1025] = 4;
    exp_55_ram[1026] = 68;
    exp_55_ram[1027] = 100;
    exp_55_ram[1028] = 20;
    exp_55_ram[1029] = 4;
    exp_55_ram[1030] = 164;
    exp_55_ram[1031] = 180;
    exp_55_ram[1032] = 196;
    exp_55_ram[1033] = 212;
    exp_55_ram[1034] = 228;
    exp_55_ram[1035] = 244;
    exp_55_ram[1036] = 4;
    exp_55_ram[1037] = 7;
    exp_55_ram[1038] = 64;
    exp_55_ram[1039] = 164;
    exp_55_ram[1040] = 180;
    exp_55_ram[1041] = 68;
    exp_55_ram[1042] = 244;
    exp_55_ram[1043] = 32;
    exp_55_ram[1044] = 244;
    exp_55_ram[1045] = 240;
    exp_55_ram[1046] = 244;
    exp_55_ram[1047] = 16;
    exp_55_ram[1048] = 244;
    exp_55_ram[1049] = 4;
    exp_55_ram[1050] = 4;
    exp_55_ram[1051] = 4;
    exp_55_ram[1052] = 4;
    exp_55_ram[1053] = 68;
    exp_55_ram[1054] = 132;
    exp_55_ram[1055] = 196;
    exp_55_ram[1056] = 4;
    exp_55_ram[1057] = 68;
    exp_55_ram[1058] = 132;
    exp_55_ram[1059] = 196;
    exp_55_ram[1060] = 4;
    exp_55_ram[1061] = 100;
    exp_55_ram[1062] = 20;
    exp_55_ram[1063] = 4;
    exp_55_ram[1064] = 164;
    exp_55_ram[1065] = 180;
    exp_55_ram[1066] = 196;
    exp_55_ram[1067] = 212;
    exp_55_ram[1068] = 228;
    exp_55_ram[1069] = 244;
    exp_55_ram[1070] = 4;
    exp_55_ram[1071] = 7;
    exp_55_ram[1072] = 192;
    exp_55_ram[1073] = 164;
    exp_55_ram[1074] = 180;
    exp_55_ram[1075] = 4;
    exp_55_ram[1076] = 4;
    exp_55_ram[1077] = 68;
    exp_55_ram[1078] = 7;
    exp_55_ram[1079] = 144;
    exp_55_ram[1080] = 196;
    exp_55_ram[1081] = 132;
    exp_55_ram[1082] = 247;
    exp_55_ram[1083] = 244;
    exp_55_ram[1084] = 4;
    exp_55_ram[1085] = 68;
    exp_55_ram[1086] = 132;
    exp_55_ram[1087] = 196;
    exp_55_ram[1088] = 4;
    exp_55_ram[1089] = 68;
    exp_55_ram[1090] = 132;
    exp_55_ram[1091] = 196;
    exp_55_ram[1092] = 4;
    exp_55_ram[1093] = 100;
    exp_55_ram[1094] = 20;
    exp_55_ram[1095] = 4;
    exp_55_ram[1096] = 164;
    exp_55_ram[1097] = 180;
    exp_55_ram[1098] = 196;
    exp_55_ram[1099] = 212;
    exp_55_ram[1100] = 228;
    exp_55_ram[1101] = 244;
    exp_55_ram[1102] = 4;
    exp_55_ram[1103] = 7;
    exp_55_ram[1104] = 192;
    exp_55_ram[1105] = 164;
    exp_55_ram[1106] = 180;
    exp_55_ram[1107] = 4;
    exp_55_ram[1108] = 68;
    exp_55_ram[1109] = 132;
    exp_55_ram[1110] = 196;
    exp_55_ram[1111] = 4;
    exp_55_ram[1112] = 68;
    exp_55_ram[1113] = 132;
    exp_55_ram[1114] = 196;
    exp_55_ram[1115] = 4;
    exp_55_ram[1116] = 100;
    exp_55_ram[1117] = 20;
    exp_55_ram[1118] = 4;
    exp_55_ram[1119] = 164;
    exp_55_ram[1120] = 180;
    exp_55_ram[1121] = 196;
    exp_55_ram[1122] = 212;
    exp_55_ram[1123] = 228;
    exp_55_ram[1124] = 244;
    exp_55_ram[1125] = 4;
    exp_55_ram[1126] = 7;
    exp_55_ram[1127] = 0;
    exp_55_ram[1128] = 164;
    exp_55_ram[1129] = 180;
    exp_55_ram[1130] = 68;
    exp_55_ram[1131] = 196;
    exp_55_ram[1132] = 231;
    exp_55_ram[1133] = 68;
    exp_55_ram[1134] = 196;
    exp_55_ram[1135] = 247;
    exp_55_ram[1136] = 4;
    exp_55_ram[1137] = 132;
    exp_55_ram[1138] = 231;
    exp_55_ram[1139] = 196;
    exp_55_ram[1140] = 196;
    exp_55_ram[1141] = 231;
    exp_55_ram[1142] = 196;
    exp_55_ram[1143] = 196;
    exp_55_ram[1144] = 247;
    exp_55_ram[1145] = 132;
    exp_55_ram[1146] = 132;
    exp_55_ram[1147] = 231;
    exp_55_ram[1148] = 16;
    exp_55_ram[1149] = 128;
    exp_55_ram[1150] = 0;
    exp_55_ram[1151] = 7;
    exp_55_ram[1152] = 193;
    exp_55_ram[1153] = 129;
    exp_55_ram[1154] = 65;
    exp_55_ram[1155] = 1;
    exp_55_ram[1156] = 0;
    exp_55_ram[1157] = 1;
    exp_55_ram[1158] = 17;
    exp_55_ram[1159] = 129;
    exp_55_ram[1160] = 1;
    exp_55_ram[1161] = 164;
    exp_55_ram[1162] = 180;
    exp_55_ram[1163] = 196;
    exp_55_ram[1164] = 132;
    exp_55_ram[1165] = 196;
    exp_55_ram[1166] = 7;
    exp_55_ram[1167] = 144;
    exp_55_ram[1168] = 196;
    exp_55_ram[1169] = 4;
    exp_55_ram[1170] = 68;
    exp_55_ram[1171] = 132;
    exp_55_ram[1172] = 196;
    exp_55_ram[1173] = 4;
    exp_55_ram[1174] = 68;
    exp_55_ram[1175] = 132;
    exp_55_ram[1176] = 196;
    exp_55_ram[1177] = 100;
    exp_55_ram[1178] = 20;
    exp_55_ram[1179] = 4;
    exp_55_ram[1180] = 164;
    exp_55_ram[1181] = 180;
    exp_55_ram[1182] = 196;
    exp_55_ram[1183] = 212;
    exp_55_ram[1184] = 228;
    exp_55_ram[1185] = 244;
    exp_55_ram[1186] = 4;
    exp_55_ram[1187] = 7;
    exp_55_ram[1188] = 95;
    exp_55_ram[1189] = 5;
    exp_55_ram[1190] = 7;
    exp_55_ram[1191] = 193;
    exp_55_ram[1192] = 129;
    exp_55_ram[1193] = 1;
    exp_55_ram[1194] = 0;
    exp_55_ram[1195] = 1;
    exp_55_ram[1196] = 129;
    exp_55_ram[1197] = 1;
    exp_55_ram[1198] = 0;
    exp_55_ram[1199] = 212;
    exp_55_ram[1200] = 0;
    exp_55_ram[1201] = 70;
    exp_55_ram[1202] = 212;
    exp_55_ram[1203] = 132;
    exp_55_ram[1204] = 6;
    exp_55_ram[1205] = 212;
    exp_55_ram[1206] = 4;
    exp_55_ram[1207] = 4;
    exp_55_ram[1208] = 6;
    exp_55_ram[1209] = 212;
    exp_55_ram[1210] = 4;
    exp_55_ram[1211] = 196;
    exp_55_ram[1212] = 6;
    exp_55_ram[1213] = 6;
    exp_55_ram[1214] = 0;
    exp_55_ram[1215] = 4;
    exp_55_ram[1216] = 230;
    exp_55_ram[1217] = 212;
    exp_55_ram[1218] = 68;
    exp_55_ram[1219] = 246;
    exp_55_ram[1220] = 244;
    exp_55_ram[1221] = 4;
    exp_55_ram[1222] = 68;
    exp_55_ram[1223] = 7;
    exp_55_ram[1224] = 7;
    exp_55_ram[1225] = 193;
    exp_55_ram[1226] = 1;
    exp_55_ram[1227] = 0;
    exp_55_ram[1228] = 1;
    exp_55_ram[1229] = 17;
    exp_55_ram[1230] = 129;
    exp_55_ram[1231] = 1;
    exp_55_ram[1232] = 164;
    exp_55_ram[1233] = 180;
    exp_55_ram[1234] = 196;
    exp_55_ram[1235] = 212;
    exp_55_ram[1236] = 132;
    exp_55_ram[1237] = 196;
    exp_55_ram[1238] = 4;
    exp_55_ram[1239] = 68;
    exp_55_ram[1240] = 167;
    exp_55_ram[1241] = 6;
    exp_55_ram[1242] = 7;
    exp_55_ram[1243] = 183;
    exp_55_ram[1244] = 6;
    exp_55_ram[1245] = 7;
    exp_55_ram[1246] = 6;
    exp_55_ram[1247] = 6;
    exp_55_ram[1248] = 7;
    exp_55_ram[1249] = 7;
    exp_55_ram[1250] = 207;
    exp_55_ram[1251] = 5;
    exp_55_ram[1252] = 5;
    exp_55_ram[1253] = 7;
    exp_55_ram[1254] = 7;
    exp_55_ram[1255] = 193;
    exp_55_ram[1256] = 129;
    exp_55_ram[1257] = 1;
    exp_55_ram[1258] = 0;
    exp_55_ram[1259] = 1;
    exp_55_ram[1260] = 129;
    exp_55_ram[1261] = 1;
    exp_55_ram[1262] = 164;
    exp_55_ram[1263] = 196;
    exp_55_ram[1264] = 55;
    exp_55_ram[1265] = 7;
    exp_55_ram[1266] = 196;
    exp_55_ram[1267] = 64;
    exp_55_ram[1268] = 247;
    exp_55_ram[1269] = 7;
    exp_55_ram[1270] = 196;
    exp_55_ram[1271] = 0;
    exp_55_ram[1272] = 247;
    exp_55_ram[1273] = 7;
    exp_55_ram[1274] = 16;
    exp_55_ram[1275] = 128;
    exp_55_ram[1276] = 0;
    exp_55_ram[1277] = 7;
    exp_55_ram[1278] = 193;
    exp_55_ram[1279] = 1;
    exp_55_ram[1280] = 0;
    exp_55_ram[1281] = 1;
    exp_55_ram[1282] = 17;
    exp_55_ram[1283] = 129;
    exp_55_ram[1284] = 1;
    exp_55_ram[1285] = 164;
    exp_55_ram[1286] = 196;
    exp_55_ram[1287] = 31;
    exp_55_ram[1288] = 5;
    exp_55_ram[1289] = 7;
    exp_55_ram[1290] = 224;
    exp_55_ram[1291] = 128;
    exp_55_ram[1292] = 208;
    exp_55_ram[1293] = 7;
    exp_55_ram[1294] = 193;
    exp_55_ram[1295] = 129;
    exp_55_ram[1296] = 1;
    exp_55_ram[1297] = 0;
    exp_55_ram[1298] = 1;
    exp_55_ram[1299] = 17;
    exp_55_ram[1300] = 129;
    exp_55_ram[1301] = 1;
    exp_55_ram[1302] = 164;
    exp_55_ram[1303] = 180;
    exp_55_ram[1304] = 132;
    exp_55_ram[1305] = 48;
    exp_55_ram[1306] = 247;
    exp_55_ram[1307] = 132;
    exp_55_ram[1308] = 128;
    exp_55_ram[1309] = 247;
    exp_55_ram[1310] = 132;
    exp_55_ram[1311] = 80;
    exp_55_ram[1312] = 247;
    exp_55_ram[1313] = 132;
    exp_55_ram[1314] = 160;
    exp_55_ram[1315] = 247;
    exp_55_ram[1316] = 224;
    exp_55_ram[1317] = 64;
    exp_55_ram[1318] = 132;
    exp_55_ram[1319] = 16;
    exp_55_ram[1320] = 247;
    exp_55_ram[1321] = 196;
    exp_55_ram[1322] = 95;
    exp_55_ram[1323] = 5;
    exp_55_ram[1324] = 7;
    exp_55_ram[1325] = 208;
    exp_55_ram[1326] = 0;
    exp_55_ram[1327] = 192;
    exp_55_ram[1328] = 128;
    exp_55_ram[1329] = 240;
    exp_55_ram[1330] = 7;
    exp_55_ram[1331] = 193;
    exp_55_ram[1332] = 129;
    exp_55_ram[1333] = 1;
    exp_55_ram[1334] = 0;
    exp_55_ram[1335] = 1;
    exp_55_ram[1336] = 17;
    exp_55_ram[1337] = 129;
    exp_55_ram[1338] = 145;
    exp_55_ram[1339] = 33;
    exp_55_ram[1340] = 49;
    exp_55_ram[1341] = 65;
    exp_55_ram[1342] = 81;
    exp_55_ram[1343] = 97;
    exp_55_ram[1344] = 113;
    exp_55_ram[1345] = 129;
    exp_55_ram[1346] = 145;
    exp_55_ram[1347] = 161;
    exp_55_ram[1348] = 177;
    exp_55_ram[1349] = 1;
    exp_55_ram[1350] = 5;
    exp_55_ram[1351] = 0;
    exp_55_ram[1352] = 0;
    exp_55_ram[1353] = 244;
    exp_55_ram[1354] = 4;
    exp_55_ram[1355] = 32;
    exp_55_ram[1356] = 244;
    exp_55_ram[1357] = 68;
    exp_55_ram[1358] = 244;
    exp_55_ram[1359] = 196;
    exp_55_ram[1360] = 199;
    exp_55_ram[1361] = 68;
    exp_55_ram[1362] = 247;
    exp_55_ram[1363] = 68;
    exp_55_ram[1364] = 95;
    exp_55_ram[1365] = 5;
    exp_55_ram[1366] = 1;
    exp_55_ram[1367] = 7;
    exp_55_ram[1368] = 247;
    exp_55_ram[1369] = 244;
    exp_55_ram[1370] = 4;
    exp_55_ram[1371] = 132;
    exp_55_ram[1372] = 196;
    exp_55_ram[1373] = 132;
    exp_55_ram[1374] = 196;
    exp_55_ram[1375] = 8;
    exp_55_ram[1376] = 182;
    exp_55_ram[1377] = 7;
    exp_55_ram[1378] = 197;
    exp_55_ram[1379] = 8;
    exp_55_ram[1380] = 166;
    exp_55_ram[1381] = 245;
    exp_55_ram[1382] = 6;
    exp_55_ram[1383] = 228;
    exp_55_ram[1384] = 244;
    exp_55_ram[1385] = 68;
    exp_55_ram[1386] = 23;
    exp_55_ram[1387] = 244;
    exp_55_ram[1388] = 223;
    exp_55_ram[1389] = 0;
    exp_55_ram[1390] = 4;
    exp_55_ram[1391] = 4;
    exp_55_ram[1392] = 7;
    exp_55_ram[1393] = 4;
    exp_55_ram[1394] = 231;
    exp_55_ram[1395] = 4;
    exp_55_ram[1396] = 68;
    exp_55_ram[1397] = 95;
    exp_55_ram[1398] = 5;
    exp_55_ram[1399] = 1;
    exp_55_ram[1400] = 7;
    exp_55_ram[1401] = 247;
    exp_55_ram[1402] = 7;
    exp_55_ram[1403] = 0;
    exp_55_ram[1404] = 132;
    exp_55_ram[1405] = 196;
    exp_55_ram[1406] = 166;
    exp_55_ram[1407] = 7;
    exp_55_ram[1408] = 197;
    exp_55_ram[1409] = 182;
    exp_55_ram[1410] = 245;
    exp_55_ram[1411] = 6;
    exp_55_ram[1412] = 228;
    exp_55_ram[1413] = 244;
    exp_55_ram[1414] = 4;
    exp_55_ram[1415] = 23;
    exp_55_ram[1416] = 244;
    exp_55_ram[1417] = 159;
    exp_55_ram[1418] = 0;
    exp_55_ram[1419] = 196;
    exp_55_ram[1420] = 247;
    exp_55_ram[1421] = 1;
    exp_55_ram[1422] = 7;
    exp_55_ram[1423] = 247;
    exp_55_ram[1424] = 7;
    exp_55_ram[1425] = 247;
    exp_55_ram[1426] = 7;
    exp_55_ram[1427] = 132;
    exp_55_ram[1428] = 196;
    exp_55_ram[1429] = 134;
    exp_55_ram[1430] = 7;
    exp_55_ram[1431] = 197;
    exp_55_ram[1432] = 150;
    exp_55_ram[1433] = 245;
    exp_55_ram[1434] = 6;
    exp_55_ram[1435] = 228;
    exp_55_ram[1436] = 244;
    exp_55_ram[1437] = 132;
    exp_55_ram[1438] = 0;
    exp_55_ram[1439] = 7;
    exp_55_ram[1440] = 247;
    exp_55_ram[1441] = 7;
    exp_55_ram[1442] = 247;
    exp_55_ram[1443] = 7;
    exp_55_ram[1444] = 132;
    exp_55_ram[1445] = 196;
    exp_55_ram[1446] = 102;
    exp_55_ram[1447] = 7;
    exp_55_ram[1448] = 197;
    exp_55_ram[1449] = 118;
    exp_55_ram[1450] = 245;
    exp_55_ram[1451] = 6;
    exp_55_ram[1452] = 228;
    exp_55_ram[1453] = 244;
    exp_55_ram[1454] = 68;
    exp_55_ram[1455] = 7;
    exp_55_ram[1456] = 71;
    exp_55_ram[1457] = 231;
    exp_55_ram[1458] = 39;
    exp_55_ram[1459] = 7;
    exp_55_ram[1460] = 247;
    exp_55_ram[1461] = 7;
    exp_55_ram[1462] = 132;
    exp_55_ram[1463] = 196;
    exp_55_ram[1464] = 70;
    exp_55_ram[1465] = 7;
    exp_55_ram[1466] = 197;
    exp_55_ram[1467] = 86;
    exp_55_ram[1468] = 245;
    exp_55_ram[1469] = 6;
    exp_55_ram[1470] = 228;
    exp_55_ram[1471] = 244;
    exp_55_ram[1472] = 4;
    exp_55_ram[1473] = 7;
    exp_55_ram[1474] = 247;
    exp_55_ram[1475] = 7;
    exp_55_ram[1476] = 132;
    exp_55_ram[1477] = 196;
    exp_55_ram[1478] = 38;
    exp_55_ram[1479] = 7;
    exp_55_ram[1480] = 197;
    exp_55_ram[1481] = 54;
    exp_55_ram[1482] = 245;
    exp_55_ram[1483] = 6;
    exp_55_ram[1484] = 228;
    exp_55_ram[1485] = 244;
    exp_55_ram[1486] = 132;
    exp_55_ram[1487] = 196;
    exp_55_ram[1488] = 7;
    exp_55_ram[1489] = 7;
    exp_55_ram[1490] = 193;
    exp_55_ram[1491] = 129;
    exp_55_ram[1492] = 65;
    exp_55_ram[1493] = 1;
    exp_55_ram[1494] = 193;
    exp_55_ram[1495] = 129;
    exp_55_ram[1496] = 65;
    exp_55_ram[1497] = 1;
    exp_55_ram[1498] = 193;
    exp_55_ram[1499] = 129;
    exp_55_ram[1500] = 65;
    exp_55_ram[1501] = 1;
    exp_55_ram[1502] = 193;
    exp_55_ram[1503] = 1;
    exp_55_ram[1504] = 0;
    exp_55_ram[1505] = 1;
    exp_55_ram[1506] = 17;
    exp_55_ram[1507] = 129;
    exp_55_ram[1508] = 145;
    exp_55_ram[1509] = 33;
    exp_55_ram[1510] = 49;
    exp_55_ram[1511] = 1;
    exp_55_ram[1512] = 164;
    exp_55_ram[1513] = 196;
    exp_55_ram[1514] = 7;
    exp_55_ram[1515] = 71;
    exp_55_ram[1516] = 135;
    exp_55_ram[1517] = 199;
    exp_55_ram[1518] = 7;
    exp_55_ram[1519] = 71;
    exp_55_ram[1520] = 135;
    exp_55_ram[1521] = 199;
    exp_55_ram[1522] = 7;
    exp_55_ram[1523] = 100;
    exp_55_ram[1524] = 20;
    exp_55_ram[1525] = 4;
    exp_55_ram[1526] = 164;
    exp_55_ram[1527] = 180;
    exp_55_ram[1528] = 196;
    exp_55_ram[1529] = 212;
    exp_55_ram[1530] = 228;
    exp_55_ram[1531] = 244;
    exp_55_ram[1532] = 196;
    exp_55_ram[1533] = 4;
    exp_55_ram[1534] = 68;
    exp_55_ram[1535] = 132;
    exp_55_ram[1536] = 196;
    exp_55_ram[1537] = 4;
    exp_55_ram[1538] = 68;
    exp_55_ram[1539] = 132;
    exp_55_ram[1540] = 196;
    exp_55_ram[1541] = 100;
    exp_55_ram[1542] = 20;
    exp_55_ram[1543] = 4;
    exp_55_ram[1544] = 164;
    exp_55_ram[1545] = 180;
    exp_55_ram[1546] = 196;
    exp_55_ram[1547] = 212;
    exp_55_ram[1548] = 228;
    exp_55_ram[1549] = 244;
    exp_55_ram[1550] = 4;
    exp_55_ram[1551] = 7;
    exp_55_ram[1552] = 223;
    exp_55_ram[1553] = 164;
    exp_55_ram[1554] = 180;
    exp_55_ram[1555] = 196;
    exp_55_ram[1556] = 240;
    exp_55_ram[1557] = 4;
    exp_55_ram[1558] = 68;
    exp_55_ram[1559] = 255;
    exp_55_ram[1560] = 5;
    exp_55_ram[1561] = 240;
    exp_55_ram[1562] = 166;
    exp_55_ram[1563] = 7;
    exp_55_ram[1564] = 200;
    exp_55_ram[1565] = 182;
    exp_55_ram[1566] = 248;
    exp_55_ram[1567] = 6;
    exp_55_ram[1568] = 228;
    exp_55_ram[1569] = 244;
    exp_55_ram[1570] = 192;
    exp_55_ram[1571] = 196;
    exp_55_ram[1572] = 7;
    exp_55_ram[1573] = 196;
    exp_55_ram[1574] = 4;
    exp_55_ram[1575] = 68;
    exp_55_ram[1576] = 132;
    exp_55_ram[1577] = 196;
    exp_55_ram[1578] = 4;
    exp_55_ram[1579] = 68;
    exp_55_ram[1580] = 132;
    exp_55_ram[1581] = 196;
    exp_55_ram[1582] = 100;
    exp_55_ram[1583] = 20;
    exp_55_ram[1584] = 4;
    exp_55_ram[1585] = 164;
    exp_55_ram[1586] = 180;
    exp_55_ram[1587] = 196;
    exp_55_ram[1588] = 212;
    exp_55_ram[1589] = 228;
    exp_55_ram[1590] = 244;
    exp_55_ram[1591] = 4;
    exp_55_ram[1592] = 7;
    exp_55_ram[1593] = 15;
    exp_55_ram[1594] = 5;
    exp_55_ram[1595] = 7;
    exp_55_ram[1596] = 0;
    exp_55_ram[1597] = 6;
    exp_55_ram[1598] = 0;
    exp_55_ram[1599] = 192;
    exp_55_ram[1600] = 0;
    exp_55_ram[1601] = 0;
    exp_55_ram[1602] = 4;
    exp_55_ram[1603] = 68;
    exp_55_ram[1604] = 197;
    exp_55_ram[1605] = 7;
    exp_55_ram[1606] = 5;
    exp_55_ram[1607] = 213;
    exp_55_ram[1608] = 7;
    exp_55_ram[1609] = 6;
    exp_55_ram[1610] = 228;
    exp_55_ram[1611] = 244;
    exp_55_ram[1612] = 64;
    exp_55_ram[1613] = 4;
    exp_55_ram[1614] = 68;
    exp_55_ram[1615] = 228;
    exp_55_ram[1616] = 244;
    exp_55_ram[1617] = 0;
    exp_55_ram[1618] = 71;
    exp_55_ram[1619] = 7;
    exp_55_ram[1620] = 247;
    exp_55_ram[1621] = 7;
    exp_55_ram[1622] = 132;
    exp_55_ram[1623] = 196;
    exp_55_ram[1624] = 38;
    exp_55_ram[1625] = 7;
    exp_55_ram[1626] = 182;
    exp_55_ram[1627] = 54;
    exp_55_ram[1628] = 183;
    exp_55_ram[1629] = 6;
    exp_55_ram[1630] = 228;
    exp_55_ram[1631] = 244;
    exp_55_ram[1632] = 196;
    exp_55_ram[1633] = 4;
    exp_55_ram[1634] = 132;
    exp_55_ram[1635] = 196;
    exp_55_ram[1636] = 7;
    exp_55_ram[1637] = 0;
    exp_55_ram[1638] = 4;
    exp_55_ram[1639] = 68;
    exp_55_ram[1640] = 132;
    exp_55_ram[1641] = 196;
    exp_55_ram[1642] = 4;
    exp_55_ram[1643] = 68;
    exp_55_ram[1644] = 132;
    exp_55_ram[1645] = 196;
    exp_55_ram[1646] = 4;
    exp_55_ram[1647] = 100;
    exp_55_ram[1648] = 20;
    exp_55_ram[1649] = 4;
    exp_55_ram[1650] = 164;
    exp_55_ram[1651] = 180;
    exp_55_ram[1652] = 196;
    exp_55_ram[1653] = 212;
    exp_55_ram[1654] = 228;
    exp_55_ram[1655] = 244;
    exp_55_ram[1656] = 196;
    exp_55_ram[1657] = 240;
    exp_55_ram[1658] = 196;
    exp_55_ram[1659] = 16;
    exp_55_ram[1660] = 231;
    exp_55_ram[1661] = 128;
    exp_55_ram[1662] = 196;
    exp_55_ram[1663] = 7;
    exp_55_ram[1664] = 196;
    exp_55_ram[1665] = 4;
    exp_55_ram[1666] = 68;
    exp_55_ram[1667] = 132;
    exp_55_ram[1668] = 196;
    exp_55_ram[1669] = 4;
    exp_55_ram[1670] = 68;
    exp_55_ram[1671] = 132;
    exp_55_ram[1672] = 196;
    exp_55_ram[1673] = 100;
    exp_55_ram[1674] = 20;
    exp_55_ram[1675] = 4;
    exp_55_ram[1676] = 164;
    exp_55_ram[1677] = 180;
    exp_55_ram[1678] = 196;
    exp_55_ram[1679] = 212;
    exp_55_ram[1680] = 228;
    exp_55_ram[1681] = 244;
    exp_55_ram[1682] = 4;
    exp_55_ram[1683] = 7;
    exp_55_ram[1684] = 79;
    exp_55_ram[1685] = 5;
    exp_55_ram[1686] = 196;
    exp_55_ram[1687] = 231;
    exp_55_ram[1688] = 192;
    exp_55_ram[1689] = 196;
    exp_55_ram[1690] = 7;
    exp_55_ram[1691] = 132;
    exp_55_ram[1692] = 196;
    exp_55_ram[1693] = 7;
    exp_55_ram[1694] = 7;
    exp_55_ram[1695] = 193;
    exp_55_ram[1696] = 129;
    exp_55_ram[1697] = 65;
    exp_55_ram[1698] = 1;
    exp_55_ram[1699] = 193;
    exp_55_ram[1700] = 1;
    exp_55_ram[1701] = 0;
    exp_55_ram[1702] = 1;
    exp_55_ram[1703] = 17;
    exp_55_ram[1704] = 129;
    exp_55_ram[1705] = 33;
    exp_55_ram[1706] = 49;
    exp_55_ram[1707] = 65;
    exp_55_ram[1708] = 81;
    exp_55_ram[1709] = 97;
    exp_55_ram[1710] = 113;
    exp_55_ram[1711] = 1;
    exp_55_ram[1712] = 164;
    exp_55_ram[1713] = 143;
    exp_55_ram[1714] = 5;
    exp_55_ram[1715] = 5;
    exp_55_ram[1716] = 0;
    exp_55_ram[1717] = 134;
    exp_55_ram[1718] = 6;
    exp_55_ram[1719] = 0;
    exp_55_ram[1720] = 10;
    exp_55_ram[1721] = 10;
    exp_55_ram[1722] = 7;
    exp_55_ram[1723] = 7;
    exp_55_ram[1724] = 207;
    exp_55_ram[1725] = 5;
    exp_55_ram[1726] = 5;
    exp_55_ram[1727] = 228;
    exp_55_ram[1728] = 0;
    exp_55_ram[1729] = 135;
    exp_55_ram[1730] = 199;
    exp_55_ram[1731] = 196;
    exp_55_ram[1732] = 231;
    exp_55_ram[1733] = 244;
    exp_55_ram[1734] = 196;
    exp_55_ram[1735] = 7;
    exp_55_ram[1736] = 196;
    exp_55_ram[1737] = 7;
    exp_55_ram[1738] = 0;
    exp_55_ram[1739] = 196;
    exp_55_ram[1740] = 39;
    exp_55_ram[1741] = 55;
    exp_55_ram[1742] = 196;
    exp_55_ram[1743] = 7;
    exp_55_ram[1744] = 0;
    exp_55_ram[1745] = 11;
    exp_55_ram[1746] = 11;
    exp_55_ram[1747] = 7;
    exp_55_ram[1748] = 7;
    exp_55_ram[1749] = 193;
    exp_55_ram[1750] = 129;
    exp_55_ram[1751] = 65;
    exp_55_ram[1752] = 1;
    exp_55_ram[1753] = 193;
    exp_55_ram[1754] = 129;
    exp_55_ram[1755] = 65;
    exp_55_ram[1756] = 1;
    exp_55_ram[1757] = 1;
    exp_55_ram[1758] = 0;
    exp_55_ram[1759] = 1;
    exp_55_ram[1760] = 17;
    exp_55_ram[1761] = 129;
    exp_55_ram[1762] = 33;
    exp_55_ram[1763] = 49;
    exp_55_ram[1764] = 1;
    exp_55_ram[1765] = 164;
    exp_55_ram[1766] = 180;
    exp_55_ram[1767] = 15;
    exp_55_ram[1768] = 5;
    exp_55_ram[1769] = 5;
    exp_55_ram[1770] = 0;
    exp_55_ram[1771] = 134;
    exp_55_ram[1772] = 6;
    exp_55_ram[1773] = 0;
    exp_55_ram[1774] = 9;
    exp_55_ram[1775] = 9;
    exp_55_ram[1776] = 7;
    exp_55_ram[1777] = 7;
    exp_55_ram[1778] = 79;
    exp_55_ram[1779] = 5;
    exp_55_ram[1780] = 5;
    exp_55_ram[1781] = 228;
    exp_55_ram[1782] = 244;
    exp_55_ram[1783] = 132;
    exp_55_ram[1784] = 196;
    exp_55_ram[1785] = 132;
    exp_55_ram[1786] = 196;
    exp_55_ram[1787] = 167;
    exp_55_ram[1788] = 6;
    exp_55_ram[1789] = 7;
    exp_55_ram[1790] = 183;
    exp_55_ram[1791] = 6;
    exp_55_ram[1792] = 7;
    exp_55_ram[1793] = 6;
    exp_55_ram[1794] = 6;
    exp_55_ram[1795] = 0;
    exp_55_ram[1796] = 230;
    exp_55_ram[1797] = 246;
    exp_55_ram[1798] = 0;
    exp_55_ram[1799] = 193;
    exp_55_ram[1800] = 129;
    exp_55_ram[1801] = 65;
    exp_55_ram[1802] = 1;
    exp_55_ram[1803] = 1;
    exp_55_ram[1804] = 0;
    exp_55_ram[1805] = 1;
    exp_55_ram[1806] = 17;
    exp_55_ram[1807] = 129;
    exp_55_ram[1808] = 1;
    exp_55_ram[1809] = 164;
    exp_55_ram[1810] = 0;
    exp_55_ram[1811] = 135;
    exp_55_ram[1812] = 7;
    exp_55_ram[1813] = 71;
    exp_55_ram[1814] = 135;
    exp_55_ram[1815] = 199;
    exp_55_ram[1816] = 7;
    exp_55_ram[1817] = 164;
    exp_55_ram[1818] = 180;
    exp_55_ram[1819] = 196;
    exp_55_ram[1820] = 212;
    exp_55_ram[1821] = 228;
    exp_55_ram[1822] = 71;
    exp_55_ram[1823] = 244;
    exp_55_ram[1824] = 0;
    exp_55_ram[1825] = 7;
    exp_55_ram[1826] = 7;
    exp_55_ram[1827] = 71;
    exp_55_ram[1828] = 135;
    exp_55_ram[1829] = 199;
    exp_55_ram[1830] = 7;
    exp_55_ram[1831] = 71;
    exp_55_ram[1832] = 135;
    exp_55_ram[1833] = 199;
    exp_55_ram[1834] = 7;
    exp_55_ram[1835] = 196;
    exp_55_ram[1836] = 100;
    exp_55_ram[1837] = 20;
    exp_55_ram[1838] = 4;
    exp_55_ram[1839] = 164;
    exp_55_ram[1840] = 180;
    exp_55_ram[1841] = 196;
    exp_55_ram[1842] = 212;
    exp_55_ram[1843] = 228;
    exp_55_ram[1844] = 71;
    exp_55_ram[1845] = 244;
    exp_55_ram[1846] = 4;
    exp_55_ram[1847] = 192;
    exp_55_ram[1848] = 196;
    exp_55_ram[1849] = 135;
    exp_55_ram[1850] = 7;
    exp_55_ram[1851] = 23;
    exp_55_ram[1852] = 231;
    exp_55_ram[1853] = 196;
    exp_55_ram[1854] = 247;
    exp_55_ram[1855] = 4;
    exp_55_ram[1856] = 247;
    exp_55_ram[1857] = 71;
    exp_55_ram[1858] = 0;
    exp_55_ram[1859] = 7;
    exp_55_ram[1860] = 196;
    exp_55_ram[1861] = 246;
    exp_55_ram[1862] = 231;
    exp_55_ram[1863] = 196;
    exp_55_ram[1864] = 23;
    exp_55_ram[1865] = 244;
    exp_55_ram[1866] = 196;
    exp_55_ram[1867] = 32;
    exp_55_ram[1868] = 231;
    exp_55_ram[1869] = 0;
    exp_55_ram[1870] = 7;
    exp_55_ram[1871] = 0;
    exp_55_ram[1872] = 231;
    exp_55_ram[1873] = 4;
    exp_55_ram[1874] = 0;
    exp_55_ram[1875] = 196;
    exp_55_ram[1876] = 7;
    exp_55_ram[1877] = 7;
    exp_55_ram[1878] = 23;
    exp_55_ram[1879] = 231;
    exp_55_ram[1880] = 196;
    exp_55_ram[1881] = 247;
    exp_55_ram[1882] = 196;
    exp_55_ram[1883] = 71;
    exp_55_ram[1884] = 4;
    exp_55_ram[1885] = 230;
    exp_55_ram[1886] = 199;
    exp_55_ram[1887] = 0;
    exp_55_ram[1888] = 6;
    exp_55_ram[1889] = 246;
    exp_55_ram[1890] = 231;
    exp_55_ram[1891] = 196;
    exp_55_ram[1892] = 23;
    exp_55_ram[1893] = 244;
    exp_55_ram[1894] = 196;
    exp_55_ram[1895] = 32;
    exp_55_ram[1896] = 231;
    exp_55_ram[1897] = 0;
    exp_55_ram[1898] = 7;
    exp_55_ram[1899] = 0;
    exp_55_ram[1900] = 231;
    exp_55_ram[1901] = 196;
    exp_55_ram[1902] = 199;
    exp_55_ram[1903] = 160;
    exp_55_ram[1904] = 7;
    exp_55_ram[1905] = 128;
    exp_55_ram[1906] = 5;
    exp_55_ram[1907] = 5;
    exp_55_ram[1908] = 228;
    exp_55_ram[1909] = 244;
    exp_55_ram[1910] = 68;
    exp_55_ram[1911] = 247;
    exp_55_ram[1912] = 7;
    exp_55_ram[1913] = 247;
    exp_55_ram[1914] = 0;
    exp_55_ram[1915] = 7;
    exp_55_ram[1916] = 231;
    exp_55_ram[1917] = 132;
    exp_55_ram[1918] = 247;
    exp_55_ram[1919] = 7;
    exp_55_ram[1920] = 247;
    exp_55_ram[1921] = 0;
    exp_55_ram[1922] = 7;
    exp_55_ram[1923] = 231;
    exp_55_ram[1924] = 0;
    exp_55_ram[1925] = 7;
    exp_55_ram[1926] = 0;
    exp_55_ram[1927] = 231;
    exp_55_ram[1928] = 196;
    exp_55_ram[1929] = 135;
    exp_55_ram[1930] = 160;
    exp_55_ram[1931] = 7;
    exp_55_ram[1932] = 192;
    exp_55_ram[1933] = 5;
    exp_55_ram[1934] = 5;
    exp_55_ram[1935] = 228;
    exp_55_ram[1936] = 244;
    exp_55_ram[1937] = 68;
    exp_55_ram[1938] = 247;
    exp_55_ram[1939] = 7;
    exp_55_ram[1940] = 247;
    exp_55_ram[1941] = 0;
    exp_55_ram[1942] = 7;
    exp_55_ram[1943] = 231;
    exp_55_ram[1944] = 132;
    exp_55_ram[1945] = 247;
    exp_55_ram[1946] = 7;
    exp_55_ram[1947] = 247;
    exp_55_ram[1948] = 0;
    exp_55_ram[1949] = 7;
    exp_55_ram[1950] = 231;
    exp_55_ram[1951] = 0;
    exp_55_ram[1952] = 7;
    exp_55_ram[1953] = 160;
    exp_55_ram[1954] = 231;
    exp_55_ram[1955] = 196;
    exp_55_ram[1956] = 71;
    exp_55_ram[1957] = 160;
    exp_55_ram[1958] = 7;
    exp_55_ram[1959] = 0;
    exp_55_ram[1960] = 5;
    exp_55_ram[1961] = 5;
    exp_55_ram[1962] = 228;
    exp_55_ram[1963] = 244;
    exp_55_ram[1964] = 68;
    exp_55_ram[1965] = 247;
    exp_55_ram[1966] = 7;
    exp_55_ram[1967] = 247;
    exp_55_ram[1968] = 0;
    exp_55_ram[1969] = 7;
    exp_55_ram[1970] = 231;
    exp_55_ram[1971] = 132;
    exp_55_ram[1972] = 247;
    exp_55_ram[1973] = 7;
    exp_55_ram[1974] = 247;
    exp_55_ram[1975] = 0;
    exp_55_ram[1976] = 7;
    exp_55_ram[1977] = 231;
    exp_55_ram[1978] = 0;
    exp_55_ram[1979] = 7;
    exp_55_ram[1980] = 160;
    exp_55_ram[1981] = 231;
    exp_55_ram[1982] = 196;
    exp_55_ram[1983] = 7;
    exp_55_ram[1984] = 160;
    exp_55_ram[1985] = 7;
    exp_55_ram[1986] = 80;
    exp_55_ram[1987] = 5;
    exp_55_ram[1988] = 5;
    exp_55_ram[1989] = 228;
    exp_55_ram[1990] = 244;
    exp_55_ram[1991] = 68;
    exp_55_ram[1992] = 247;
    exp_55_ram[1993] = 7;
    exp_55_ram[1994] = 247;
    exp_55_ram[1995] = 0;
    exp_55_ram[1996] = 7;
    exp_55_ram[1997] = 231;
    exp_55_ram[1998] = 132;
    exp_55_ram[1999] = 247;
    exp_55_ram[2000] = 7;
    exp_55_ram[2001] = 247;
    exp_55_ram[2002] = 0;
    exp_55_ram[2003] = 7;
    exp_55_ram[2004] = 231;
    exp_55_ram[2005] = 0;
    exp_55_ram[2006] = 7;
    exp_55_ram[2007] = 0;
    exp_55_ram[2008] = 231;
    exp_55_ram[2009] = 196;
    exp_55_ram[2010] = 71;
    exp_55_ram[2011] = 199;
    exp_55_ram[2012] = 128;
    exp_55_ram[2013] = 7;
    exp_55_ram[2014] = 80;
    exp_55_ram[2015] = 5;
    exp_55_ram[2016] = 5;
    exp_55_ram[2017] = 228;
    exp_55_ram[2018] = 244;
    exp_55_ram[2019] = 68;
    exp_55_ram[2020] = 247;
    exp_55_ram[2021] = 7;
    exp_55_ram[2022] = 247;
    exp_55_ram[2023] = 0;
    exp_55_ram[2024] = 7;
    exp_55_ram[2025] = 231;
    exp_55_ram[2026] = 132;
    exp_55_ram[2027] = 64;
    exp_55_ram[2028] = 7;
    exp_55_ram[2029] = 144;
    exp_55_ram[2030] = 5;
    exp_55_ram[2031] = 5;
    exp_55_ram[2032] = 228;
    exp_55_ram[2033] = 244;
    exp_55_ram[2034] = 68;
    exp_55_ram[2035] = 247;
    exp_55_ram[2036] = 7;
    exp_55_ram[2037] = 247;
    exp_55_ram[2038] = 0;
    exp_55_ram[2039] = 7;
    exp_55_ram[2040] = 231;
    exp_55_ram[2041] = 132;
    exp_55_ram[2042] = 160;
    exp_55_ram[2043] = 7;
    exp_55_ram[2044] = 208;
    exp_55_ram[2045] = 5;
    exp_55_ram[2046] = 5;
    exp_55_ram[2047] = 228;
    exp_55_ram[2048] = 244;
    exp_55_ram[2049] = 68;
    exp_55_ram[2050] = 247;
    exp_55_ram[2051] = 7;
    exp_55_ram[2052] = 247;
    exp_55_ram[2053] = 0;
    exp_55_ram[2054] = 7;
    exp_55_ram[2055] = 231;
    exp_55_ram[2056] = 132;
    exp_55_ram[2057] = 247;
    exp_55_ram[2058] = 7;
    exp_55_ram[2059] = 247;
    exp_55_ram[2060] = 0;
    exp_55_ram[2061] = 7;
    exp_55_ram[2062] = 231;
    exp_55_ram[2063] = 0;
    exp_55_ram[2064] = 7;
    exp_55_ram[2065] = 160;
    exp_55_ram[2066] = 231;
    exp_55_ram[2067] = 0;
    exp_55_ram[2068] = 7;
    exp_55_ram[2069] = 7;
    exp_55_ram[2070] = 0;
    exp_55_ram[2071] = 7;
    exp_55_ram[2072] = 7;
    exp_55_ram[2073] = 193;
    exp_55_ram[2074] = 129;
    exp_55_ram[2075] = 1;
    exp_55_ram[2076] = 0;
    exp_55_ram[2077] = 1;
    exp_55_ram[2078] = 17;
    exp_55_ram[2079] = 129;
    exp_55_ram[2080] = 1;
    exp_55_ram[2081] = 164;
    exp_55_ram[2082] = 196;
    exp_55_ram[2083] = 64;
    exp_55_ram[2084] = 5;
    exp_55_ram[2085] = 7;
    exp_55_ram[2086] = 223;
    exp_55_ram[2087] = 5;
    exp_55_ram[2088] = 7;
    exp_55_ram[2089] = 193;
    exp_55_ram[2090] = 129;
    exp_55_ram[2091] = 1;
    exp_55_ram[2092] = 0;
    exp_55_ram[2093] = 1;
    exp_55_ram[2094] = 17;
    exp_55_ram[2095] = 129;
    exp_55_ram[2096] = 33;
    exp_55_ram[2097] = 49;
    exp_55_ram[2098] = 65;
    exp_55_ram[2099] = 81;
    exp_55_ram[2100] = 97;
    exp_55_ram[2101] = 113;
    exp_55_ram[2102] = 129;
    exp_55_ram[2103] = 145;
    exp_55_ram[2104] = 1;
    exp_55_ram[2105] = 164;
    exp_55_ram[2106] = 180;
    exp_55_ram[2107] = 196;
    exp_55_ram[2108] = 32;
    exp_55_ram[2109] = 244;
    exp_55_ram[2110] = 64;
    exp_55_ram[2111] = 244;
    exp_55_ram[2112] = 132;
    exp_55_ram[2113] = 7;
    exp_55_ram[2114] = 207;
    exp_55_ram[2115] = 164;
    exp_55_ram[2116] = 196;
    exp_55_ram[2117] = 1;
    exp_55_ram[2118] = 7;
    exp_55_ram[2119] = 247;
    exp_55_ram[2120] = 244;
    exp_55_ram[2121] = 132;
    exp_55_ram[2122] = 7;
    exp_55_ram[2123] = 0;
    exp_55_ram[2124] = 68;
    exp_55_ram[2125] = 12;
    exp_55_ram[2126] = 231;
    exp_55_ram[2127] = 68;
    exp_55_ram[2128] = 12;
    exp_55_ram[2129] = 231;
    exp_55_ram[2130] = 4;
    exp_55_ram[2131] = 12;
    exp_55_ram[2132] = 231;
    exp_55_ram[2133] = 132;
    exp_55_ram[2134] = 23;
    exp_55_ram[2135] = 244;
    exp_55_ram[2136] = 196;
    exp_55_ram[2137] = 7;
    exp_55_ram[2138] = 196;
    exp_55_ram[2139] = 247;
    exp_55_ram[2140] = 244;
    exp_55_ram[2141] = 132;
    exp_55_ram[2142] = 7;
    exp_55_ram[2143] = 0;
    exp_55_ram[2144] = 4;
    exp_55_ram[2145] = 68;
    exp_55_ram[2146] = 70;
    exp_55_ram[2147] = 7;
    exp_55_ram[2148] = 182;
    exp_55_ram[2149] = 86;
    exp_55_ram[2150] = 183;
    exp_55_ram[2151] = 6;
    exp_55_ram[2152] = 228;
    exp_55_ram[2153] = 244;
    exp_55_ram[2154] = 159;
    exp_55_ram[2155] = 0;
    exp_55_ram[2156] = 4;
    exp_55_ram[2157] = 4;
    exp_55_ram[2158] = 132;
    exp_55_ram[2159] = 7;
    exp_55_ram[2160] = 68;
    exp_55_ram[2161] = 7;
    exp_55_ram[2162] = 7;
    exp_55_ram[2163] = 207;
    exp_55_ram[2164] = 164;
    exp_55_ram[2165] = 196;
    exp_55_ram[2166] = 1;
    exp_55_ram[2167] = 7;
    exp_55_ram[2168] = 247;
    exp_55_ram[2169] = 244;
    exp_55_ram[2170] = 132;
    exp_55_ram[2171] = 7;
    exp_55_ram[2172] = 0;
    exp_55_ram[2173] = 68;
    exp_55_ram[2174] = 11;
    exp_55_ram[2175] = 231;
    exp_55_ram[2176] = 68;
    exp_55_ram[2177] = 11;
    exp_55_ram[2178] = 231;
    exp_55_ram[2179] = 4;
    exp_55_ram[2180] = 11;
    exp_55_ram[2181] = 231;
    exp_55_ram[2182] = 68;
    exp_55_ram[2183] = 23;
    exp_55_ram[2184] = 244;
    exp_55_ram[2185] = 196;
    exp_55_ram[2186] = 7;
    exp_55_ram[2187] = 196;
    exp_55_ram[2188] = 247;
    exp_55_ram[2189] = 244;
    exp_55_ram[2190] = 4;
    exp_55_ram[2191] = 7;
    exp_55_ram[2192] = 196;
    exp_55_ram[2193] = 247;
    exp_55_ram[2194] = 244;
    exp_55_ram[2195] = 132;
    exp_55_ram[2196] = 7;
    exp_55_ram[2197] = 0;
    exp_55_ram[2198] = 4;
    exp_55_ram[2199] = 68;
    exp_55_ram[2200] = 38;
    exp_55_ram[2201] = 7;
    exp_55_ram[2202] = 182;
    exp_55_ram[2203] = 54;
    exp_55_ram[2204] = 183;
    exp_55_ram[2205] = 6;
    exp_55_ram[2206] = 228;
    exp_55_ram[2207] = 244;
    exp_55_ram[2208] = 159;
    exp_55_ram[2209] = 0;
    exp_55_ram[2210] = 132;
    exp_55_ram[2211] = 71;
    exp_55_ram[2212] = 244;
    exp_55_ram[2213] = 4;
    exp_55_ram[2214] = 1;
    exp_55_ram[2215] = 7;
    exp_55_ram[2216] = 7;
    exp_55_ram[2217] = 144;
    exp_55_ram[2218] = 5;
    exp_55_ram[2219] = 5;
    exp_55_ram[2220] = 228;
    exp_55_ram[2221] = 244;
    exp_55_ram[2222] = 196;
    exp_55_ram[2223] = 23;
    exp_55_ram[2224] = 244;
    exp_55_ram[2225] = 196;
    exp_55_ram[2226] = 196;
    exp_55_ram[2227] = 247;
    exp_55_ram[2228] = 244;
    exp_55_ram[2229] = 196;
    exp_55_ram[2230] = 112;
    exp_55_ram[2231] = 247;
    exp_55_ram[2232] = 244;
    exp_55_ram[2233] = 4;
    exp_55_ram[2234] = 196;
    exp_55_ram[2235] = 247;
    exp_55_ram[2236] = 244;
    exp_55_ram[2237] = 4;
    exp_55_ram[2238] = 244;
    exp_55_ram[2239] = 247;
    exp_55_ram[2240] = 244;
    exp_55_ram[2241] = 4;
    exp_55_ram[2242] = 0;
    exp_55_ram[2243] = 7;
    exp_55_ram[2244] = 7;
    exp_55_ram[2245] = 144;
    exp_55_ram[2246] = 5;
    exp_55_ram[2247] = 5;
    exp_55_ram[2248] = 228;
    exp_55_ram[2249] = 244;
    exp_55_ram[2250] = 196;
    exp_55_ram[2251] = 244;
    exp_55_ram[2252] = 4;
    exp_55_ram[2253] = 244;
    exp_55_ram[2254] = 247;
    exp_55_ram[2255] = 244;
    exp_55_ram[2256] = 4;
    exp_55_ram[2257] = 192;
    exp_55_ram[2258] = 7;
    exp_55_ram[2259] = 16;
    exp_55_ram[2260] = 5;
    exp_55_ram[2261] = 5;
    exp_55_ram[2262] = 228;
    exp_55_ram[2263] = 244;
    exp_55_ram[2264] = 196;
    exp_55_ram[2265] = 244;
    exp_55_ram[2266] = 4;
    exp_55_ram[2267] = 244;
    exp_55_ram[2268] = 247;
    exp_55_ram[2269] = 244;
    exp_55_ram[2270] = 4;
    exp_55_ram[2271] = 244;
    exp_55_ram[2272] = 196;
    exp_55_ram[2273] = 68;
    exp_55_ram[2274] = 132;
    exp_55_ram[2275] = 196;
    exp_55_ram[2276] = 4;
    exp_55_ram[2277] = 68;
    exp_55_ram[2278] = 132;
    exp_55_ram[2279] = 196;
    exp_55_ram[2280] = 4;
    exp_55_ram[2281] = 68;
    exp_55_ram[2282] = 199;
    exp_55_ram[2283] = 103;
    exp_55_ram[2284] = 23;
    exp_55_ram[2285] = 7;
    exp_55_ram[2286] = 167;
    exp_55_ram[2287] = 183;
    exp_55_ram[2288] = 199;
    exp_55_ram[2289] = 215;
    exp_55_ram[2290] = 231;
    exp_55_ram[2291] = 196;
    exp_55_ram[2292] = 193;
    exp_55_ram[2293] = 129;
    exp_55_ram[2294] = 65;
    exp_55_ram[2295] = 1;
    exp_55_ram[2296] = 193;
    exp_55_ram[2297] = 129;
    exp_55_ram[2298] = 65;
    exp_55_ram[2299] = 1;
    exp_55_ram[2300] = 193;
    exp_55_ram[2301] = 129;
    exp_55_ram[2302] = 1;
    exp_55_ram[2303] = 0;
    exp_55_ram[2304] = 1;
    exp_55_ram[2305] = 17;
    exp_55_ram[2306] = 129;
    exp_55_ram[2307] = 145;
    exp_55_ram[2308] = 33;
    exp_55_ram[2309] = 49;
    exp_55_ram[2310] = 1;
    exp_55_ram[2311] = 164;
    exp_55_ram[2312] = 0;
    exp_55_ram[2313] = 0;
    exp_55_ram[2314] = 244;
    exp_55_ram[2315] = 4;
    exp_55_ram[2316] = 196;
    exp_55_ram[2317] = 7;
    exp_55_ram[2318] = 71;
    exp_55_ram[2319] = 228;
    exp_55_ram[2320] = 244;
    exp_55_ram[2321] = 4;
    exp_55_ram[2322] = 68;
    exp_55_ram[2323] = 159;
    exp_55_ram[2324] = 5;
    exp_55_ram[2325] = 7;
    exp_55_ram[2326] = 0;
    exp_55_ram[2327] = 7;
    exp_55_ram[2328] = 0;
    exp_55_ram[2329] = 228;
    exp_55_ram[2330] = 244;
    exp_55_ram[2331] = 0;
    exp_55_ram[2332] = 71;
    exp_55_ram[2333] = 7;
    exp_55_ram[2334] = 247;
    exp_55_ram[2335] = 7;
    exp_55_ram[2336] = 4;
    exp_55_ram[2337] = 68;
    exp_55_ram[2338] = 201;
    exp_55_ram[2339] = 7;
    exp_55_ram[2340] = 37;
    exp_55_ram[2341] = 217;
    exp_55_ram[2342] = 245;
    exp_55_ram[2343] = 6;
    exp_55_ram[2344] = 7;
    exp_55_ram[2345] = 7;
    exp_55_ram[2346] = 132;
    exp_55_ram[2347] = 196;
    exp_55_ram[2348] = 166;
    exp_55_ram[2349] = 7;
    exp_55_ram[2350] = 200;
    exp_55_ram[2351] = 182;
    exp_55_ram[2352] = 248;
    exp_55_ram[2353] = 6;
    exp_55_ram[2354] = 228;
    exp_55_ram[2355] = 244;
    exp_55_ram[2356] = 0;
    exp_55_ram[2357] = 199;
    exp_55_ram[2358] = 4;
    exp_55_ram[2359] = 132;
    exp_55_ram[2360] = 196;
    exp_55_ram[2361] = 7;
    exp_55_ram[2362] = 223;
    exp_55_ram[2363] = 4;
    exp_55_ram[2364] = 68;
    exp_55_ram[2365] = 132;
    exp_55_ram[2366] = 196;
    exp_55_ram[2367] = 4;
    exp_55_ram[2368] = 68;
    exp_55_ram[2369] = 132;
    exp_55_ram[2370] = 196;
    exp_55_ram[2371] = 4;
    exp_55_ram[2372] = 100;
    exp_55_ram[2373] = 20;
    exp_55_ram[2374] = 4;
    exp_55_ram[2375] = 164;
    exp_55_ram[2376] = 180;
    exp_55_ram[2377] = 196;
    exp_55_ram[2378] = 212;
    exp_55_ram[2379] = 228;
    exp_55_ram[2380] = 244;
    exp_55_ram[2381] = 4;
    exp_55_ram[2382] = 68;
    exp_55_ram[2383] = 159;
    exp_55_ram[2384] = 5;
    exp_55_ram[2385] = 0;
    exp_55_ram[2386] = 199;
    exp_55_ram[2387] = 231;
    exp_55_ram[2388] = 0;
    exp_55_ram[2389] = 199;
    exp_55_ram[2390] = 7;
    exp_55_ram[2391] = 193;
    exp_55_ram[2392] = 129;
    exp_55_ram[2393] = 65;
    exp_55_ram[2394] = 1;
    exp_55_ram[2395] = 193;
    exp_55_ram[2396] = 1;
    exp_55_ram[2397] = 0;
    exp_55_ram[2398] = 1;
    exp_55_ram[2399] = 17;
    exp_55_ram[2400] = 129;
    exp_55_ram[2401] = 1;
    exp_55_ram[2402] = 164;
    exp_55_ram[2403] = 4;
    exp_55_ram[2404] = 196;
    exp_55_ram[2405] = 15;
    exp_55_ram[2406] = 5;
    exp_55_ram[2407] = 244;
    exp_55_ram[2408] = 180;
    exp_55_ram[2409] = 7;
    exp_55_ram[2410] = 144;
    exp_55_ram[2411] = 231;
    exp_55_ram[2412] = 196;
    exp_55_ram[2413] = 7;
    exp_55_ram[2414] = 39;
    exp_55_ram[2415] = 231;
    exp_55_ram[2416] = 23;
    exp_55_ram[2417] = 244;
    exp_55_ram[2418] = 180;
    exp_55_ram[2419] = 196;
    exp_55_ram[2420] = 247;
    exp_55_ram[2421] = 7;
    exp_55_ram[2422] = 244;
    exp_55_ram[2423] = 95;
    exp_55_ram[2424] = 0;
    exp_55_ram[2425] = 196;
    exp_55_ram[2426] = 7;
    exp_55_ram[2427] = 193;
    exp_55_ram[2428] = 129;
    exp_55_ram[2429] = 1;
    exp_55_ram[2430] = 0;
    exp_55_ram[2431] = 1;
    exp_55_ram[2432] = 17;
    exp_55_ram[2433] = 129;
    exp_55_ram[2434] = 1;
    exp_55_ram[2435] = 0;
    exp_55_ram[2436] = 199;
    exp_55_ram[2437] = 7;
    exp_55_ram[2438] = 31;
    exp_55_ram[2439] = 5;
    exp_55_ram[2440] = 7;
    exp_55_ram[2441] = 193;
    exp_55_ram[2442] = 129;
    exp_55_ram[2443] = 1;
    exp_55_ram[2444] = 0;
    exp_55_ram[2445] = 1;
    exp_55_ram[2446] = 17;
    exp_55_ram[2447] = 129;
    exp_55_ram[2448] = 1;
    exp_55_ram[2449] = 164;
    exp_55_ram[2450] = 180;
    exp_55_ram[2451] = 196;
    exp_55_ram[2452] = 154;
    exp_55_ram[2453] = 7;
    exp_55_ram[2454] = 244;
    exp_55_ram[2455] = 160;
    exp_55_ram[2456] = 244;
    exp_55_ram[2457] = 4;
    exp_55_ram[2458] = 192;
    exp_55_ram[2459] = 196;
    exp_55_ram[2460] = 196;
    exp_55_ram[2461] = 247;
    exp_55_ram[2462] = 244;
    exp_55_ram[2463] = 52;
    exp_55_ram[2464] = 7;
    exp_55_ram[2465] = 68;
    exp_55_ram[2466] = 7;
    exp_55_ram[2467] = 132;
    exp_55_ram[2468] = 16;
    exp_55_ram[2469] = 247;
    exp_55_ram[2470] = 52;
    exp_55_ram[2471] = 7;
    exp_55_ram[2472] = 68;
    exp_55_ram[2473] = 7;
    exp_55_ram[2474] = 207;
    exp_55_ram[2475] = 16;
    exp_55_ram[2476] = 244;
    exp_55_ram[2477] = 64;
    exp_55_ram[2478] = 132;
    exp_55_ram[2479] = 132;
    exp_55_ram[2480] = 247;
    exp_55_ram[2481] = 52;
    exp_55_ram[2482] = 7;
    exp_55_ram[2483] = 68;
    exp_55_ram[2484] = 7;
    exp_55_ram[2485] = 15;
    exp_55_ram[2486] = 196;
    exp_55_ram[2487] = 196;
    exp_55_ram[2488] = 247;
    exp_55_ram[2489] = 244;
    exp_55_ram[2490] = 196;
    exp_55_ram[2491] = 160;
    exp_55_ram[2492] = 247;
    exp_55_ram[2493] = 244;
    exp_55_ram[2494] = 132;
    exp_55_ram[2495] = 247;
    exp_55_ram[2496] = 244;
    exp_55_ram[2497] = 196;
    exp_55_ram[2498] = 7;
    exp_55_ram[2499] = 0;
    exp_55_ram[2500] = 0;
    exp_55_ram[2501] = 193;
    exp_55_ram[2502] = 129;
    exp_55_ram[2503] = 1;
    exp_55_ram[2504] = 0;
    exp_55_ram[2505] = 1;
    exp_55_ram[2506] = 17;
    exp_55_ram[2507] = 129;
    exp_55_ram[2508] = 1;
    exp_55_ram[2509] = 164;
    exp_55_ram[2510] = 180;
    exp_55_ram[2511] = 196;
    exp_55_ram[2512] = 132;
    exp_55_ram[2513] = 0;
    exp_55_ram[2514] = 7;
    exp_55_ram[2515] = 7;
    exp_55_ram[2516] = 6;
    exp_55_ram[2517] = 7;
    exp_55_ram[2518] = 223;
    exp_55_ram[2519] = 0;
    exp_55_ram[2520] = 193;
    exp_55_ram[2521] = 129;
    exp_55_ram[2522] = 1;
    exp_55_ram[2523] = 0;
    exp_55_ram[2524] = 1;
    exp_55_ram[2525] = 17;
    exp_55_ram[2526] = 129;
    exp_55_ram[2527] = 33;
    exp_55_ram[2528] = 49;
    exp_55_ram[2529] = 1;
    exp_55_ram[2530] = 164;
    exp_55_ram[2531] = 31;
    exp_55_ram[2532] = 164;
    exp_55_ram[2533] = 180;
    exp_55_ram[2534] = 0;
    exp_55_ram[2535] = 31;
    exp_55_ram[2536] = 5;
    exp_55_ram[2537] = 5;
    exp_55_ram[2538] = 132;
    exp_55_ram[2539] = 196;
    exp_55_ram[2540] = 166;
    exp_55_ram[2541] = 7;
    exp_55_ram[2542] = 6;
    exp_55_ram[2543] = 182;
    exp_55_ram[2544] = 7;
    exp_55_ram[2545] = 6;
    exp_55_ram[2546] = 196;
    exp_55_ram[2547] = 6;
    exp_55_ram[2548] = 0;
    exp_55_ram[2549] = 9;
    exp_55_ram[2550] = 7;
    exp_55_ram[2551] = 198;
    exp_55_ram[2552] = 9;
    exp_55_ram[2553] = 7;
    exp_55_ram[2554] = 214;
    exp_55_ram[2555] = 9;
    exp_55_ram[2556] = 7;
    exp_55_ram[2557] = 215;
    exp_55_ram[2558] = 0;
    exp_55_ram[2559] = 7;
    exp_55_ram[2560] = 193;
    exp_55_ram[2561] = 129;
    exp_55_ram[2562] = 65;
    exp_55_ram[2563] = 1;
    exp_55_ram[2564] = 1;
    exp_55_ram[2565] = 0;
    exp_55_ram[2566] = 1;
    exp_55_ram[2567] = 17;
    exp_55_ram[2568] = 129;
    exp_55_ram[2569] = 1;
    exp_55_ram[2570] = 0;
    exp_55_ram[2571] = 135;
    exp_55_ram[2572] = 143;
    exp_55_ram[2573] = 0;
    exp_55_ram[2574] = 193;
    exp_55_ram[2575] = 129;
    exp_55_ram[2576] = 1;
    exp_55_ram[2577] = 0;
    exp_55_ram[2578] = 1;
    exp_55_ram[2579] = 17;
    exp_55_ram[2580] = 129;
    exp_55_ram[2581] = 1;
    exp_55_ram[2582] = 0;
    exp_55_ram[2583] = 135;
    exp_55_ram[2584] = 143;
    exp_55_ram[2585] = 16;
    exp_55_ram[2586] = 244;
    exp_55_ram[2587] = 4;
    exp_55_ram[2588] = 64;
    exp_55_ram[2589] = 0;
    exp_55_ram[2590] = 132;
    exp_55_ram[2591] = 159;
    exp_55_ram[2592] = 160;
    exp_55_ram[2593] = 207;
    exp_55_ram[2594] = 192;
    exp_55_ram[2595] = 196;
    exp_55_ram[2596] = 23;
    exp_55_ram[2597] = 244;
    exp_55_ram[2598] = 0;
    exp_55_ram[2599] = 71;
    exp_55_ram[2600] = 7;
    exp_55_ram[2601] = 196;
    exp_55_ram[2602] = 207;
    exp_55_ram[2603] = 0;
    exp_55_ram[2604] = 135;
    exp_55_ram[2605] = 160;
    exp_55_ram[2606] = 247;
    exp_55_ram[2607] = 7;
    exp_55_ram[2608] = 31;
    exp_55_ram[2609] = 196;
    exp_55_ram[2610] = 240;
    exp_55_ram[2611] = 231;
    exp_55_ram[2612] = 192;
    exp_55_ram[2613] = 196;
    exp_55_ram[2614] = 23;
    exp_55_ram[2615] = 244;
    exp_55_ram[2616] = 0;
    exp_55_ram[2617] = 71;
    exp_55_ram[2618] = 7;
    exp_55_ram[2619] = 196;
    exp_55_ram[2620] = 79;
    exp_55_ram[2621] = 0;
    exp_55_ram[2622] = 135;
    exp_55_ram[2623] = 160;
    exp_55_ram[2624] = 247;
    exp_55_ram[2625] = 7;
    exp_55_ram[2626] = 159;
    exp_55_ram[2627] = 196;
    exp_55_ram[2628] = 16;
    exp_55_ram[2629] = 231;
    exp_55_ram[2630] = 132;
    exp_55_ram[2631] = 23;
    exp_55_ram[2632] = 244;
    exp_55_ram[2633] = 132;
    exp_55_ram[2634] = 144;
    exp_55_ram[2635] = 231;
    exp_55_ram[2636] = 0;
    exp_55_ram[2637] = 71;
    exp_55_ram[2638] = 7;
    exp_55_ram[2639] = 0;
    exp_55_ram[2640] = 79;
    exp_55_ram[2641] = 0;
    exp_55_ram[2642] = 193;
    exp_55_ram[2643] = 129;
    exp_55_ram[2644] = 1;
    exp_55_ram[2645] = 0;
    exp_55_ram[2646] = 1;
    exp_55_ram[2647] = 17;
    exp_55_ram[2648] = 129;
    exp_55_ram[2649] = 1;
    exp_55_ram[2650] = 0;
    exp_55_ram[2651] = 135;
    exp_55_ram[2652] = 143;
    exp_55_ram[2653] = 4;
    exp_55_ram[2654] = 192;
    exp_55_ram[2655] = 0;
    exp_55_ram[2656] = 132;
    exp_55_ram[2657] = 31;
    exp_55_ram[2658] = 160;
    exp_55_ram[2659] = 79;
    exp_55_ram[2660] = 4;
    exp_55_ram[2661] = 192;
    exp_55_ram[2662] = 0;
    exp_55_ram[2663] = 135;
    exp_55_ram[2664] = 7;
    exp_55_ram[2665] = 196;
    exp_55_ram[2666] = 207;
    exp_55_ram[2667] = 0;
    exp_55_ram[2668] = 135;
    exp_55_ram[2669] = 128;
    exp_55_ram[2670] = 247;
    exp_55_ram[2671] = 7;
    exp_55_ram[2672] = 31;
    exp_55_ram[2673] = 196;
    exp_55_ram[2674] = 23;
    exp_55_ram[2675] = 244;
    exp_55_ram[2676] = 196;
    exp_55_ram[2677] = 240;
    exp_55_ram[2678] = 231;
    exp_55_ram[2679] = 240;
    exp_55_ram[2680] = 244;
    exp_55_ram[2681] = 192;
    exp_55_ram[2682] = 0;
    exp_55_ram[2683] = 135;
    exp_55_ram[2684] = 7;
    exp_55_ram[2685] = 196;
    exp_55_ram[2686] = 207;
    exp_55_ram[2687] = 0;
    exp_55_ram[2688] = 135;
    exp_55_ram[2689] = 128;
    exp_55_ram[2690] = 247;
    exp_55_ram[2691] = 7;
    exp_55_ram[2692] = 31;
    exp_55_ram[2693] = 196;
    exp_55_ram[2694] = 247;
    exp_55_ram[2695] = 244;
    exp_55_ram[2696] = 196;
    exp_55_ram[2697] = 7;
    exp_55_ram[2698] = 132;
    exp_55_ram[2699] = 23;
    exp_55_ram[2700] = 244;
    exp_55_ram[2701] = 132;
    exp_55_ram[2702] = 144;
    exp_55_ram[2703] = 231;
    exp_55_ram[2704] = 0;
    exp_55_ram[2705] = 135;
    exp_55_ram[2706] = 7;
    exp_55_ram[2707] = 0;
    exp_55_ram[2708] = 79;
    exp_55_ram[2709] = 0;
    exp_55_ram[2710] = 193;
    exp_55_ram[2711] = 129;
    exp_55_ram[2712] = 1;
    exp_55_ram[2713] = 0;
    exp_55_ram[2714] = 1;
    exp_55_ram[2715] = 17;
    exp_55_ram[2716] = 129;
    exp_55_ram[2717] = 33;
    exp_55_ram[2718] = 49;
    exp_55_ram[2719] = 65;
    exp_55_ram[2720] = 81;
    exp_55_ram[2721] = 97;
    exp_55_ram[2722] = 113;
    exp_55_ram[2723] = 129;
    exp_55_ram[2724] = 145;
    exp_55_ram[2725] = 161;
    exp_55_ram[2726] = 177;
    exp_55_ram[2727] = 1;
    exp_55_ram[2728] = 16;
    exp_55_ram[2729] = 244;
    exp_55_ram[2730] = 16;
    exp_55_ram[2731] = 0;
    exp_55_ram[2732] = 228;
    exp_55_ram[2733] = 244;
    exp_55_ram[2734] = 79;
    exp_55_ram[2735] = 164;
    exp_55_ram[2736] = 180;
    exp_55_ram[2737] = 4;
    exp_55_ram[2738] = 0;
    exp_55_ram[2739] = 196;
    exp_55_ram[2740] = 52;
    exp_55_ram[2741] = 135;
    exp_55_ram[2742] = 247;
    exp_55_ram[2743] = 244;
    exp_55_ram[2744] = 196;
    exp_55_ram[2745] = 52;
    exp_55_ram[2746] = 135;
    exp_55_ram[2747] = 247;
    exp_55_ram[2748] = 244;
    exp_55_ram[2749] = 196;
    exp_55_ram[2750] = 52;
    exp_55_ram[2751] = 135;
    exp_55_ram[2752] = 247;
    exp_55_ram[2753] = 244;
    exp_55_ram[2754] = 196;
    exp_55_ram[2755] = 52;
    exp_55_ram[2756] = 135;
    exp_55_ram[2757] = 247;
    exp_55_ram[2758] = 244;
    exp_55_ram[2759] = 196;
    exp_55_ram[2760] = 71;
    exp_55_ram[2761] = 244;
    exp_55_ram[2762] = 79;
    exp_55_ram[2763] = 5;
    exp_55_ram[2764] = 5;
    exp_55_ram[2765] = 4;
    exp_55_ram[2766] = 68;
    exp_55_ram[2767] = 166;
    exp_55_ram[2768] = 7;
    exp_55_ram[2769] = 6;
    exp_55_ram[2770] = 182;
    exp_55_ram[2771] = 7;
    exp_55_ram[2772] = 6;
    exp_55_ram[2773] = 0;
    exp_55_ram[2774] = 134;
    exp_55_ram[2775] = 212;
    exp_55_ram[2776] = 4;
    exp_55_ram[2777] = 132;
    exp_55_ram[2778] = 196;
    exp_55_ram[2779] = 5;
    exp_55_ram[2780] = 7;
    exp_55_ram[2781] = 198;
    exp_55_ram[2782] = 5;
    exp_55_ram[2783] = 7;
    exp_55_ram[2784] = 214;
    exp_55_ram[2785] = 5;
    exp_55_ram[2786] = 7;
    exp_55_ram[2787] = 215;
    exp_55_ram[2788] = 196;
    exp_55_ram[2789] = 0;
    exp_55_ram[2790] = 7;
    exp_55_ram[2791] = 159;
    exp_55_ram[2792] = 0;
    exp_55_ram[2793] = 199;
    exp_55_ram[2794] = 15;
    exp_55_ram[2795] = 15;
    exp_55_ram[2796] = 164;
    exp_55_ram[2797] = 180;
    exp_55_ram[2798] = 4;
    exp_55_ram[2799] = 0;
    exp_55_ram[2800] = 4;
    exp_55_ram[2801] = 68;
    exp_55_ram[2802] = 52;
    exp_55_ram[2803] = 134;
    exp_55_ram[2804] = 215;
    exp_55_ram[2805] = 0;
    exp_55_ram[2806] = 215;
    exp_55_ram[2807] = 214;
    exp_55_ram[2808] = 52;
    exp_55_ram[2809] = 134;
    exp_55_ram[2810] = 215;
    exp_55_ram[2811] = 215;
    exp_55_ram[2812] = 5;
    exp_55_ram[2813] = 54;
    exp_55_ram[2814] = 7;
    exp_55_ram[2815] = 36;
    exp_55_ram[2816] = 52;
    exp_55_ram[2817] = 4;
    exp_55_ram[2818] = 68;
    exp_55_ram[2819] = 52;
    exp_55_ram[2820] = 134;
    exp_55_ram[2821] = 215;
    exp_55_ram[2822] = 0;
    exp_55_ram[2823] = 215;
    exp_55_ram[2824] = 214;
    exp_55_ram[2825] = 52;
    exp_55_ram[2826] = 134;
    exp_55_ram[2827] = 215;
    exp_55_ram[2828] = 215;
    exp_55_ram[2829] = 5;
    exp_55_ram[2830] = 86;
    exp_55_ram[2831] = 7;
    exp_55_ram[2832] = 68;
    exp_55_ram[2833] = 84;
    exp_55_ram[2834] = 4;
    exp_55_ram[2835] = 68;
    exp_55_ram[2836] = 52;
    exp_55_ram[2837] = 134;
    exp_55_ram[2838] = 215;
    exp_55_ram[2839] = 0;
    exp_55_ram[2840] = 215;
    exp_55_ram[2841] = 214;
    exp_55_ram[2842] = 52;
    exp_55_ram[2843] = 134;
    exp_55_ram[2844] = 215;
    exp_55_ram[2845] = 215;
    exp_55_ram[2846] = 5;
    exp_55_ram[2847] = 118;
    exp_55_ram[2848] = 7;
    exp_55_ram[2849] = 100;
    exp_55_ram[2850] = 116;
    exp_55_ram[2851] = 4;
    exp_55_ram[2852] = 68;
    exp_55_ram[2853] = 52;
    exp_55_ram[2854] = 134;
    exp_55_ram[2855] = 215;
    exp_55_ram[2856] = 0;
    exp_55_ram[2857] = 215;
    exp_55_ram[2858] = 214;
    exp_55_ram[2859] = 52;
    exp_55_ram[2860] = 134;
    exp_55_ram[2861] = 215;
    exp_55_ram[2862] = 215;
    exp_55_ram[2863] = 5;
    exp_55_ram[2864] = 150;
    exp_55_ram[2865] = 7;
    exp_55_ram[2866] = 132;
    exp_55_ram[2867] = 148;
    exp_55_ram[2868] = 196;
    exp_55_ram[2869] = 71;
    exp_55_ram[2870] = 244;
    exp_55_ram[2871] = 15;
    exp_55_ram[2872] = 5;
    exp_55_ram[2873] = 5;
    exp_55_ram[2874] = 4;
    exp_55_ram[2875] = 68;
    exp_55_ram[2876] = 166;
    exp_55_ram[2877] = 7;
    exp_55_ram[2878] = 6;
    exp_55_ram[2879] = 182;
    exp_55_ram[2880] = 7;
    exp_55_ram[2881] = 6;
    exp_55_ram[2882] = 0;
    exp_55_ram[2883] = 134;
    exp_55_ram[2884] = 212;
    exp_55_ram[2885] = 4;
    exp_55_ram[2886] = 4;
    exp_55_ram[2887] = 68;
    exp_55_ram[2888] = 5;
    exp_55_ram[2889] = 7;
    exp_55_ram[2890] = 198;
    exp_55_ram[2891] = 5;
    exp_55_ram[2892] = 7;
    exp_55_ram[2893] = 214;
    exp_55_ram[2894] = 5;
    exp_55_ram[2895] = 7;
    exp_55_ram[2896] = 215;
    exp_55_ram[2897] = 196;
    exp_55_ram[2898] = 0;
    exp_55_ram[2899] = 7;
    exp_55_ram[2900] = 95;
    exp_55_ram[2901] = 0;
    exp_55_ram[2902] = 71;
    exp_55_ram[2903] = 207;
    exp_55_ram[2904] = 207;
    exp_55_ram[2905] = 164;
    exp_55_ram[2906] = 180;
    exp_55_ram[2907] = 4;
    exp_55_ram[2908] = 0;
    exp_55_ram[2909] = 196;
    exp_55_ram[2910] = 52;
    exp_55_ram[2911] = 135;
    exp_55_ram[2912] = 247;
    exp_55_ram[2913] = 244;
    exp_55_ram[2914] = 196;
    exp_55_ram[2915] = 52;
    exp_55_ram[2916] = 135;
    exp_55_ram[2917] = 247;
    exp_55_ram[2918] = 244;
    exp_55_ram[2919] = 196;
    exp_55_ram[2920] = 52;
    exp_55_ram[2921] = 135;
    exp_55_ram[2922] = 247;
    exp_55_ram[2923] = 244;
    exp_55_ram[2924] = 196;
    exp_55_ram[2925] = 52;
    exp_55_ram[2926] = 135;
    exp_55_ram[2927] = 247;
    exp_55_ram[2928] = 244;
    exp_55_ram[2929] = 196;
    exp_55_ram[2930] = 71;
    exp_55_ram[2931] = 244;
    exp_55_ram[2932] = 207;
    exp_55_ram[2933] = 5;
    exp_55_ram[2934] = 5;
    exp_55_ram[2935] = 4;
    exp_55_ram[2936] = 68;
    exp_55_ram[2937] = 166;
    exp_55_ram[2938] = 7;
    exp_55_ram[2939] = 6;
    exp_55_ram[2940] = 182;
    exp_55_ram[2941] = 7;
    exp_55_ram[2942] = 6;
    exp_55_ram[2943] = 0;
    exp_55_ram[2944] = 134;
    exp_55_ram[2945] = 212;
    exp_55_ram[2946] = 4;
    exp_55_ram[2947] = 132;
    exp_55_ram[2948] = 196;
    exp_55_ram[2949] = 5;
    exp_55_ram[2950] = 7;
    exp_55_ram[2951] = 198;
    exp_55_ram[2952] = 5;
    exp_55_ram[2953] = 7;
    exp_55_ram[2954] = 214;
    exp_55_ram[2955] = 5;
    exp_55_ram[2956] = 7;
    exp_55_ram[2957] = 215;
    exp_55_ram[2958] = 196;
    exp_55_ram[2959] = 0;
    exp_55_ram[2960] = 7;
    exp_55_ram[2961] = 31;
    exp_55_ram[2962] = 0;
    exp_55_ram[2963] = 199;
    exp_55_ram[2964] = 159;
    exp_55_ram[2965] = 143;
    exp_55_ram[2966] = 164;
    exp_55_ram[2967] = 180;
    exp_55_ram[2968] = 4;
    exp_55_ram[2969] = 0;
    exp_55_ram[2970] = 4;
    exp_55_ram[2971] = 68;
    exp_55_ram[2972] = 52;
    exp_55_ram[2973] = 134;
    exp_55_ram[2974] = 0;
    exp_55_ram[2975] = 7;
    exp_55_ram[2976] = 7;
    exp_55_ram[2977] = 143;
    exp_55_ram[2978] = 5;
    exp_55_ram[2979] = 5;
    exp_55_ram[2980] = 228;
    exp_55_ram[2981] = 244;
    exp_55_ram[2982] = 4;
    exp_55_ram[2983] = 68;
    exp_55_ram[2984] = 52;
    exp_55_ram[2985] = 134;
    exp_55_ram[2986] = 0;
    exp_55_ram[2987] = 7;
    exp_55_ram[2988] = 7;
    exp_55_ram[2989] = 143;
    exp_55_ram[2990] = 5;
    exp_55_ram[2991] = 5;
    exp_55_ram[2992] = 228;
    exp_55_ram[2993] = 244;
    exp_55_ram[2994] = 4;
    exp_55_ram[2995] = 68;
    exp_55_ram[2996] = 52;
    exp_55_ram[2997] = 134;
    exp_55_ram[2998] = 0;
    exp_55_ram[2999] = 7;
    exp_55_ram[3000] = 7;
    exp_55_ram[3001] = 143;
    exp_55_ram[3002] = 5;
    exp_55_ram[3003] = 5;
    exp_55_ram[3004] = 228;
    exp_55_ram[3005] = 244;
    exp_55_ram[3006] = 4;
    exp_55_ram[3007] = 68;
    exp_55_ram[3008] = 52;
    exp_55_ram[3009] = 134;
    exp_55_ram[3010] = 0;
    exp_55_ram[3011] = 7;
    exp_55_ram[3012] = 7;
    exp_55_ram[3013] = 143;
    exp_55_ram[3014] = 5;
    exp_55_ram[3015] = 5;
    exp_55_ram[3016] = 228;
    exp_55_ram[3017] = 244;
    exp_55_ram[3018] = 196;
    exp_55_ram[3019] = 71;
    exp_55_ram[3020] = 244;
    exp_55_ram[3021] = 143;
    exp_55_ram[3022] = 5;
    exp_55_ram[3023] = 5;
    exp_55_ram[3024] = 4;
    exp_55_ram[3025] = 68;
    exp_55_ram[3026] = 166;
    exp_55_ram[3027] = 7;
    exp_55_ram[3028] = 6;
    exp_55_ram[3029] = 182;
    exp_55_ram[3030] = 7;
    exp_55_ram[3031] = 6;
    exp_55_ram[3032] = 0;
    exp_55_ram[3033] = 134;
    exp_55_ram[3034] = 6;
    exp_55_ram[3035] = 0;
    exp_55_ram[3036] = 13;
    exp_55_ram[3037] = 7;
    exp_55_ram[3038] = 198;
    exp_55_ram[3039] = 13;
    exp_55_ram[3040] = 7;
    exp_55_ram[3041] = 214;
    exp_55_ram[3042] = 13;
    exp_55_ram[3043] = 7;
    exp_55_ram[3044] = 215;
    exp_55_ram[3045] = 196;
    exp_55_ram[3046] = 0;
    exp_55_ram[3047] = 7;
    exp_55_ram[3048] = 79;
    exp_55_ram[3049] = 0;
    exp_55_ram[3050] = 7;
    exp_55_ram[3051] = 223;
    exp_55_ram[3052] = 0;
    exp_55_ram[3053] = 193;
    exp_55_ram[3054] = 129;
    exp_55_ram[3055] = 65;
    exp_55_ram[3056] = 1;
    exp_55_ram[3057] = 193;
    exp_55_ram[3058] = 129;
    exp_55_ram[3059] = 65;
    exp_55_ram[3060] = 1;
    exp_55_ram[3061] = 193;
    exp_55_ram[3062] = 129;
    exp_55_ram[3063] = 65;
    exp_55_ram[3064] = 1;
    exp_55_ram[3065] = 1;
    exp_55_ram[3066] = 0;
    exp_55_ram[3067] = 1;
    exp_55_ram[3068] = 17;
    exp_55_ram[3069] = 129;
    exp_55_ram[3070] = 33;
    exp_55_ram[3071] = 49;
    exp_55_ram[3072] = 65;
    exp_55_ram[3073] = 81;
    exp_55_ram[3074] = 1;
    exp_55_ram[3075] = 0;
    exp_55_ram[3076] = 71;
    exp_55_ram[3077] = 95;
    exp_55_ram[3078] = 79;
    exp_55_ram[3079] = 5;
    exp_55_ram[3080] = 71;
    exp_55_ram[3081] = 244;
    exp_55_ram[3082] = 0;
    exp_55_ram[3083] = 199;
    exp_55_ram[3084] = 159;
    exp_55_ram[3085] = 143;
    exp_55_ram[3086] = 5;
    exp_55_ram[3087] = 247;
    exp_55_ram[3088] = 244;
    exp_55_ram[3089] = 0;
    exp_55_ram[3090] = 71;
    exp_55_ram[3091] = 223;
    exp_55_ram[3092] = 207;
    exp_55_ram[3093] = 5;
    exp_55_ram[3094] = 244;
    exp_55_ram[3095] = 0;
    exp_55_ram[3096] = 199;
    exp_55_ram[3097] = 95;
    exp_55_ram[3098] = 79;
    exp_55_ram[3099] = 5;
    exp_55_ram[3100] = 244;
    exp_55_ram[3101] = 0;
    exp_55_ram[3102] = 71;
    exp_55_ram[3103] = 223;
    exp_55_ram[3104] = 207;
    exp_55_ram[3105] = 5;
    exp_55_ram[3106] = 244;
    exp_55_ram[3107] = 112;
    exp_55_ram[3108] = 244;
    exp_55_ram[3109] = 16;
    exp_55_ram[3110] = 244;
    exp_55_ram[3111] = 4;
    exp_55_ram[3112] = 7;
    exp_55_ram[3113] = 15;
    exp_55_ram[3114] = 5;
    exp_55_ram[3115] = 5;
    exp_55_ram[3116] = 228;
    exp_55_ram[3117] = 244;
    exp_55_ram[3118] = 132;
    exp_55_ram[3119] = 196;
    exp_55_ram[3120] = 7;
    exp_55_ram[3121] = 7;
    exp_55_ram[3122] = 95;
    exp_55_ram[3123] = 15;
    exp_55_ram[3124] = 164;
    exp_55_ram[3125] = 180;
    exp_55_ram[3126] = 4;
    exp_55_ram[3127] = 128;
    exp_55_ram[3128] = 0;
    exp_55_ram[3129] = 143;
    exp_55_ram[3130] = 5;
    exp_55_ram[3131] = 5;
    exp_55_ram[3132] = 132;
    exp_55_ram[3133] = 196;
    exp_55_ram[3134] = 7;
    exp_55_ram[3135] = 7;
    exp_55_ram[3136] = 15;
    exp_55_ram[3137] = 5;
    exp_55_ram[3138] = 5;
    exp_55_ram[3139] = 0;
    exp_55_ram[3140] = 135;
    exp_55_ram[3141] = 7;
    exp_55_ram[3142] = 207;
    exp_55_ram[3143] = 5;
    exp_55_ram[3144] = 5;
    exp_55_ram[3145] = 7;
    exp_55_ram[3146] = 7;
    exp_55_ram[3147] = 10;
    exp_55_ram[3148] = 10;
    exp_55_ram[3149] = 207;
    exp_55_ram[3150] = 5;
    exp_55_ram[3151] = 7;
    exp_55_ram[3152] = 0;
    exp_55_ram[3153] = 135;
    exp_55_ram[3154] = 7;
    exp_55_ram[3155] = 0;
    exp_55_ram[3156] = 132;
    exp_55_ram[3157] = 196;
    exp_55_ram[3158] = 38;
    exp_55_ram[3159] = 7;
    exp_55_ram[3160] = 197;
    exp_55_ram[3161] = 54;
    exp_55_ram[3162] = 245;
    exp_55_ram[3163] = 6;
    exp_55_ram[3164] = 228;
    exp_55_ram[3165] = 244;
    exp_55_ram[3166] = 0;
    exp_55_ram[3167] = 223;
    exp_55_ram[3168] = 5;
    exp_55_ram[3169] = 5;
    exp_55_ram[3170] = 228;
    exp_55_ram[3171] = 244;
    exp_55_ram[3172] = 132;
    exp_55_ram[3173] = 7;
    exp_55_ram[3174] = 223;
    exp_55_ram[3175] = 5;
    exp_55_ram[3176] = 7;
    exp_55_ram[3177] = 95;
    exp_55_ram[3178] = 68;
    exp_55_ram[3179] = 23;
    exp_55_ram[3180] = 244;
    exp_55_ram[3181] = 68;
    exp_55_ram[3182] = 48;
    exp_55_ram[3183] = 231;
    exp_55_ram[3184] = 0;
    exp_55_ram[3185] = 0;
    exp_55_ram[3186] = 193;
    exp_55_ram[3187] = 129;
    exp_55_ram[3188] = 65;
    exp_55_ram[3189] = 1;
    exp_55_ram[3190] = 193;
    exp_55_ram[3191] = 129;
    exp_55_ram[3192] = 1;
    exp_55_ram[3193] = 0;
    exp_55_ram[3194] = 1;
    exp_55_ram[3195] = 17;
    exp_55_ram[3196] = 129;
    exp_55_ram[3197] = 1;
    exp_55_ram[3198] = 0;
    exp_55_ram[3199] = 199;
    exp_55_ram[3200] = 159;
    exp_55_ram[3201] = 0;
    exp_55_ram[3202] = 199;
    exp_55_ram[3203] = 223;
    exp_55_ram[3204] = 0;
    exp_55_ram[3205] = 199;
    exp_55_ram[3206] = 31;
    exp_55_ram[3207] = 0;
    exp_55_ram[3208] = 199;
    exp_55_ram[3209] = 95;
    exp_55_ram[3210] = 0;
    exp_55_ram[3211] = 71;
    exp_55_ram[3212] = 159;
    exp_55_ram[3213] = 0;
    exp_55_ram[3214] = 71;
    exp_55_ram[3215] = 223;
    exp_55_ram[3216] = 0;
    exp_55_ram[3217] = 135;
    exp_55_ram[3218] = 31;
    exp_55_ram[3219] = 95;
    exp_55_ram[3220] = 5;
    exp_55_ram[3221] = 244;
    exp_55_ram[3222] = 244;
    exp_55_ram[3223] = 247;
    exp_55_ram[3224] = 80;
    exp_55_ram[3225] = 247;
    exp_55_ram[3226] = 39;
    exp_55_ram[3227] = 0;
    exp_55_ram[3228] = 199;
    exp_55_ram[3229] = 247;
    exp_55_ram[3230] = 7;
    exp_55_ram[3231] = 7;
    exp_55_ram[3232] = 143;
    exp_55_ram[3233] = 192;
    exp_55_ram[3234] = 15;
    exp_55_ram[3235] = 64;
    exp_55_ram[3236] = 143;
    exp_55_ram[3237] = 192;
    exp_55_ram[3238] = 95;
    exp_55_ram[3239] = 64;
    exp_55_ram[3240] = 144;
    exp_55_ram[3241] = 192;
    exp_55_ram[3242] = 15;
    exp_55_ram[3243] = 0;
    exp_55_ram[3244] = 159;
    exp_55_ram[3245] = 1;
    exp_55_ram[3246] = 129;
    exp_55_ram[3247] = 1;
    exp_55_ram[3248] = 5;
    exp_55_ram[3249] = 244;
    exp_55_ram[3250] = 244;
    exp_55_ram[3251] = 167;
    exp_55_ram[3252] = 160;
    exp_55_ram[3253] = 247;
    exp_55_ram[3254] = 247;
    exp_55_ram[3255] = 7;
    exp_55_ram[3256] = 193;
    exp_55_ram[3257] = 1;
    exp_55_ram[3258] = 0;
    exp_55_ram[3259] = 1;
    exp_55_ram[3260] = 17;
    exp_55_ram[3261] = 129;
    exp_55_ram[3262] = 145;
    exp_55_ram[3263] = 1;
    exp_55_ram[3264] = 164;
    exp_55_ram[3265] = 180;
    exp_55_ram[3266] = 196;
    exp_55_ram[3267] = 212;
    exp_55_ram[3268] = 228;
    exp_55_ram[3269] = 8;
    exp_55_ram[3270] = 8;
    exp_55_ram[3271] = 244;
    exp_55_ram[3272] = 6;
    exp_55_ram[3273] = 244;
    exp_55_ram[3274] = 7;
    exp_55_ram[3275] = 244;
    exp_55_ram[3276] = 4;
    exp_55_ram[3277] = 247;
    exp_55_ram[3278] = 247;
    exp_55_ram[3279] = 196;
    exp_55_ram[3280] = 231;
    exp_55_ram[3281] = 68;
    exp_55_ram[3282] = 247;
    exp_55_ram[3283] = 247;
    exp_55_ram[3284] = 196;
    exp_55_ram[3285] = 231;
    exp_55_ram[3286] = 132;
    exp_55_ram[3287] = 247;
    exp_55_ram[3288] = 247;
    exp_55_ram[3289] = 196;
    exp_55_ram[3290] = 231;
    exp_55_ram[3291] = 68;
    exp_55_ram[3292] = 167;
    exp_55_ram[3293] = 7;
    exp_55_ram[3294] = 247;
    exp_55_ram[3295] = 247;
    exp_55_ram[3296] = 196;
    exp_55_ram[3297] = 231;
    exp_55_ram[3298] = 4;
    exp_55_ram[3299] = 167;
    exp_55_ram[3300] = 7;
    exp_55_ram[3301] = 247;
    exp_55_ram[3302] = 247;
    exp_55_ram[3303] = 196;
    exp_55_ram[3304] = 231;
    exp_55_ram[3305] = 180;
    exp_55_ram[3306] = 247;
    exp_55_ram[3307] = 247;
    exp_55_ram[3308] = 196;
    exp_55_ram[3309] = 231;
    exp_55_ram[3310] = 164;
    exp_55_ram[3311] = 247;
    exp_55_ram[3312] = 247;
    exp_55_ram[3313] = 196;
    exp_55_ram[3314] = 231;
    exp_55_ram[3315] = 148;
    exp_55_ram[3316] = 247;
    exp_55_ram[3317] = 247;
    exp_55_ram[3318] = 196;
    exp_55_ram[3319] = 231;
    exp_55_ram[3320] = 4;
    exp_55_ram[3321] = 192;
    exp_55_ram[3322] = 244;
    exp_55_ram[3323] = 132;
    exp_55_ram[3324] = 247;
    exp_55_ram[3325] = 7;
    exp_55_ram[3326] = 247;
    exp_55_ram[3327] = 244;
    exp_55_ram[3328] = 244;
    exp_55_ram[3329] = 68;
    exp_55_ram[3330] = 247;
    exp_55_ram[3331] = 7;
    exp_55_ram[3332] = 247;
    exp_55_ram[3333] = 244;
    exp_55_ram[3334] = 244;
    exp_55_ram[3335] = 4;
    exp_55_ram[3336] = 247;
    exp_55_ram[3337] = 7;
    exp_55_ram[3338] = 247;
    exp_55_ram[3339] = 244;
    exp_55_ram[3340] = 244;
    exp_55_ram[3341] = 196;
    exp_55_ram[3342] = 247;
    exp_55_ram[3343] = 7;
    exp_55_ram[3344] = 247;
    exp_55_ram[3345] = 244;
    exp_55_ram[3346] = 244;
    exp_55_ram[3347] = 7;
    exp_55_ram[3348] = 95;
    exp_55_ram[3349] = 5;
    exp_55_ram[3350] = 7;
    exp_55_ram[3351] = 196;
    exp_55_ram[3352] = 231;
    exp_55_ram[3353] = 228;
    exp_55_ram[3354] = 231;
    exp_55_ram[3355] = 244;
    exp_55_ram[3356] = 7;
    exp_55_ram[3357] = 31;
    exp_55_ram[3358] = 5;
    exp_55_ram[3359] = 7;
    exp_55_ram[3360] = 196;
    exp_55_ram[3361] = 231;
    exp_55_ram[3362] = 212;
    exp_55_ram[3363] = 231;
    exp_55_ram[3364] = 244;
    exp_55_ram[3365] = 7;
    exp_55_ram[3366] = 223;
    exp_55_ram[3367] = 5;
    exp_55_ram[3368] = 7;
    exp_55_ram[3369] = 196;
    exp_55_ram[3370] = 231;
    exp_55_ram[3371] = 196;
    exp_55_ram[3372] = 231;
    exp_55_ram[3373] = 244;
    exp_55_ram[3374] = 196;
    exp_55_ram[3375] = 247;
    exp_55_ram[3376] = 180;
    exp_55_ram[3377] = 231;
    exp_55_ram[3378] = 228;
    exp_55_ram[3379] = 244;
    exp_55_ram[3380] = 7;
    exp_55_ram[3381] = 31;
    exp_55_ram[3382] = 5;
    exp_55_ram[3383] = 7;
    exp_55_ram[3384] = 196;
    exp_55_ram[3385] = 151;
    exp_55_ram[3386] = 231;
    exp_55_ram[3387] = 212;
    exp_55_ram[3388] = 244;
    exp_55_ram[3389] = 7;
    exp_55_ram[3390] = 223;
    exp_55_ram[3391] = 5;
    exp_55_ram[3392] = 7;
    exp_55_ram[3393] = 196;
    exp_55_ram[3394] = 151;
    exp_55_ram[3395] = 231;
    exp_55_ram[3396] = 196;
    exp_55_ram[3397] = 244;
    exp_55_ram[3398] = 7;
    exp_55_ram[3399] = 159;
    exp_55_ram[3400] = 5;
    exp_55_ram[3401] = 7;
    exp_55_ram[3402] = 196;
    exp_55_ram[3403] = 151;
    exp_55_ram[3404] = 231;
    exp_55_ram[3405] = 244;
    exp_55_ram[3406] = 23;
    exp_55_ram[3407] = 244;
    exp_55_ram[3408] = 244;
    exp_55_ram[3409] = 144;
    exp_55_ram[3410] = 231;
    exp_55_ram[3411] = 0;
    exp_55_ram[3412] = 0;
    exp_55_ram[3413] = 193;
    exp_55_ram[3414] = 129;
    exp_55_ram[3415] = 65;
    exp_55_ram[3416] = 1;
    exp_55_ram[3417] = 0;
    exp_55_ram[3418] = 1;
    exp_55_ram[3419] = 17;
    exp_55_ram[3420] = 129;
    exp_55_ram[3421] = 1;
    exp_55_ram[3422] = 164;
    exp_55_ram[3423] = 5;
    exp_55_ram[3424] = 244;
    exp_55_ram[3425] = 196;
    exp_55_ram[3426] = 199;
    exp_55_ram[3427] = 196;
    exp_55_ram[3428] = 151;
    exp_55_ram[3429] = 247;
    exp_55_ram[3430] = 196;
    exp_55_ram[3431] = 183;
    exp_55_ram[3432] = 23;
    exp_55_ram[3433] = 247;
    exp_55_ram[3434] = 7;
    exp_55_ram[3435] = 159;
    exp_55_ram[3436] = 5;
    exp_55_ram[3437] = 7;
    exp_55_ram[3438] = 196;
    exp_55_ram[3439] = 231;
    exp_55_ram[3440] = 196;
    exp_55_ram[3441] = 215;
    exp_55_ram[3442] = 196;
    exp_55_ram[3443] = 167;
    exp_55_ram[3444] = 247;
    exp_55_ram[3445] = 196;
    exp_55_ram[3446] = 199;
    exp_55_ram[3447] = 23;
    exp_55_ram[3448] = 247;
    exp_55_ram[3449] = 7;
    exp_55_ram[3450] = 223;
    exp_55_ram[3451] = 5;
    exp_55_ram[3452] = 7;
    exp_55_ram[3453] = 196;
    exp_55_ram[3454] = 231;
    exp_55_ram[3455] = 196;
    exp_55_ram[3456] = 215;
    exp_55_ram[3457] = 23;
    exp_55_ram[3458] = 247;
    exp_55_ram[3459] = 7;
    exp_55_ram[3460] = 95;
    exp_55_ram[3461] = 5;
    exp_55_ram[3462] = 7;
    exp_55_ram[3463] = 196;
    exp_55_ram[3464] = 231;
    exp_55_ram[3465] = 180;
    exp_55_ram[3466] = 247;
    exp_55_ram[3467] = 244;
    exp_55_ram[3468] = 196;
    exp_55_ram[3469] = 215;
    exp_55_ram[3470] = 244;
    exp_55_ram[3471] = 247;
    exp_55_ram[3472] = 247;
    exp_55_ram[3473] = 196;
    exp_55_ram[3474] = 135;
    exp_55_ram[3475] = 247;
    exp_55_ram[3476] = 247;
    exp_55_ram[3477] = 7;
    exp_55_ram[3478] = 223;
    exp_55_ram[3479] = 5;
    exp_55_ram[3480] = 7;
    exp_55_ram[3481] = 196;
    exp_55_ram[3482] = 231;
    exp_55_ram[3483] = 71;
    exp_55_ram[3484] = 196;
    exp_55_ram[3485] = 215;
    exp_55_ram[3486] = 247;
    exp_55_ram[3487] = 247;
    exp_55_ram[3488] = 196;
    exp_55_ram[3489] = 135;
    exp_55_ram[3490] = 247;
    exp_55_ram[3491] = 247;
    exp_55_ram[3492] = 7;
    exp_55_ram[3493] = 31;
    exp_55_ram[3494] = 5;
    exp_55_ram[3495] = 244;
    exp_55_ram[3496] = 196;
    exp_55_ram[3497] = 199;
    exp_55_ram[3498] = 244;
    exp_55_ram[3499] = 247;
    exp_55_ram[3500] = 247;
    exp_55_ram[3501] = 196;
    exp_55_ram[3502] = 119;
    exp_55_ram[3503] = 247;
    exp_55_ram[3504] = 247;
    exp_55_ram[3505] = 7;
    exp_55_ram[3506] = 223;
    exp_55_ram[3507] = 5;
    exp_55_ram[3508] = 7;
    exp_55_ram[3509] = 196;
    exp_55_ram[3510] = 231;
    exp_55_ram[3511] = 231;
    exp_55_ram[3512] = 196;
    exp_55_ram[3513] = 199;
    exp_55_ram[3514] = 247;
    exp_55_ram[3515] = 247;
    exp_55_ram[3516] = 196;
    exp_55_ram[3517] = 119;
    exp_55_ram[3518] = 247;
    exp_55_ram[3519] = 247;
    exp_55_ram[3520] = 7;
    exp_55_ram[3521] = 31;
    exp_55_ram[3522] = 5;
    exp_55_ram[3523] = 244;
    exp_55_ram[3524] = 196;
    exp_55_ram[3525] = 183;
    exp_55_ram[3526] = 244;
    exp_55_ram[3527] = 247;
    exp_55_ram[3528] = 247;
    exp_55_ram[3529] = 196;
    exp_55_ram[3530] = 103;
    exp_55_ram[3531] = 247;
    exp_55_ram[3532] = 247;
    exp_55_ram[3533] = 7;
    exp_55_ram[3534] = 223;
    exp_55_ram[3535] = 5;
    exp_55_ram[3536] = 7;
    exp_55_ram[3537] = 196;
    exp_55_ram[3538] = 231;
    exp_55_ram[3539] = 167;
    exp_55_ram[3540] = 196;
    exp_55_ram[3541] = 183;
    exp_55_ram[3542] = 247;
    exp_55_ram[3543] = 247;
    exp_55_ram[3544] = 196;
    exp_55_ram[3545] = 103;
    exp_55_ram[3546] = 247;
    exp_55_ram[3547] = 247;
    exp_55_ram[3548] = 7;
    exp_55_ram[3549] = 31;
    exp_55_ram[3550] = 5;
    exp_55_ram[3551] = 244;
    exp_55_ram[3552] = 244;
    exp_55_ram[3553] = 196;
    exp_55_ram[3554] = 247;
    exp_55_ram[3555] = 7;
    exp_55_ram[3556] = 244;
    exp_55_ram[3557] = 196;
    exp_55_ram[3558] = 183;
    exp_55_ram[3559] = 244;
    exp_55_ram[3560] = 247;
    exp_55_ram[3561] = 247;
    exp_55_ram[3562] = 196;
    exp_55_ram[3563] = 103;
    exp_55_ram[3564] = 247;
    exp_55_ram[3565] = 247;
    exp_55_ram[3566] = 7;
    exp_55_ram[3567] = 159;
    exp_55_ram[3568] = 5;
    exp_55_ram[3569] = 7;
    exp_55_ram[3570] = 196;
    exp_55_ram[3571] = 231;
    exp_55_ram[3572] = 135;
    exp_55_ram[3573] = 196;
    exp_55_ram[3574] = 183;
    exp_55_ram[3575] = 247;
    exp_55_ram[3576] = 247;
    exp_55_ram[3577] = 196;
    exp_55_ram[3578] = 103;
    exp_55_ram[3579] = 247;
    exp_55_ram[3580] = 247;
    exp_55_ram[3581] = 7;
    exp_55_ram[3582] = 223;
    exp_55_ram[3583] = 5;
    exp_55_ram[3584] = 244;
    exp_55_ram[3585] = 196;
    exp_55_ram[3586] = 199;
    exp_55_ram[3587] = 244;
    exp_55_ram[3588] = 247;
    exp_55_ram[3589] = 247;
    exp_55_ram[3590] = 196;
    exp_55_ram[3591] = 119;
    exp_55_ram[3592] = 247;
    exp_55_ram[3593] = 247;
    exp_55_ram[3594] = 7;
    exp_55_ram[3595] = 159;
    exp_55_ram[3596] = 5;
    exp_55_ram[3597] = 7;
    exp_55_ram[3598] = 196;
    exp_55_ram[3599] = 231;
    exp_55_ram[3600] = 199;
    exp_55_ram[3601] = 196;
    exp_55_ram[3602] = 199;
    exp_55_ram[3603] = 247;
    exp_55_ram[3604] = 247;
    exp_55_ram[3605] = 196;
    exp_55_ram[3606] = 119;
    exp_55_ram[3607] = 247;
    exp_55_ram[3608] = 247;
    exp_55_ram[3609] = 7;
    exp_55_ram[3610] = 223;
    exp_55_ram[3611] = 5;
    exp_55_ram[3612] = 244;
    exp_55_ram[3613] = 196;
    exp_55_ram[3614] = 215;
    exp_55_ram[3615] = 244;
    exp_55_ram[3616] = 247;
    exp_55_ram[3617] = 247;
    exp_55_ram[3618] = 196;
    exp_55_ram[3619] = 135;
    exp_55_ram[3620] = 247;
    exp_55_ram[3621] = 247;
    exp_55_ram[3622] = 7;
    exp_55_ram[3623] = 159;
    exp_55_ram[3624] = 5;
    exp_55_ram[3625] = 7;
    exp_55_ram[3626] = 196;
    exp_55_ram[3627] = 231;
    exp_55_ram[3628] = 39;
    exp_55_ram[3629] = 196;
    exp_55_ram[3630] = 215;
    exp_55_ram[3631] = 247;
    exp_55_ram[3632] = 247;
    exp_55_ram[3633] = 196;
    exp_55_ram[3634] = 135;
    exp_55_ram[3635] = 247;
    exp_55_ram[3636] = 247;
    exp_55_ram[3637] = 7;
    exp_55_ram[3638] = 223;
    exp_55_ram[3639] = 5;
    exp_55_ram[3640] = 244;
    exp_55_ram[3641] = 244;
    exp_55_ram[3642] = 23;
    exp_55_ram[3643] = 247;
    exp_55_ram[3644] = 7;
    exp_55_ram[3645] = 193;
    exp_55_ram[3646] = 129;
    exp_55_ram[3647] = 1;
    exp_55_ram[3648] = 0;
    exp_55_ram[3649] = 1;
    exp_55_ram[3650] = 17;
    exp_55_ram[3651] = 129;
    exp_55_ram[3652] = 1;
    exp_55_ram[3653] = 207;
    exp_55_ram[3654] = 5;
    exp_55_ram[3655] = 244;
    exp_55_ram[3656] = 244;
    exp_55_ram[3657] = 16;
    exp_55_ram[3658] = 247;
    exp_55_ram[3659] = 0;
    exp_55_ram[3660] = 71;
    exp_55_ram[3661] = 0;
    exp_55_ram[3662] = 244;
    exp_55_ram[3663] = 32;
    exp_55_ram[3664] = 247;
    exp_55_ram[3665] = 0;
    exp_55_ram[3666] = 7;
    exp_55_ram[3667] = 128;
    exp_55_ram[3668] = 244;
    exp_55_ram[3669] = 48;
    exp_55_ram[3670] = 247;
    exp_55_ram[3671] = 0;
    exp_55_ram[3672] = 199;
    exp_55_ram[3673] = 0;
    exp_55_ram[3674] = 244;
    exp_55_ram[3675] = 64;
    exp_55_ram[3676] = 247;
    exp_55_ram[3677] = 0;
    exp_55_ram[3678] = 135;
    exp_55_ram[3679] = 128;
    exp_55_ram[3680] = 244;
    exp_55_ram[3681] = 80;
    exp_55_ram[3682] = 247;
    exp_55_ram[3683] = 0;
    exp_55_ram[3684] = 71;
    exp_55_ram[3685] = 7;
    exp_55_ram[3686] = 193;
    exp_55_ram[3687] = 129;
    exp_55_ram[3688] = 1;
    exp_55_ram[3689] = 0;
    exp_55_ram[3690] = 1;
    exp_55_ram[3691] = 17;
    exp_55_ram[3692] = 129;
    exp_55_ram[3693] = 1;
    exp_55_ram[3694] = 143;
    exp_55_ram[3695] = 5;
    exp_55_ram[3696] = 244;
    exp_55_ram[3697] = 244;
    exp_55_ram[3698] = 7;
    exp_55_ram[3699] = 15;
    exp_55_ram[3700] = 5;
    exp_55_ram[3701] = 16;
    exp_55_ram[3702] = 247;
    exp_55_ram[3703] = 0;
    exp_55_ram[3704] = 7;
    exp_55_ram[3705] = 128;
    exp_55_ram[3706] = 244;
    exp_55_ram[3707] = 7;
    exp_55_ram[3708] = 207;
    exp_55_ram[3709] = 5;
    exp_55_ram[3710] = 32;
    exp_55_ram[3711] = 247;
    exp_55_ram[3712] = 0;
    exp_55_ram[3713] = 199;
    exp_55_ram[3714] = 64;
    exp_55_ram[3715] = 244;
    exp_55_ram[3716] = 7;
    exp_55_ram[3717] = 143;
    exp_55_ram[3718] = 5;
    exp_55_ram[3719] = 48;
    exp_55_ram[3720] = 247;
    exp_55_ram[3721] = 0;
    exp_55_ram[3722] = 135;
    exp_55_ram[3723] = 7;
    exp_55_ram[3724] = 193;
    exp_55_ram[3725] = 129;
    exp_55_ram[3726] = 1;
    exp_55_ram[3727] = 0;
    exp_55_ram[3728] = 1;
    exp_55_ram[3729] = 17;
    exp_55_ram[3730] = 129;
    exp_55_ram[3731] = 1;
    exp_55_ram[3732] = 15;
    exp_55_ram[3733] = 5;
    exp_55_ram[3734] = 244;
    exp_55_ram[3735] = 244;
    exp_55_ram[3736] = 7;
    exp_55_ram[3737] = 143;
    exp_55_ram[3738] = 5;
    exp_55_ram[3739] = 7;
    exp_55_ram[3740] = 244;
    exp_55_ram[3741] = 7;
    exp_55_ram[3742] = 79;
    exp_55_ram[3743] = 5;
    exp_55_ram[3744] = 247;
    exp_55_ram[3745] = 7;
    exp_55_ram[3746] = 193;
    exp_55_ram[3747] = 129;
    exp_55_ram[3748] = 1;
    exp_55_ram[3749] = 0;
    exp_55_ram[3750] = 1;
    exp_55_ram[3751] = 17;
    exp_55_ram[3752] = 129;
    exp_55_ram[3753] = 1;
    exp_55_ram[3754] = 0;
    exp_55_ram[3755] = 7;
    exp_55_ram[3756] = 0;
    exp_55_ram[3757] = 71;
    exp_55_ram[3758] = 0;
    exp_55_ram[3759] = 135;
    exp_55_ram[3760] = 0;
    exp_55_ram[3761] = 199;
    exp_55_ram[3762] = 0;
    exp_55_ram[3763] = 7;
    exp_55_ram[3764] = 0;
    exp_55_ram[3765] = 23;
    exp_55_ram[3766] = 0;
    exp_55_ram[3767] = 39;
    exp_55_ram[3768] = 0;
    exp_55_ram[3769] = 55;
    exp_55_ram[3770] = 0;
    exp_55_ram[3771] = 71;
    exp_55_ram[3772] = 0;
    exp_55_ram[3773] = 86;
    exp_55_ram[3774] = 209;
    exp_55_ram[3775] = 225;
    exp_55_ram[3776] = 241;
    exp_55_ram[3777] = 14;
    exp_55_ram[3778] = 3;
    exp_55_ram[3779] = 5;
    exp_55_ram[3780] = 0;
    exp_55_ram[3781] = 5;
    exp_55_ram[3782] = 79;
    exp_55_ram[3783] = 0;
    exp_55_ram[3784] = 71;
    exp_55_ram[3785] = 79;
    exp_55_ram[3786] = 0;
    exp_55_ram[3787] = 55;
    exp_55_ram[3788] = 7;
    exp_55_ram[3789] = 207;
    exp_55_ram[3790] = 0;
    exp_55_ram[3791] = 71;
    exp_55_ram[3792] = 7;
    exp_55_ram[3793] = 207;
    exp_55_ram[3794] = 0;
    exp_55_ram[3795] = 87;
    exp_55_ram[3796] = 7;
    exp_55_ram[3797] = 207;
    exp_55_ram[3798] = 0;
    exp_55_ram[3799] = 135;
    exp_55_ram[3800] = 143;
    exp_55_ram[3801] = 0;
    exp_55_ram[3802] = 193;
    exp_55_ram[3803] = 129;
    exp_55_ram[3804] = 1;
    exp_55_ram[3805] = 0;
    exp_55_ram[3806] = 1;
    exp_55_ram[3807] = 17;
    exp_55_ram[3808] = 129;
    exp_55_ram[3809] = 1;
    exp_55_ram[3810] = 0;
    exp_55_ram[3811] = 0;
    exp_55_ram[3812] = 71;
    exp_55_ram[3813] = 231;
    exp_55_ram[3814] = 0;
    exp_55_ram[3815] = 0;
    exp_55_ram[3816] = 7;
    exp_55_ram[3817] = 231;
    exp_55_ram[3818] = 0;
    exp_55_ram[3819] = 0;
    exp_55_ram[3820] = 199;
    exp_55_ram[3821] = 231;
    exp_55_ram[3822] = 0;
    exp_55_ram[3823] = 0;
    exp_55_ram[3824] = 199;
    exp_55_ram[3825] = 231;
    exp_55_ram[3826] = 0;
    exp_55_ram[3827] = 16;
    exp_55_ram[3828] = 231;
    exp_55_ram[3829] = 0;
    exp_55_ram[3830] = 16;
    exp_55_ram[3831] = 231;
    exp_55_ram[3832] = 0;
    exp_55_ram[3833] = 16;
    exp_55_ram[3834] = 231;
    exp_55_ram[3835] = 0;
    exp_55_ram[3836] = 16;
    exp_55_ram[3837] = 231;
    exp_55_ram[3838] = 0;
    exp_55_ram[3839] = 16;
    exp_55_ram[3840] = 231;
    exp_55_ram[3841] = 0;
    exp_55_ram[3842] = 16;
    exp_55_ram[3843] = 231;
    exp_55_ram[3844] = 159;
    exp_55_ram[3845] = 0;
    exp_55_ram[3846] = 199;
    exp_55_ram[3847] = 207;
    exp_55_ram[3848] = 0;
    exp_55_ram[3849] = 199;
    exp_55_ram[3850] = 15;
    exp_55_ram[3851] = 0;
    exp_55_ram[3852] = 7;
    exp_55_ram[3853] = 79;
    exp_55_ram[3854] = 0;
    exp_55_ram[3855] = 71;
    exp_55_ram[3856] = 143;
    exp_55_ram[3857] = 0;
    exp_55_ram[3858] = 7;
    exp_55_ram[3859] = 207;
    exp_55_ram[3860] = 0;
    exp_55_ram[3861] = 135;
    exp_55_ram[3862] = 15;
    exp_55_ram[3863] = 0;
    exp_55_ram[3864] = 7;
    exp_55_ram[3865] = 79;
    exp_55_ram[3866] = 4;
    exp_55_ram[3867] = 79;
    exp_55_ram[3868] = 5;
    exp_55_ram[3869] = 244;
    exp_55_ram[3870] = 180;
    exp_55_ram[3871] = 7;
    exp_55_ram[3872] = 207;
    exp_55_ram[3873] = 5;
    exp_55_ram[3874] = 7;
    exp_55_ram[3875] = 196;
    exp_55_ram[3876] = 7;
    exp_55_ram[3877] = 0;
    exp_55_ram[3878] = 7;
    exp_55_ram[3879] = 183;
    exp_55_ram[3880] = 23;
    exp_55_ram[3881] = 7;
    exp_55_ram[3882] = 143;
    exp_55_ram[3883] = 0;
    exp_55_ram[3884] = 7;
    exp_55_ram[3885] = 199;
    exp_55_ram[3886] = 23;
    exp_55_ram[3887] = 7;
    exp_55_ram[3888] = 15;
    exp_55_ram[3889] = 0;
    exp_55_ram[3890] = 7;
    exp_55_ram[3891] = 215;
    exp_55_ram[3892] = 23;
    exp_55_ram[3893] = 7;
    exp_55_ram[3894] = 143;
    exp_55_ram[3895] = 0;
    exp_55_ram[3896] = 199;
    exp_55_ram[3897] = 79;
    exp_55_ram[3898] = 180;
    exp_55_ram[3899] = 7;
    exp_55_ram[3900] = 207;
    exp_55_ram[3901] = 5;
    exp_55_ram[3902] = 247;
    exp_55_ram[3903] = 7;
    exp_55_ram[3904] = 0;
    exp_55_ram[3905] = 7;
    exp_55_ram[3906] = 31;
    exp_55_ram[3907] = 5;
    exp_55_ram[3908] = 7;
    exp_55_ram[3909] = 223;
    exp_55_ram[3910] = 196;
    exp_55_ram[3911] = 96;
    exp_55_ram[3912] = 247;
    exp_55_ram[3913] = 4;
    exp_55_ram[3914] = 160;
    exp_55_ram[3915] = 95;
    exp_55_ram[3916] = 223;
    exp_55_ram[3917] = 196;
    exp_55_ram[3918] = 23;
    exp_55_ram[3919] = 244;
    exp_55_ram[3920] = 223;
    exp_55_ram[3921] = 180;
    exp_55_ram[3922] = 7;
    exp_55_ram[3923] = 144;
    exp_55_ram[3924] = 231;
    exp_55_ram[3925] = 180;
    exp_55_ram[3926] = 16;
    exp_55_ram[3927] = 247;
    exp_55_ram[3928] = 0;
    exp_55_ram[3929] = 7;
    exp_55_ram[3930] = 15;
    exp_55_ram[3931] = 159;
    exp_55_ram[3932] = 5;
    exp_55_ram[3933] = 0;
    exp_55_ram[3934] = 231;
    exp_55_ram[3935] = 159;
    exp_55_ram[3936] = 5;
    exp_55_ram[3937] = 0;
    exp_55_ram[3938] = 231;
    exp_55_ram[3939] = 159;
    exp_55_ram[3940] = 5;
    exp_55_ram[3941] = 0;
    exp_55_ram[3942] = 231;
    exp_55_ram[3943] = 223;
    exp_55_ram[3944] = 4;
    exp_55_ram[3945] = 159;
    exp_55_ram[3946] = 180;
    exp_55_ram[3947] = 32;
    exp_55_ram[3948] = 247;
    exp_55_ram[3949] = 0;
    exp_55_ram[3950] = 7;
    exp_55_ram[3951] = 207;
    exp_55_ram[3952] = 159;
    exp_55_ram[3953] = 5;
    exp_55_ram[3954] = 0;
    exp_55_ram[3955] = 231;
    exp_55_ram[3956] = 159;
    exp_55_ram[3957] = 4;
    exp_55_ram[3958] = 95;
    exp_55_ram[3959] = 180;
    exp_55_ram[3960] = 48;
    exp_55_ram[3961] = 247;
    exp_55_ram[3962] = 0;
    exp_55_ram[3963] = 7;
    exp_55_ram[3964] = 159;
    exp_55_ram[3965] = 223;
    exp_55_ram[3966] = 5;
    exp_55_ram[3967] = 7;
    exp_55_ram[3968] = 0;
    exp_55_ram[3969] = 231;
    exp_55_ram[3970] = 159;
    exp_55_ram[3971] = 5;
    exp_55_ram[3972] = 7;
    exp_55_ram[3973] = 0;
    exp_55_ram[3974] = 231;
    exp_55_ram[3975] = 95;
    exp_55_ram[3976] = 5;
    exp_55_ram[3977] = 7;
    exp_55_ram[3978] = 0;
    exp_55_ram[3979] = 231;
    exp_55_ram[3980] = 159;
    exp_55_ram[3981] = 4;
    exp_55_ram[3982] = 95;
    exp_55_ram[3983] = 180;
    exp_55_ram[3984] = 64;
    exp_55_ram[3985] = 247;
    exp_55_ram[3986] = 0;
    exp_55_ram[3987] = 7;
    exp_55_ram[3988] = 159;
    exp_55_ram[3989] = 223;
    exp_55_ram[3990] = 5;
    exp_55_ram[3991] = 7;
    exp_55_ram[3992] = 0;
    exp_55_ram[3993] = 231;
    exp_55_ram[3994] = 159;
    exp_55_ram[3995] = 5;
    exp_55_ram[3996] = 7;
    exp_55_ram[3997] = 0;
    exp_55_ram[3998] = 231;
    exp_55_ram[3999] = 95;
    exp_55_ram[4000] = 5;
    exp_55_ram[4001] = 7;
    exp_55_ram[4002] = 0;
    exp_55_ram[4003] = 231;
    exp_55_ram[4004] = 159;
    exp_55_ram[4005] = 4;
    exp_55_ram[4006] = 95;
    exp_55_ram[4007] = 5;
    exp_55_ram[4008] = 5;
    exp_55_ram[4009] = 181;
    exp_55_ram[4010] = 1;
    exp_55_ram[4011] = 183;
    exp_55_ram[4012] = 7;
    exp_55_ram[4013] = 5;
    exp_55_ram[4014] = 21;
    exp_55_ram[4015] = 245;
    exp_55_ram[4016] = 1;
    exp_55_ram[4017] = 0;
    exp_55_ram[4018] = 176;
    exp_55_ram[4019] = 245;
    exp_55_ram[4020] = 245;
    exp_55_ram[4021] = 223;
    exp_55_ram[4022] = 250;
    exp_55_ram[4023] = 0;
    exp_55_ram[4024] = 0;
    exp_55_ram[4025] = 0;
    exp_55_ram[4026] = 0;
    exp_55_ram[4027] = 0;
    exp_55_ram[4028] = 0;
    exp_55_ram[4029] = 0;
    exp_55_ram[4030] = 0;
    exp_55_ram[4031] = 0;
    exp_55_ram[4032] = 0;
    exp_55_ram[4033] = 77;
    exp_55_ram[4034] = 68;
    exp_55_ram[4035] = 78;
    exp_55_ram[4036] = 89;
    exp_55_ram[4037] = 83;
    exp_55_ram[4038] = 66;
    exp_55_ram[4039] = 81;
    exp_55_ram[4040] = 68;
    exp_55_ram[4041] = 82;
    exp_55_ram[4042] = 76;
    exp_55_ram[4043] = 77;
    exp_55_ram[4044] = 90;
    exp_55_ram[4045] = 70;
    exp_55_ram[4046] = 69;
    exp_55_ram[4047] = 70;
    exp_55_ram[4048] = 67;
    exp_55_ram[4049] = 88;
    exp_55_ram[4050] = 89;
    exp_55_ram[4051] = 71;
    exp_55_ram[4052] = 85;
    exp_55_ram[4053] = 86;
    exp_55_ram[4054] = 79;
    exp_55_ram[4055] = 74;
    exp_55_ram[4056] = 85;
    exp_55_ram[4057] = 88;
    exp_55_ram[4058] = 84;
    exp_55_ram[4059] = 67;
    exp_55_ram[4060] = 74;
    exp_55_ram[4061] = 66;
    exp_55_ram[4062] = 84;
    exp_55_ram[4063] = 83;
    exp_55_ram[4064] = 76;
    exp_55_ram[4065] = 77;
    exp_55_ram[4066] = 70;
    exp_55_ram[4067] = 90;
    exp_55_ram[4068] = 77;
    exp_55_ram[4069] = 89;
    exp_55_ram[4070] = 87;
    exp_55_ram[4071] = 81;
    exp_55_ram[4072] = 84;
    exp_55_ram[4073] = 75;
    exp_55_ram[4074] = 0;
    exp_55_ram[4075] = 85;
    exp_55_ram[4076] = 76;
    exp_55_ram[4077] = 78;
    exp_55_ram[4078] = 77;
    exp_55_ram[4079] = 70;
    exp_55_ram[4080] = 86;
    exp_55_ram[4081] = 0;
    exp_55_ram[4082] = 80;
    exp_55_ram[4083] = 79;
    exp_55_ram[4084] = 82;
    exp_55_ram[4085] = 71;
    exp_55_ram[4086] = 85;
    exp_55_ram[4087] = 78;
    exp_55_ram[4088] = 0;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_53) begin
      exp_55_ram[exp_49] <= exp_51;
    end
  end
  assign exp_55 = exp_55_ram[exp_50];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_81) begin
        exp_55_ram[exp_77] <= exp_79;
    end
  end
  assign exp_83 = exp_55_ram[exp_78];
  assign exp_82 = exp_96;
  assign exp_96 = 1;
  assign exp_78 = exp_95;
  assign exp_95 = exp_16[31:2];
  assign exp_81 = exp_92;
  assign exp_92 = 0;
  assign exp_77 = exp_91;
  assign exp_91 = 0;
  assign exp_79 = exp_91;
  assign exp_54 = exp_131;
  assign exp_131 = 1;
  assign exp_50 = exp_130;
  assign exp_130 = exp_18[31:2];
  assign exp_53 = exp_119;
  assign exp_119 = exp_117 & exp_118;
  assign exp_117 = exp_22 & exp_23;
  assign exp_118 = exp_24[2:2];
  assign exp_49 = exp_115;
  assign exp_115 = exp_18[31:2];
  assign exp_51 = exp_116;
  assign exp_116 = exp_19[23:16];

  //Create RAM
  reg [7:0] exp_48_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_48_ram[0] = 0;
    exp_48_ram[1] = 1;
    exp_48_ram[2] = 1;
    exp_48_ram[3] = 2;
    exp_48_ram[4] = 2;
    exp_48_ram[5] = 3;
    exp_48_ram[6] = 3;
    exp_48_ram[7] = 4;
    exp_48_ram[8] = 4;
    exp_48_ram[9] = 5;
    exp_48_ram[10] = 5;
    exp_48_ram[11] = 6;
    exp_48_ram[12] = 6;
    exp_48_ram[13] = 7;
    exp_48_ram[14] = 7;
    exp_48_ram[15] = 8;
    exp_48_ram[16] = 8;
    exp_48_ram[17] = 9;
    exp_48_ram[18] = 9;
    exp_48_ram[19] = 10;
    exp_48_ram[20] = 10;
    exp_48_ram[21] = 11;
    exp_48_ram[22] = 11;
    exp_48_ram[23] = 12;
    exp_48_ram[24] = 12;
    exp_48_ram[25] = 13;
    exp_48_ram[26] = 13;
    exp_48_ram[27] = 14;
    exp_48_ram[28] = 14;
    exp_48_ram[29] = 15;
    exp_48_ram[30] = 15;
    exp_48_ram[31] = 81;
    exp_48_ram[32] = 1;
    exp_48_ram[33] = 48;
    exp_48_ram[34] = 0;
    exp_48_ram[35] = 8;
    exp_48_ram[36] = 135;
    exp_48_ram[37] = 8;
    exp_48_ram[38] = 133;
    exp_48_ram[39] = 131;
    exp_48_ram[40] = 148;
    exp_48_ram[41] = 22;
    exp_48_ram[42] = 134;
    exp_48_ram[43] = 246;
    exp_48_ram[44] = 7;
    exp_48_ram[45] = 120;
    exp_48_ram[46] = 7;
    exp_48_ram[47] = 55;
    exp_48_ram[48] = 23;
    exp_48_ram[49] = 85;
    exp_48_ram[50] = 134;
    exp_48_ram[51] = 198;
    exp_48_ram[52] = 5;
    exp_48_ram[53] = 135;
    exp_48_ram[54] = 6;
    exp_48_ram[55] = 12;
    exp_48_ram[56] = 149;
    exp_48_ram[57] = 215;
    exp_48_ram[58] = 24;
    exp_48_ram[59] = 101;
    exp_48_ram[60] = 147;
    exp_48_ram[61] = 88;
    exp_48_ram[62] = 214;
    exp_48_ram[63] = 22;
    exp_48_ram[64] = 86;
    exp_48_ram[65] = 87;
    exp_48_ram[66] = 247;
    exp_48_ram[67] = 133;
    exp_48_ram[68] = 5;
    exp_48_ram[69] = 23;
    exp_48_ram[70] = 103;
    exp_48_ram[71] = 254;
    exp_48_ram[72] = 135;
    exp_48_ram[73] = 133;
    exp_48_ram[74] = 232;
    exp_48_ram[75] = 246;
    exp_48_ram[76] = 133;
    exp_48_ram[77] = 135;
    exp_48_ram[78] = 135;
    exp_48_ram[79] = 247;
    exp_48_ram[80] = 19;
    exp_48_ram[81] = 83;
    exp_48_ram[82] = 215;
    exp_48_ram[83] = 23;
    exp_48_ram[84] = 99;
    exp_48_ram[85] = 6;
    exp_48_ram[86] = 134;
    exp_48_ram[87] = 124;
    exp_48_ram[88] = 3;
    exp_48_ram[89] = 134;
    exp_48_ram[90] = 102;
    exp_48_ram[91] = 116;
    exp_48_ram[92] = 134;
    exp_48_ram[93] = 21;
    exp_48_ram[94] = 101;
    exp_48_ram[95] = 5;
    exp_48_ram[96] = 0;
    exp_48_ram[97] = 5;
    exp_48_ram[98] = 7;
    exp_48_ram[99] = 108;
    exp_48_ram[100] = 7;
    exp_48_ram[101] = 240;
    exp_48_ram[102] = 22;
    exp_48_ram[103] = 7;
    exp_48_ram[104] = 88;
    exp_48_ram[105] = 7;
    exp_48_ram[106] = 112;
    exp_48_ram[107] = 7;
    exp_48_ram[108] = 116;
    exp_48_ram[109] = 5;
    exp_48_ram[110] = 87;
    exp_48_ram[111] = 134;
    exp_48_ram[112] = 199;
    exp_48_ram[113] = 6;
    exp_48_ram[114] = 7;
    exp_48_ram[115] = 6;
    exp_48_ram[116] = 22;
    exp_48_ram[117] = 135;
    exp_48_ram[118] = 5;
    exp_48_ram[119] = 88;
    exp_48_ram[120] = 22;
    exp_48_ram[121] = 86;
    exp_48_ram[122] = 87;
    exp_48_ram[123] = 246;
    exp_48_ram[124] = 215;
    exp_48_ram[125] = 150;
    exp_48_ram[126] = 231;
    exp_48_ram[127] = 14;
    exp_48_ram[128] = 133;
    exp_48_ram[129] = 126;
    exp_48_ram[130] = 7;
    exp_48_ram[131] = 133;
    exp_48_ram[132] = 104;
    exp_48_ram[133] = 118;
    exp_48_ram[134] = 133;
    exp_48_ram[135] = 7;
    exp_48_ram[136] = 7;
    exp_48_ram[137] = 119;
    exp_48_ram[138] = 19;
    exp_48_ram[139] = 83;
    exp_48_ram[140] = 87;
    exp_48_ram[141] = 151;
    exp_48_ram[142] = 227;
    exp_48_ram[143] = 6;
    exp_48_ram[144] = 6;
    exp_48_ram[145] = 124;
    exp_48_ram[146] = 3;
    exp_48_ram[147] = 6;
    exp_48_ram[148] = 102;
    exp_48_ram[149] = 116;
    exp_48_ram[150] = 6;
    exp_48_ram[151] = 21;
    exp_48_ram[152] = 101;
    exp_48_ram[153] = 128;
    exp_48_ram[154] = 7;
    exp_48_ram[155] = 5;
    exp_48_ram[156] = 100;
    exp_48_ram[157] = 5;
    exp_48_ram[158] = 240;
    exp_48_ram[159] = 24;
    exp_48_ram[160] = 213;
    exp_48_ram[161] = 147;
    exp_48_ram[162] = 151;
    exp_48_ram[163] = 215;
    exp_48_ram[164] = 88;
    exp_48_ram[165] = 102;
    exp_48_ram[166] = 119;
    exp_48_ram[167] = 23;
    exp_48_ram[168] = 215;
    exp_48_ram[169] = 85;
    exp_48_ram[170] = 85;
    exp_48_ram[171] = 23;
    exp_48_ram[172] = 103;
    exp_48_ram[173] = 134;
    exp_48_ram[174] = 5;
    exp_48_ram[175] = 126;
    exp_48_ram[176] = 7;
    exp_48_ram[177] = 5;
    exp_48_ram[178] = 104;
    exp_48_ram[179] = 118;
    exp_48_ram[180] = 5;
    exp_48_ram[181] = 7;
    exp_48_ram[182] = 6;
    exp_48_ram[183] = 247;
    exp_48_ram[184] = 22;
    exp_48_ram[185] = 86;
    exp_48_ram[186] = 214;
    exp_48_ram[187] = 23;
    exp_48_ram[188] = 133;
    exp_48_ram[189] = 103;
    exp_48_ram[190] = 135;
    exp_48_ram[191] = 254;
    exp_48_ram[192] = 135;
    exp_48_ram[193] = 135;
    exp_48_ram[194] = 232;
    exp_48_ram[195] = 246;
    exp_48_ram[196] = 135;
    exp_48_ram[197] = 135;
    exp_48_ram[198] = 149;
    exp_48_ram[199] = 135;
    exp_48_ram[200] = 229;
    exp_48_ram[201] = 240;
    exp_48_ram[202] = 230;
    exp_48_ram[203] = 7;
    exp_48_ram[204] = 244;
    exp_48_ram[205] = 7;
    exp_48_ram[206] = 53;
    exp_48_ram[207] = 149;
    exp_48_ram[208] = 23;
    exp_48_ram[209] = 213;
    exp_48_ram[210] = 7;
    exp_48_ram[211] = 7;
    exp_48_ram[212] = 71;
    exp_48_ram[213] = 5;
    exp_48_ram[214] = 7;
    exp_48_ram[215] = 5;
    exp_48_ram[216] = 22;
    exp_48_ram[217] = 5;
    exp_48_ram[218] = 238;
    exp_48_ram[219] = 181;
    exp_48_ram[220] = 69;
    exp_48_ram[221] = 240;
    exp_48_ram[222] = 7;
    exp_48_ram[223] = 5;
    exp_48_ram[224] = 224;
    exp_48_ram[225] = 5;
    exp_48_ram[226] = 240;
    exp_48_ram[227] = 88;
    exp_48_ram[228] = 150;
    exp_48_ram[229] = 104;
    exp_48_ram[230] = 222;
    exp_48_ram[231] = 94;
    exp_48_ram[232] = 118;
    exp_48_ram[233] = 151;
    exp_48_ram[234] = 215;
    exp_48_ram[235] = 19;
    exp_48_ram[236] = 102;
    exp_48_ram[237] = 23;
    exp_48_ram[238] = 215;
    exp_48_ram[239] = 87;
    exp_48_ram[240] = 94;
    exp_48_ram[241] = 150;
    exp_48_ram[242] = 231;
    exp_48_ram[243] = 143;
    exp_48_ram[244] = 5;
    exp_48_ram[245] = 126;
    exp_48_ram[246] = 7;
    exp_48_ram[247] = 5;
    exp_48_ram[248] = 104;
    exp_48_ram[249] = 118;
    exp_48_ram[250] = 5;
    exp_48_ram[251] = 7;
    exp_48_ram[252] = 7;
    exp_48_ram[253] = 118;
    exp_48_ram[254] = 87;
    exp_48_ram[255] = 150;
    exp_48_ram[256] = 142;
    exp_48_ram[257] = 23;
    exp_48_ram[258] = 215;
    exp_48_ram[259] = 231;
    exp_48_ram[260] = 6;
    exp_48_ram[261] = 254;
    exp_48_ram[262] = 135;
    exp_48_ram[263] = 6;
    exp_48_ram[264] = 232;
    exp_48_ram[265] = 246;
    exp_48_ram[266] = 6;
    exp_48_ram[267] = 135;
    exp_48_ram[268] = 21;
    exp_48_ram[269] = 14;
    exp_48_ram[270] = 101;
    exp_48_ram[271] = 134;
    exp_48_ram[272] = 120;
    exp_48_ram[273] = 86;
    exp_48_ram[274] = 118;
    exp_48_ram[275] = 83;
    exp_48_ram[276] = 135;
    exp_48_ram[277] = 14;
    exp_48_ram[278] = 6;
    exp_48_ram[279] = 87;
    exp_48_ram[280] = 8;
    exp_48_ram[281] = 8;
    exp_48_ram[282] = 7;
    exp_48_ram[283] = 6;
    exp_48_ram[284] = 116;
    exp_48_ram[285] = 6;
    exp_48_ram[286] = 86;
    exp_48_ram[287] = 134;
    exp_48_ram[288] = 230;
    exp_48_ram[289] = 156;
    exp_48_ram[290] = 7;
    exp_48_ram[291] = 135;
    exp_48_ram[292] = 119;
    exp_48_ram[293] = 23;
    exp_48_ram[294] = 126;
    exp_48_ram[295] = 152;
    exp_48_ram[296] = 7;
    exp_48_ram[297] = 5;
    exp_48_ram[298] = 254;
    exp_48_ram[299] = 5;
    exp_48_ram[300] = 240;
    exp_48_ram[301] = 5;
    exp_48_ram[302] = 5;
    exp_48_ram[303] = 240;
    exp_48_ram[304] = 7;
    exp_48_ram[305] = 7;
    exp_48_ram[306] = 216;
    exp_48_ram[307] = 120;
    exp_48_ram[308] = 7;
    exp_48_ram[309] = 3;
    exp_48_ram[310] = 120;
    exp_48_ram[311] = 213;
    exp_48_ram[312] = 14;
    exp_48_ram[313] = 213;
    exp_48_ram[314] = 119;
    exp_48_ram[315] = 14;
    exp_48_ram[316] = 245;
    exp_48_ram[317] = 214;
    exp_48_ram[318] = 26;
    exp_48_ram[319] = 238;
    exp_48_ram[320] = 138;
    exp_48_ram[321] = 5;
    exp_48_ram[322] = 128;
    exp_48_ram[323] = 150;
    exp_48_ram[324] = 110;
    exp_48_ram[325] = 152;
    exp_48_ram[326] = 16;
    exp_48_ram[327] = 231;
    exp_48_ram[328] = 183;
    exp_48_ram[329] = 150;
    exp_48_ram[330] = 102;
    exp_48_ram[331] = 12;
    exp_48_ram[332] = 156;
    exp_48_ram[333] = 20;
    exp_48_ram[334] = 208;
    exp_48_ram[335] = 0;
    exp_48_ram[336] = 5;
    exp_48_ram[337] = 128;
    exp_48_ram[338] = 5;
    exp_48_ram[339] = 138;
    exp_48_ram[340] = 133;
    exp_48_ram[341] = 128;
    exp_48_ram[342] = 86;
    exp_48_ram[343] = 2;
    exp_48_ram[344] = 128;
    exp_48_ram[345] = 108;
    exp_48_ram[346] = 146;
    exp_48_ram[347] = 104;
    exp_48_ram[348] = 102;
    exp_48_ram[349] = 5;
    exp_48_ram[350] = 128;
    exp_48_ram[351] = 5;
    exp_48_ram[352] = 128;
    exp_48_ram[353] = 152;
    exp_48_ram[354] = 240;
    exp_48_ram[355] = 232;
    exp_48_ram[356] = 240;
    exp_48_ram[357] = 142;
    exp_48_ram[358] = 158;
    exp_48_ram[359] = 7;
    exp_48_ram[360] = 240;
    exp_48_ram[361] = 1;
    exp_48_ram[362] = 36;
    exp_48_ram[363] = 38;
    exp_48_ram[364] = 4;
    exp_48_ram[365] = 2;
    exp_48_ram[366] = 0;
    exp_48_ram[367] = 7;
    exp_48_ram[368] = 7;
    exp_48_ram[369] = 7;
    exp_48_ram[370] = 192;
    exp_48_ram[371] = 7;
    exp_48_ram[372] = 135;
    exp_48_ram[373] = 5;
    exp_48_ram[374] = 87;
    exp_48_ram[375] = 20;
    exp_48_ram[376] = 32;
    exp_48_ram[377] = 5;
    exp_48_ram[378] = 151;
    exp_48_ram[379] = 36;
    exp_48_ram[380] = 23;
    exp_48_ram[381] = 215;
    exp_48_ram[382] = 102;
    exp_48_ram[383] = 133;
    exp_48_ram[384] = 1;
    exp_48_ram[385] = 128;
    exp_48_ram[386] = 7;
    exp_48_ram[387] = 23;
    exp_48_ram[388] = 4;
    exp_48_ram[389] = 240;
    exp_48_ram[390] = 7;
    exp_48_ram[391] = 7;
    exp_48_ram[392] = 240;
    exp_48_ram[393] = 1;
    exp_48_ram[394] = 46;
    exp_48_ram[395] = 44;
    exp_48_ram[396] = 42;
    exp_48_ram[397] = 40;
    exp_48_ram[398] = 38;
    exp_48_ram[399] = 36;
    exp_48_ram[400] = 103;
    exp_48_ram[401] = 140;
    exp_48_ram[402] = 4;
    exp_48_ram[403] = 137;
    exp_48_ram[404] = 132;
    exp_48_ram[405] = 132;
    exp_48_ram[406] = 133;
    exp_48_ram[407] = 0;
    exp_48_ram[408] = 9;
    exp_48_ram[409] = 10;
    exp_48_ram[410] = 10;
    exp_48_ram[411] = 7;
    exp_48_ram[412] = 196;
    exp_48_ram[413] = 7;
    exp_48_ram[414] = 7;
    exp_48_ram[415] = 84;
    exp_48_ram[416] = 7;
    exp_48_ram[417] = 66;
    exp_48_ram[418] = 4;
    exp_48_ram[419] = 135;
    exp_48_ram[420] = 132;
    exp_48_ram[421] = 84;
    exp_48_ram[422] = 21;
    exp_48_ram[423] = 228;
    exp_48_ram[424] = 23;
    exp_48_ram[425] = 32;
    exp_48_ram[426] = 36;
    exp_48_ram[427] = 149;
    exp_48_ram[428] = 26;
    exp_48_ram[429] = 213;
    exp_48_ram[430] = 103;
    exp_48_ram[431] = 36;
    exp_48_ram[432] = 41;
    exp_48_ram[433] = 41;
    exp_48_ram[434] = 42;
    exp_48_ram[435] = 133;
    exp_48_ram[436] = 5;
    exp_48_ram[437] = 1;
    exp_48_ram[438] = 128;
    exp_48_ram[439] = 0;
    exp_48_ram[440] = 9;
    exp_48_ram[441] = 240;
    exp_48_ram[442] = 133;
    exp_48_ram[443] = 20;
    exp_48_ram[444] = 7;
    exp_48_ram[445] = 240;
    exp_48_ram[446] = 7;
    exp_48_ram[447] = 220;
    exp_48_ram[448] = 134;
    exp_48_ram[449] = 5;
    exp_48_ram[450] = 5;
    exp_48_ram[451] = 0;
    exp_48_ram[452] = 101;
    exp_48_ram[453] = 6;
    exp_48_ram[454] = 52;
    exp_48_ram[455] = 5;
    exp_48_ram[456] = 5;
    exp_48_ram[457] = 6;
    exp_48_ram[458] = 0;
    exp_48_ram[459] = 228;
    exp_48_ram[460] = 137;
    exp_48_ram[461] = 7;
    exp_48_ram[462] = 7;
    exp_48_ram[463] = 5;
    exp_48_ram[464] = 84;
    exp_48_ram[465] = 7;
    exp_48_ram[466] = 66;
    exp_48_ram[467] = 135;
    exp_48_ram[468] = 21;
    exp_48_ram[469] = 9;
    exp_48_ram[470] = 9;
    exp_48_ram[471] = 89;
    exp_48_ram[472] = 101;
    exp_48_ram[473] = 23;
    exp_48_ram[474] = 7;
    exp_48_ram[475] = 7;
    exp_48_ram[476] = 245;
    exp_48_ram[477] = 247;
    exp_48_ram[478] = 0;
    exp_48_ram[479] = 247;
    exp_48_ram[480] = 6;
    exp_48_ram[481] = 10;
    exp_48_ram[482] = 135;
    exp_48_ram[483] = 55;
    exp_48_ram[484] = 133;
    exp_48_ram[485] = 7;
    exp_48_ram[486] = 7;
    exp_48_ram[487] = 247;
    exp_48_ram[488] = 12;
    exp_48_ram[489] = 7;
    exp_48_ram[490] = 7;
    exp_48_ram[491] = 10;
    exp_48_ram[492] = 245;
    exp_48_ram[493] = 10;
    exp_48_ram[494] = 215;
    exp_48_ram[495] = 149;
    exp_48_ram[496] = 103;
    exp_48_ram[497] = 212;
    exp_48_ram[498] = 240;
    exp_48_ram[499] = 133;
    exp_48_ram[500] = 21;
    exp_48_ram[501] = 7;
    exp_48_ram[502] = 240;
    exp_48_ram[503] = 4;
    exp_48_ram[504] = 7;
    exp_48_ram[505] = 10;
    exp_48_ram[506] = 240;
    exp_48_ram[507] = 0;
    exp_48_ram[508] = 7;
    exp_48_ram[509] = 135;
    exp_48_ram[510] = 76;
    exp_48_ram[511] = 5;
    exp_48_ram[512] = 7;
    exp_48_ram[513] = 213;
    exp_48_ram[514] = 5;
    exp_48_ram[515] = 128;
    exp_48_ram[516] = 215;
    exp_48_ram[517] = 85;
    exp_48_ram[518] = 149;
    exp_48_ram[519] = 101;
    exp_48_ram[520] = 240;
    exp_48_ram[521] = 0;
    exp_48_ram[522] = 7;
    exp_48_ram[523] = 135;
    exp_48_ram[524] = 76;
    exp_48_ram[525] = 5;
    exp_48_ram[526] = 7;
    exp_48_ram[527] = 21;
    exp_48_ram[528] = 5;
    exp_48_ram[529] = 128;
    exp_48_ram[530] = 23;
    exp_48_ram[531] = 149;
    exp_48_ram[532] = 85;
    exp_48_ram[533] = 229;
    exp_48_ram[534] = 240;
    exp_48_ram[535] = 7;
    exp_48_ram[536] = 122;
    exp_48_ram[537] = 7;
    exp_48_ram[538] = 183;
    exp_48_ram[539] = 151;
    exp_48_ram[540] = 23;
    exp_48_ram[541] = 6;
    exp_48_ram[542] = 134;
    exp_48_ram[543] = 85;
    exp_48_ram[544] = 7;
    exp_48_ram[545] = 133;
    exp_48_ram[546] = 69;
    exp_48_ram[547] = 133;
    exp_48_ram[548] = 128;
    exp_48_ram[549] = 7;
    exp_48_ram[550] = 7;
    exp_48_ram[551] = 106;
    exp_48_ram[552] = 7;
    exp_48_ram[553] = 240;
    exp_48_ram[554] = 117;
    exp_48_ram[555] = 110;
    exp_48_ram[556] = 87;
    exp_48_ram[557] = 104;
    exp_48_ram[558] = 105;
    exp_48_ram[559] = 0;
    exp_48_ram[560] = 97;
    exp_48_ram[561] = 98;
    exp_48_ram[562] = 65;
    exp_48_ram[563] = 97;
    exp_48_ram[564] = 110;
    exp_48_ram[565] = 65;
    exp_48_ram[566] = 101;
    exp_48_ram[567] = 116;
    exp_48_ram[568] = 68;
    exp_48_ram[569] = 0;
    exp_48_ram[570] = 101;
    exp_48_ram[571] = 32;
    exp_48_ram[572] = 108;
    exp_48_ram[573] = 0;
    exp_48_ram[574] = 117;
    exp_48_ram[575] = 110;
    exp_48_ram[576] = 110;
    exp_48_ram[577] = 116;
    exp_48_ram[578] = 100;
    exp_48_ram[579] = 100;
    exp_48_ram[580] = 46;
    exp_48_ram[581] = 0;
    exp_48_ram[582] = 117;
    exp_48_ram[583] = 110;
    exp_48_ram[584] = 87;
    exp_48_ram[585] = 101;
    exp_48_ram[586] = 46;
    exp_48_ram[587] = 51;
    exp_48_ram[588] = 105;
    exp_48_ram[589] = 110;
    exp_48_ram[590] = 101;
    exp_48_ram[591] = 117;
    exp_48_ram[592] = 112;
    exp_48_ram[593] = 115;
    exp_48_ram[594] = 32;
    exp_48_ram[595] = 101;
    exp_48_ram[596] = 100;
    exp_48_ram[597] = 54;
    exp_48_ram[598] = 105;
    exp_48_ram[599] = 110;
    exp_48_ram[600] = 101;
    exp_48_ram[601] = 117;
    exp_48_ram[602] = 112;
    exp_48_ram[603] = 115;
    exp_48_ram[604] = 32;
    exp_48_ram[605] = 101;
    exp_48_ram[606] = 100;
    exp_48_ram[607] = 51;
    exp_48_ram[608] = 105;
    exp_48_ram[609] = 110;
    exp_48_ram[610] = 101;
    exp_48_ram[611] = 105;
    exp_48_ram[612] = 101;
    exp_48_ram[613] = 110;
    exp_48_ram[614] = 115;
    exp_48_ram[615] = 110;
    exp_48_ram[616] = 54;
    exp_48_ram[617] = 105;
    exp_48_ram[618] = 110;
    exp_48_ram[619] = 101;
    exp_48_ram[620] = 105;
    exp_48_ram[621] = 101;
    exp_48_ram[622] = 110;
    exp_48_ram[623] = 115;
    exp_48_ram[624] = 110;
    exp_48_ram[625] = 101;
    exp_48_ram[626] = 0;
    exp_48_ram[627] = 111;
    exp_48_ram[628] = 58;
    exp_48_ram[629] = 97;
    exp_48_ram[630] = 0;
    exp_48_ram[631] = 111;
    exp_48_ram[632] = 0;
    exp_48_ram[633] = 105;
    exp_48_ram[634] = 101;
    exp_48_ram[635] = 67;
    exp_48_ram[636] = 115;
    exp_48_ram[637] = 68;
    exp_48_ram[638] = 0;
    exp_48_ram[639] = 97;
    exp_48_ram[640] = 101;
    exp_48_ram[641] = 32;
    exp_48_ram[642] = 108;
    exp_48_ram[643] = 41;
    exp_48_ram[644] = 105;
    exp_48_ram[645] = 32;
    exp_48_ram[646] = 101;
    exp_48_ram[647] = 41;
    exp_48_ram[648] = 115;
    exp_48_ram[649] = 117;
    exp_48_ram[650] = 112;
    exp_48_ram[651] = 97;
    exp_48_ram[652] = 110;
    exp_48_ram[653] = 41;
    exp_48_ram[654] = 108;
    exp_48_ram[655] = 108;
    exp_48_ram[656] = 0;
    exp_48_ram[657] = 41;
    exp_48_ram[658] = 105;
    exp_48_ram[659] = 32;
    exp_48_ram[660] = 104;
    exp_48_ram[661] = 0;
    exp_48_ram[662] = 41;
    exp_48_ram[663] = 77;
    exp_48_ram[664] = 109;
    exp_48_ram[665] = 111;
    exp_48_ram[666] = 32;
    exp_48_ram[667] = 105;
    exp_48_ram[668] = 110;
    exp_48_ram[669] = 0;
    exp_48_ram[670] = 0;
    exp_48_ram[671] = 110;
    exp_48_ram[672] = 97;
    exp_48_ram[673] = 99;
    exp_48_ram[674] = 101;
    exp_48_ram[675] = 61;
    exp_48_ram[676] = 61;
    exp_48_ram[677] = 61;
    exp_48_ram[678] = 61;
    exp_48_ram[679] = 0;
    exp_48_ram[680] = 46;
    exp_48_ram[681] = 101;
    exp_48_ram[682] = 115;
    exp_48_ram[683] = 105;
    exp_48_ram[684] = 32;
    exp_48_ram[685] = 108;
    exp_48_ram[686] = 108;
    exp_48_ram[687] = 41;
    exp_48_ram[688] = 45;
    exp_48_ram[689] = 32;
    exp_48_ram[690] = 116;
    exp_48_ram[691] = 105;
    exp_48_ram[692] = 101;
    exp_48_ram[693] = 105;
    exp_48_ram[694] = 32;
    exp_48_ram[695] = 46;
    exp_48_ram[696] = 51;
    exp_48_ram[697] = 46;
    exp_48_ram[698] = 102;
    exp_48_ram[699] = 116;
    exp_48_ram[700] = 40;
    exp_48_ram[701] = 99;
    exp_48_ram[702] = 46;
    exp_48_ram[703] = 98;
    exp_48_ram[704] = 46;
    exp_48_ram[705] = 110;
    exp_48_ram[706] = 101;
    exp_48_ram[707] = 110;
    exp_48_ram[708] = 40;
    exp_48_ram[709] = 103;
    exp_48_ram[710] = 108;
    exp_48_ram[711] = 103;
    exp_48_ram[712] = 97;
    exp_48_ram[713] = 41;
    exp_48_ram[714] = 102;
    exp_48_ram[715] = 109;
    exp_48_ram[716] = 108;
    exp_48_ram[717] = 114;
    exp_48_ram[718] = 116;
    exp_48_ram[719] = 103;
    exp_48_ram[720] = 97;
    exp_48_ram[721] = 0;
    exp_48_ram[722] = 46;
    exp_48_ram[723] = 116;
    exp_48_ram[724] = 112;
    exp_48_ram[725] = 116;
    exp_48_ram[726] = 115;
    exp_48_ram[727] = 45;
    exp_48_ram[728] = 32;
    exp_48_ram[729] = 116;
    exp_48_ram[730] = 105;
    exp_48_ram[731] = 101;
    exp_48_ram[732] = 105;
    exp_48_ram[733] = 32;
    exp_48_ram[734] = 46;
    exp_48_ram[735] = 97;
    exp_48_ram[736] = 101;
    exp_48_ram[737] = 32;
    exp_48_ram[738] = 10;
    exp_48_ram[739] = 32;
    exp_48_ram[740] = 62;
    exp_48_ram[741] = 1;
    exp_48_ram[742] = 3;
    exp_48_ram[743] = 4;
    exp_48_ram[744] = 4;
    exp_48_ram[745] = 5;
    exp_48_ram[746] = 5;
    exp_48_ram[747] = 5;
    exp_48_ram[748] = 5;
    exp_48_ram[749] = 6;
    exp_48_ram[750] = 6;
    exp_48_ram[751] = 6;
    exp_48_ram[752] = 6;
    exp_48_ram[753] = 6;
    exp_48_ram[754] = 6;
    exp_48_ram[755] = 6;
    exp_48_ram[756] = 6;
    exp_48_ram[757] = 7;
    exp_48_ram[758] = 7;
    exp_48_ram[759] = 7;
    exp_48_ram[760] = 7;
    exp_48_ram[761] = 7;
    exp_48_ram[762] = 7;
    exp_48_ram[763] = 7;
    exp_48_ram[764] = 7;
    exp_48_ram[765] = 7;
    exp_48_ram[766] = 7;
    exp_48_ram[767] = 7;
    exp_48_ram[768] = 7;
    exp_48_ram[769] = 7;
    exp_48_ram[770] = 7;
    exp_48_ram[771] = 7;
    exp_48_ram[772] = 7;
    exp_48_ram[773] = 8;
    exp_48_ram[774] = 8;
    exp_48_ram[775] = 8;
    exp_48_ram[776] = 8;
    exp_48_ram[777] = 8;
    exp_48_ram[778] = 8;
    exp_48_ram[779] = 8;
    exp_48_ram[780] = 8;
    exp_48_ram[781] = 8;
    exp_48_ram[782] = 8;
    exp_48_ram[783] = 8;
    exp_48_ram[784] = 8;
    exp_48_ram[785] = 8;
    exp_48_ram[786] = 8;
    exp_48_ram[787] = 8;
    exp_48_ram[788] = 8;
    exp_48_ram[789] = 8;
    exp_48_ram[790] = 8;
    exp_48_ram[791] = 8;
    exp_48_ram[792] = 8;
    exp_48_ram[793] = 8;
    exp_48_ram[794] = 8;
    exp_48_ram[795] = 8;
    exp_48_ram[796] = 8;
    exp_48_ram[797] = 8;
    exp_48_ram[798] = 8;
    exp_48_ram[799] = 8;
    exp_48_ram[800] = 8;
    exp_48_ram[801] = 8;
    exp_48_ram[802] = 8;
    exp_48_ram[803] = 8;
    exp_48_ram[804] = 8;
    exp_48_ram[805] = 1;
    exp_48_ram[806] = 38;
    exp_48_ram[807] = 4;
    exp_48_ram[808] = 46;
    exp_48_ram[809] = 39;
    exp_48_ram[810] = 38;
    exp_48_ram[811] = 39;
    exp_48_ram[812] = 167;
    exp_48_ram[813] = 133;
    exp_48_ram[814] = 36;
    exp_48_ram[815] = 1;
    exp_48_ram[816] = 128;
    exp_48_ram[817] = 1;
    exp_48_ram[818] = 38;
    exp_48_ram[819] = 4;
    exp_48_ram[820] = 46;
    exp_48_ram[821] = 44;
    exp_48_ram[822] = 39;
    exp_48_ram[823] = 38;
    exp_48_ram[824] = 39;
    exp_48_ram[825] = 39;
    exp_48_ram[826] = 160;
    exp_48_ram[827] = 39;
    exp_48_ram[828] = 133;
    exp_48_ram[829] = 36;
    exp_48_ram[830] = 1;
    exp_48_ram[831] = 128;
    exp_48_ram[832] = 1;
    exp_48_ram[833] = 46;
    exp_48_ram[834] = 44;
    exp_48_ram[835] = 4;
    exp_48_ram[836] = 38;
    exp_48_ram[837] = 71;
    exp_48_ram[838] = 167;
    exp_48_ram[839] = 133;
    exp_48_ram[840] = 37;
    exp_48_ram[841] = 240;
    exp_48_ram[842] = 7;
    exp_48_ram[843] = 133;
    exp_48_ram[844] = 32;
    exp_48_ram[845] = 36;
    exp_48_ram[846] = 1;
    exp_48_ram[847] = 128;
    exp_48_ram[848] = 1;
    exp_48_ram[849] = 38;
    exp_48_ram[850] = 36;
    exp_48_ram[851] = 4;
    exp_48_ram[852] = 71;
    exp_48_ram[853] = 167;
    exp_48_ram[854] = 133;
    exp_48_ram[855] = 240;
    exp_48_ram[856] = 7;
    exp_48_ram[857] = 133;
    exp_48_ram[858] = 32;
    exp_48_ram[859] = 36;
    exp_48_ram[860] = 1;
    exp_48_ram[861] = 128;
    exp_48_ram[862] = 1;
    exp_48_ram[863] = 38;
    exp_48_ram[864] = 36;
    exp_48_ram[865] = 4;
    exp_48_ram[866] = 46;
    exp_48_ram[867] = 44;
    exp_48_ram[868] = 38;
    exp_48_ram[869] = 0;
    exp_48_ram[870] = 39;
    exp_48_ram[871] = 135;
    exp_48_ram[872] = 38;
    exp_48_ram[873] = 39;
    exp_48_ram[874] = 7;
    exp_48_ram[875] = 199;
    exp_48_ram[876] = 37;
    exp_48_ram[877] = 133;
    exp_48_ram[878] = 240;
    exp_48_ram[879] = 39;
    exp_48_ram[880] = 39;
    exp_48_ram[881] = 7;
    exp_48_ram[882] = 199;
    exp_48_ram[883] = 150;
    exp_48_ram[884] = 39;
    exp_48_ram[885] = 133;
    exp_48_ram[886] = 32;
    exp_48_ram[887] = 36;
    exp_48_ram[888] = 1;
    exp_48_ram[889] = 128;
    exp_48_ram[890] = 1;
    exp_48_ram[891] = 46;
    exp_48_ram[892] = 44;
    exp_48_ram[893] = 4;
    exp_48_ram[894] = 38;
    exp_48_ram[895] = 71;
    exp_48_ram[896] = 167;
    exp_48_ram[897] = 133;
    exp_48_ram[898] = 37;
    exp_48_ram[899] = 240;
    exp_48_ram[900] = 71;
    exp_48_ram[901] = 167;
    exp_48_ram[902] = 133;
    exp_48_ram[903] = 5;
    exp_48_ram[904] = 240;
    exp_48_ram[905] = 7;
    exp_48_ram[906] = 133;
    exp_48_ram[907] = 32;
    exp_48_ram[908] = 36;
    exp_48_ram[909] = 1;
    exp_48_ram[910] = 128;
    exp_48_ram[911] = 1;
    exp_48_ram[912] = 46;
    exp_48_ram[913] = 4;
    exp_48_ram[914] = 38;
    exp_48_ram[915] = 39;
    exp_48_ram[916] = 7;
    exp_48_ram[917] = 216;
    exp_48_ram[918] = 39;
    exp_48_ram[919] = 7;
    exp_48_ram[920] = 222;
    exp_48_ram[921] = 39;
    exp_48_ram[922] = 7;
    exp_48_ram[923] = 220;
    exp_48_ram[924] = 39;
    exp_48_ram[925] = 7;
    exp_48_ram[926] = 198;
    exp_48_ram[927] = 7;
    exp_48_ram[928] = 0;
    exp_48_ram[929] = 7;
    exp_48_ram[930] = 133;
    exp_48_ram[931] = 36;
    exp_48_ram[932] = 1;
    exp_48_ram[933] = 128;
    exp_48_ram[934] = 1;
    exp_48_ram[935] = 46;
    exp_48_ram[936] = 4;
    exp_48_ram[937] = 38;
    exp_48_ram[938] = 39;
    exp_48_ram[939] = 7;
    exp_48_ram[940] = 220;
    exp_48_ram[941] = 39;
    exp_48_ram[942] = 7;
    exp_48_ram[943] = 198;
    exp_48_ram[944] = 7;
    exp_48_ram[945] = 0;
    exp_48_ram[946] = 7;
    exp_48_ram[947] = 133;
    exp_48_ram[948] = 36;
    exp_48_ram[949] = 1;
    exp_48_ram[950] = 128;
    exp_48_ram[951] = 1;
    exp_48_ram[952] = 46;
    exp_48_ram[953] = 44;
    exp_48_ram[954] = 4;
    exp_48_ram[955] = 38;
    exp_48_ram[956] = 37;
    exp_48_ram[957] = 240;
    exp_48_ram[958] = 7;
    exp_48_ram[959] = 136;
    exp_48_ram[960] = 39;
    exp_48_ram[961] = 135;
    exp_48_ram[962] = 0;
    exp_48_ram[963] = 39;
    exp_48_ram[964] = 133;
    exp_48_ram[965] = 32;
    exp_48_ram[966] = 36;
    exp_48_ram[967] = 1;
    exp_48_ram[968] = 128;
    exp_48_ram[969] = 1;
    exp_48_ram[970] = 46;
    exp_48_ram[971] = 44;
    exp_48_ram[972] = 42;
    exp_48_ram[973] = 4;
    exp_48_ram[974] = 4;
    exp_48_ram[975] = 167;
    exp_48_ram[976] = 36;
    exp_48_ram[977] = 7;
    exp_48_ram[978] = 34;
    exp_48_ram[979] = 7;
    exp_48_ram[980] = 32;
    exp_48_ram[981] = 7;
    exp_48_ram[982] = 46;
    exp_48_ram[983] = 44;
    exp_48_ram[984] = 42;
    exp_48_ram[985] = 42;
    exp_48_ram[986] = 35;
    exp_48_ram[987] = 40;
    exp_48_ram[988] = 40;
    exp_48_ram[989] = 37;
    exp_48_ram[990] = 37;
    exp_48_ram[991] = 38;
    exp_48_ram[992] = 38;
    exp_48_ram[993] = 39;
    exp_48_ram[994] = 39;
    exp_48_ram[995] = 32;
    exp_48_ram[996] = 34;
    exp_48_ram[997] = 36;
    exp_48_ram[998] = 38;
    exp_48_ram[999] = 40;
    exp_48_ram[1000] = 42;
    exp_48_ram[1001] = 44;
    exp_48_ram[1002] = 46;
    exp_48_ram[1003] = 32;
    exp_48_ram[1004] = 7;
    exp_48_ram[1005] = 133;
    exp_48_ram[1006] = 0;
    exp_48_ram[1007] = 36;
    exp_48_ram[1008] = 38;
    exp_48_ram[1009] = 7;
    exp_48_ram[1010] = 37;
    exp_48_ram[1011] = 38;
    exp_48_ram[1012] = 133;
    exp_48_ram[1013] = 16;
    exp_48_ram[1014] = 39;
    exp_48_ram[1015] = 39;
    exp_48_ram[1016] = 7;
    exp_48_ram[1017] = 32;
    exp_48_ram[1018] = 35;
    exp_48_ram[1019] = 40;
    exp_48_ram[1020] = 40;
    exp_48_ram[1021] = 37;
    exp_48_ram[1022] = 37;
    exp_48_ram[1023] = 38;
    exp_48_ram[1024] = 38;
    exp_48_ram[1025] = 39;
    exp_48_ram[1026] = 39;
    exp_48_ram[1027] = 32;
    exp_48_ram[1028] = 34;
    exp_48_ram[1029] = 36;
    exp_48_ram[1030] = 38;
    exp_48_ram[1031] = 40;
    exp_48_ram[1032] = 42;
    exp_48_ram[1033] = 44;
    exp_48_ram[1034] = 46;
    exp_48_ram[1035] = 32;
    exp_48_ram[1036] = 7;
    exp_48_ram[1037] = 133;
    exp_48_ram[1038] = 0;
    exp_48_ram[1039] = 36;
    exp_48_ram[1040] = 38;
    exp_48_ram[1041] = 167;
    exp_48_ram[1042] = 34;
    exp_48_ram[1043] = 7;
    exp_48_ram[1044] = 32;
    exp_48_ram[1045] = 7;
    exp_48_ram[1046] = 46;
    exp_48_ram[1047] = 7;
    exp_48_ram[1048] = 44;
    exp_48_ram[1049] = 42;
    exp_48_ram[1050] = 40;
    exp_48_ram[1051] = 42;
    exp_48_ram[1052] = 35;
    exp_48_ram[1053] = 40;
    exp_48_ram[1054] = 40;
    exp_48_ram[1055] = 37;
    exp_48_ram[1056] = 37;
    exp_48_ram[1057] = 38;
    exp_48_ram[1058] = 38;
    exp_48_ram[1059] = 39;
    exp_48_ram[1060] = 39;
    exp_48_ram[1061] = 32;
    exp_48_ram[1062] = 34;
    exp_48_ram[1063] = 36;
    exp_48_ram[1064] = 38;
    exp_48_ram[1065] = 40;
    exp_48_ram[1066] = 42;
    exp_48_ram[1067] = 44;
    exp_48_ram[1068] = 46;
    exp_48_ram[1069] = 32;
    exp_48_ram[1070] = 7;
    exp_48_ram[1071] = 133;
    exp_48_ram[1072] = 0;
    exp_48_ram[1073] = 32;
    exp_48_ram[1074] = 34;
    exp_48_ram[1075] = 7;
    exp_48_ram[1076] = 37;
    exp_48_ram[1077] = 38;
    exp_48_ram[1078] = 133;
    exp_48_ram[1079] = 0;
    exp_48_ram[1080] = 39;
    exp_48_ram[1081] = 39;
    exp_48_ram[1082] = 7;
    exp_48_ram[1083] = 46;
    exp_48_ram[1084] = 35;
    exp_48_ram[1085] = 40;
    exp_48_ram[1086] = 40;
    exp_48_ram[1087] = 37;
    exp_48_ram[1088] = 37;
    exp_48_ram[1089] = 38;
    exp_48_ram[1090] = 38;
    exp_48_ram[1091] = 39;
    exp_48_ram[1092] = 39;
    exp_48_ram[1093] = 32;
    exp_48_ram[1094] = 34;
    exp_48_ram[1095] = 36;
    exp_48_ram[1096] = 38;
    exp_48_ram[1097] = 40;
    exp_48_ram[1098] = 42;
    exp_48_ram[1099] = 44;
    exp_48_ram[1100] = 46;
    exp_48_ram[1101] = 32;
    exp_48_ram[1102] = 7;
    exp_48_ram[1103] = 133;
    exp_48_ram[1104] = 0;
    exp_48_ram[1105] = 32;
    exp_48_ram[1106] = 34;
    exp_48_ram[1107] = 163;
    exp_48_ram[1108] = 168;
    exp_48_ram[1109] = 168;
    exp_48_ram[1110] = 165;
    exp_48_ram[1111] = 165;
    exp_48_ram[1112] = 166;
    exp_48_ram[1113] = 166;
    exp_48_ram[1114] = 167;
    exp_48_ram[1115] = 167;
    exp_48_ram[1116] = 32;
    exp_48_ram[1117] = 34;
    exp_48_ram[1118] = 36;
    exp_48_ram[1119] = 38;
    exp_48_ram[1120] = 40;
    exp_48_ram[1121] = 42;
    exp_48_ram[1122] = 44;
    exp_48_ram[1123] = 46;
    exp_48_ram[1124] = 32;
    exp_48_ram[1125] = 7;
    exp_48_ram[1126] = 133;
    exp_48_ram[1127] = 0;
    exp_48_ram[1128] = 44;
    exp_48_ram[1129] = 46;
    exp_48_ram[1130] = 39;
    exp_48_ram[1131] = 39;
    exp_48_ram[1132] = 228;
    exp_48_ram[1133] = 39;
    exp_48_ram[1134] = 39;
    exp_48_ram[1135] = 24;
    exp_48_ram[1136] = 39;
    exp_48_ram[1137] = 39;
    exp_48_ram[1138] = 232;
    exp_48_ram[1139] = 39;
    exp_48_ram[1140] = 39;
    exp_48_ram[1141] = 238;
    exp_48_ram[1142] = 39;
    exp_48_ram[1143] = 39;
    exp_48_ram[1144] = 28;
    exp_48_ram[1145] = 39;
    exp_48_ram[1146] = 39;
    exp_48_ram[1147] = 246;
    exp_48_ram[1148] = 7;
    exp_48_ram[1149] = 0;
    exp_48_ram[1150] = 7;
    exp_48_ram[1151] = 133;
    exp_48_ram[1152] = 32;
    exp_48_ram[1153] = 36;
    exp_48_ram[1154] = 36;
    exp_48_ram[1155] = 1;
    exp_48_ram[1156] = 128;
    exp_48_ram[1157] = 1;
    exp_48_ram[1158] = 46;
    exp_48_ram[1159] = 44;
    exp_48_ram[1160] = 4;
    exp_48_ram[1161] = 44;
    exp_48_ram[1162] = 46;
    exp_48_ram[1163] = 7;
    exp_48_ram[1164] = 37;
    exp_48_ram[1165] = 38;
    exp_48_ram[1166] = 133;
    exp_48_ram[1167] = 0;
    exp_48_ram[1168] = 35;
    exp_48_ram[1169] = 40;
    exp_48_ram[1170] = 40;
    exp_48_ram[1171] = 37;
    exp_48_ram[1172] = 37;
    exp_48_ram[1173] = 38;
    exp_48_ram[1174] = 38;
    exp_48_ram[1175] = 39;
    exp_48_ram[1176] = 39;
    exp_48_ram[1177] = 32;
    exp_48_ram[1178] = 34;
    exp_48_ram[1179] = 36;
    exp_48_ram[1180] = 38;
    exp_48_ram[1181] = 40;
    exp_48_ram[1182] = 42;
    exp_48_ram[1183] = 44;
    exp_48_ram[1184] = 46;
    exp_48_ram[1185] = 32;
    exp_48_ram[1186] = 7;
    exp_48_ram[1187] = 133;
    exp_48_ram[1188] = 240;
    exp_48_ram[1189] = 7;
    exp_48_ram[1190] = 133;
    exp_48_ram[1191] = 32;
    exp_48_ram[1192] = 36;
    exp_48_ram[1193] = 1;
    exp_48_ram[1194] = 128;
    exp_48_ram[1195] = 1;
    exp_48_ram[1196] = 46;
    exp_48_ram[1197] = 4;
    exp_48_ram[1198] = 6;
    exp_48_ram[1199] = 38;
    exp_48_ram[1200] = 6;
    exp_48_ram[1201] = 134;
    exp_48_ram[1202] = 36;
    exp_48_ram[1203] = 38;
    exp_48_ram[1204] = 166;
    exp_48_ram[1205] = 32;
    exp_48_ram[1206] = 34;
    exp_48_ram[1207] = 38;
    exp_48_ram[1208] = 150;
    exp_48_ram[1209] = 34;
    exp_48_ram[1210] = 32;
    exp_48_ram[1211] = 38;
    exp_48_ram[1212] = 166;
    exp_48_ram[1213] = 135;
    exp_48_ram[1214] = 7;
    exp_48_ram[1215] = 38;
    exp_48_ram[1216] = 230;
    exp_48_ram[1217] = 32;
    exp_48_ram[1218] = 38;
    exp_48_ram[1219] = 231;
    exp_48_ram[1220] = 34;
    exp_48_ram[1221] = 39;
    exp_48_ram[1222] = 39;
    exp_48_ram[1223] = 5;
    exp_48_ram[1224] = 133;
    exp_48_ram[1225] = 36;
    exp_48_ram[1226] = 1;
    exp_48_ram[1227] = 128;
    exp_48_ram[1228] = 1;
    exp_48_ram[1229] = 46;
    exp_48_ram[1230] = 44;
    exp_48_ram[1231] = 4;
    exp_48_ram[1232] = 36;
    exp_48_ram[1233] = 38;
    exp_48_ram[1234] = 32;
    exp_48_ram[1235] = 34;
    exp_48_ram[1236] = 39;
    exp_48_ram[1237] = 39;
    exp_48_ram[1238] = 37;
    exp_48_ram[1239] = 37;
    exp_48_ram[1240] = 6;
    exp_48_ram[1241] = 8;
    exp_48_ram[1242] = 56;
    exp_48_ram[1243] = 134;
    exp_48_ram[1244] = 135;
    exp_48_ram[1245] = 134;
    exp_48_ram[1246] = 7;
    exp_48_ram[1247] = 135;
    exp_48_ram[1248] = 5;
    exp_48_ram[1249] = 133;
    exp_48_ram[1250] = 240;
    exp_48_ram[1251] = 7;
    exp_48_ram[1252] = 135;
    exp_48_ram[1253] = 5;
    exp_48_ram[1254] = 133;
    exp_48_ram[1255] = 32;
    exp_48_ram[1256] = 36;
    exp_48_ram[1257] = 1;
    exp_48_ram[1258] = 128;
    exp_48_ram[1259] = 1;
    exp_48_ram[1260] = 46;
    exp_48_ram[1261] = 4;
    exp_48_ram[1262] = 38;
    exp_48_ram[1263] = 39;
    exp_48_ram[1264] = 247;
    exp_48_ram[1265] = 150;
    exp_48_ram[1266] = 39;
    exp_48_ram[1267] = 7;
    exp_48_ram[1268] = 119;
    exp_48_ram[1269] = 154;
    exp_48_ram[1270] = 39;
    exp_48_ram[1271] = 7;
    exp_48_ram[1272] = 119;
    exp_48_ram[1273] = 150;
    exp_48_ram[1274] = 7;
    exp_48_ram[1275] = 0;
    exp_48_ram[1276] = 7;
    exp_48_ram[1277] = 133;
    exp_48_ram[1278] = 36;
    exp_48_ram[1279] = 1;
    exp_48_ram[1280] = 128;
    exp_48_ram[1281] = 1;
    exp_48_ram[1282] = 46;
    exp_48_ram[1283] = 44;
    exp_48_ram[1284] = 4;
    exp_48_ram[1285] = 38;
    exp_48_ram[1286] = 37;
    exp_48_ram[1287] = 240;
    exp_48_ram[1288] = 7;
    exp_48_ram[1289] = 134;
    exp_48_ram[1290] = 7;
    exp_48_ram[1291] = 0;
    exp_48_ram[1292] = 7;
    exp_48_ram[1293] = 133;
    exp_48_ram[1294] = 32;
    exp_48_ram[1295] = 36;
    exp_48_ram[1296] = 1;
    exp_48_ram[1297] = 128;
    exp_48_ram[1298] = 1;
    exp_48_ram[1299] = 46;
    exp_48_ram[1300] = 44;
    exp_48_ram[1301] = 4;
    exp_48_ram[1302] = 38;
    exp_48_ram[1303] = 36;
    exp_48_ram[1304] = 39;
    exp_48_ram[1305] = 7;
    exp_48_ram[1306] = 4;
    exp_48_ram[1307] = 39;
    exp_48_ram[1308] = 7;
    exp_48_ram[1309] = 14;
    exp_48_ram[1310] = 39;
    exp_48_ram[1311] = 7;
    exp_48_ram[1312] = 8;
    exp_48_ram[1313] = 39;
    exp_48_ram[1314] = 7;
    exp_48_ram[1315] = 22;
    exp_48_ram[1316] = 7;
    exp_48_ram[1317] = 0;
    exp_48_ram[1318] = 39;
    exp_48_ram[1319] = 7;
    exp_48_ram[1320] = 18;
    exp_48_ram[1321] = 37;
    exp_48_ram[1322] = 240;
    exp_48_ram[1323] = 7;
    exp_48_ram[1324] = 134;
    exp_48_ram[1325] = 7;
    exp_48_ram[1326] = 0;
    exp_48_ram[1327] = 7;
    exp_48_ram[1328] = 0;
    exp_48_ram[1329] = 7;
    exp_48_ram[1330] = 133;
    exp_48_ram[1331] = 32;
    exp_48_ram[1332] = 36;
    exp_48_ram[1333] = 1;
    exp_48_ram[1334] = 128;
    exp_48_ram[1335] = 1;
    exp_48_ram[1336] = 38;
    exp_48_ram[1337] = 36;
    exp_48_ram[1338] = 34;
    exp_48_ram[1339] = 32;
    exp_48_ram[1340] = 46;
    exp_48_ram[1341] = 44;
    exp_48_ram[1342] = 42;
    exp_48_ram[1343] = 40;
    exp_48_ram[1344] = 38;
    exp_48_ram[1345] = 36;
    exp_48_ram[1346] = 34;
    exp_48_ram[1347] = 32;
    exp_48_ram[1348] = 46;
    exp_48_ram[1349] = 4;
    exp_48_ram[1350] = 4;
    exp_48_ram[1351] = 7;
    exp_48_ram[1352] = 8;
    exp_48_ram[1353] = 44;
    exp_48_ram[1354] = 46;
    exp_48_ram[1355] = 7;
    exp_48_ram[1356] = 42;
    exp_48_ram[1357] = 167;
    exp_48_ram[1358] = 38;
    exp_48_ram[1359] = 39;
    exp_48_ram[1360] = 135;
    exp_48_ram[1361] = 39;
    exp_48_ram[1362] = 6;
    exp_48_ram[1363] = 37;
    exp_48_ram[1364] = 240;
    exp_48_ram[1365] = 7;
    exp_48_ram[1366] = 87;
    exp_48_ram[1367] = 135;
    exp_48_ram[1368] = 7;
    exp_48_ram[1369] = 44;
    exp_48_ram[1370] = 46;
    exp_48_ram[1371] = 38;
    exp_48_ram[1372] = 38;
    exp_48_ram[1373] = 40;
    exp_48_ram[1374] = 40;
    exp_48_ram[1375] = 5;
    exp_48_ram[1376] = 7;
    exp_48_ram[1377] = 5;
    exp_48_ram[1378] = 181;
    exp_48_ram[1379] = 133;
    exp_48_ram[1380] = 135;
    exp_48_ram[1381] = 134;
    exp_48_ram[1382] = 135;
    exp_48_ram[1383] = 44;
    exp_48_ram[1384] = 46;
    exp_48_ram[1385] = 39;
    exp_48_ram[1386] = 135;
    exp_48_ram[1387] = 42;
    exp_48_ram[1388] = 240;
    exp_48_ram[1389] = 0;
    exp_48_ram[1390] = 40;
    exp_48_ram[1391] = 167;
    exp_48_ram[1392] = 135;
    exp_48_ram[1393] = 39;
    exp_48_ram[1394] = 128;
    exp_48_ram[1395] = 37;
    exp_48_ram[1396] = 37;
    exp_48_ram[1397] = 240;
    exp_48_ram[1398] = 7;
    exp_48_ram[1399] = 87;
    exp_48_ram[1400] = 135;
    exp_48_ram[1401] = 7;
    exp_48_ram[1402] = 141;
    exp_48_ram[1403] = 13;
    exp_48_ram[1404] = 38;
    exp_48_ram[1405] = 38;
    exp_48_ram[1406] = 7;
    exp_48_ram[1407] = 5;
    exp_48_ram[1408] = 181;
    exp_48_ram[1409] = 135;
    exp_48_ram[1410] = 134;
    exp_48_ram[1411] = 135;
    exp_48_ram[1412] = 44;
    exp_48_ram[1413] = 46;
    exp_48_ram[1414] = 39;
    exp_48_ram[1415] = 135;
    exp_48_ram[1416] = 40;
    exp_48_ram[1417] = 240;
    exp_48_ram[1418] = 0;
    exp_48_ram[1419] = 167;
    exp_48_ram[1420] = 135;
    exp_48_ram[1421] = 87;
    exp_48_ram[1422] = 135;
    exp_48_ram[1423] = 7;
    exp_48_ram[1424] = 140;
    exp_48_ram[1425] = 215;
    exp_48_ram[1426] = 140;
    exp_48_ram[1427] = 38;
    exp_48_ram[1428] = 38;
    exp_48_ram[1429] = 7;
    exp_48_ram[1430] = 5;
    exp_48_ram[1431] = 181;
    exp_48_ram[1432] = 135;
    exp_48_ram[1433] = 134;
    exp_48_ram[1434] = 135;
    exp_48_ram[1435] = 44;
    exp_48_ram[1436] = 46;
    exp_48_ram[1437] = 167;
    exp_48_ram[1438] = 23;
    exp_48_ram[1439] = 135;
    exp_48_ram[1440] = 7;
    exp_48_ram[1441] = 139;
    exp_48_ram[1442] = 215;
    exp_48_ram[1443] = 139;
    exp_48_ram[1444] = 38;
    exp_48_ram[1445] = 38;
    exp_48_ram[1446] = 7;
    exp_48_ram[1447] = 5;
    exp_48_ram[1448] = 181;
    exp_48_ram[1449] = 135;
    exp_48_ram[1450] = 134;
    exp_48_ram[1451] = 135;
    exp_48_ram[1452] = 44;
    exp_48_ram[1453] = 46;
    exp_48_ram[1454] = 167;
    exp_48_ram[1455] = 7;
    exp_48_ram[1456] = 151;
    exp_48_ram[1457] = 135;
    exp_48_ram[1458] = 151;
    exp_48_ram[1459] = 138;
    exp_48_ram[1460] = 215;
    exp_48_ram[1461] = 138;
    exp_48_ram[1462] = 38;
    exp_48_ram[1463] = 38;
    exp_48_ram[1464] = 7;
    exp_48_ram[1465] = 5;
    exp_48_ram[1466] = 181;
    exp_48_ram[1467] = 135;
    exp_48_ram[1468] = 134;
    exp_48_ram[1469] = 135;
    exp_48_ram[1470] = 44;
    exp_48_ram[1471] = 46;
    exp_48_ram[1472] = 167;
    exp_48_ram[1473] = 137;
    exp_48_ram[1474] = 215;
    exp_48_ram[1475] = 137;
    exp_48_ram[1476] = 38;
    exp_48_ram[1477] = 38;
    exp_48_ram[1478] = 7;
    exp_48_ram[1479] = 5;
    exp_48_ram[1480] = 181;
    exp_48_ram[1481] = 135;
    exp_48_ram[1482] = 134;
    exp_48_ram[1483] = 135;
    exp_48_ram[1484] = 44;
    exp_48_ram[1485] = 46;
    exp_48_ram[1486] = 39;
    exp_48_ram[1487] = 39;
    exp_48_ram[1488] = 5;
    exp_48_ram[1489] = 133;
    exp_48_ram[1490] = 32;
    exp_48_ram[1491] = 36;
    exp_48_ram[1492] = 36;
    exp_48_ram[1493] = 41;
    exp_48_ram[1494] = 41;
    exp_48_ram[1495] = 42;
    exp_48_ram[1496] = 42;
    exp_48_ram[1497] = 43;
    exp_48_ram[1498] = 43;
    exp_48_ram[1499] = 44;
    exp_48_ram[1500] = 44;
    exp_48_ram[1501] = 45;
    exp_48_ram[1502] = 45;
    exp_48_ram[1503] = 1;
    exp_48_ram[1504] = 128;
    exp_48_ram[1505] = 1;
    exp_48_ram[1506] = 46;
    exp_48_ram[1507] = 44;
    exp_48_ram[1508] = 42;
    exp_48_ram[1509] = 40;
    exp_48_ram[1510] = 38;
    exp_48_ram[1511] = 4;
    exp_48_ram[1512] = 46;
    exp_48_ram[1513] = 39;
    exp_48_ram[1514] = 163;
    exp_48_ram[1515] = 168;
    exp_48_ram[1516] = 168;
    exp_48_ram[1517] = 165;
    exp_48_ram[1518] = 165;
    exp_48_ram[1519] = 166;
    exp_48_ram[1520] = 166;
    exp_48_ram[1521] = 167;
    exp_48_ram[1522] = 167;
    exp_48_ram[1523] = 38;
    exp_48_ram[1524] = 40;
    exp_48_ram[1525] = 42;
    exp_48_ram[1526] = 44;
    exp_48_ram[1527] = 46;
    exp_48_ram[1528] = 32;
    exp_48_ram[1529] = 34;
    exp_48_ram[1530] = 36;
    exp_48_ram[1531] = 38;
    exp_48_ram[1532] = 35;
    exp_48_ram[1533] = 40;
    exp_48_ram[1534] = 40;
    exp_48_ram[1535] = 37;
    exp_48_ram[1536] = 37;
    exp_48_ram[1537] = 38;
    exp_48_ram[1538] = 38;
    exp_48_ram[1539] = 39;
    exp_48_ram[1540] = 39;
    exp_48_ram[1541] = 32;
    exp_48_ram[1542] = 34;
    exp_48_ram[1543] = 36;
    exp_48_ram[1544] = 38;
    exp_48_ram[1545] = 40;
    exp_48_ram[1546] = 42;
    exp_48_ram[1547] = 44;
    exp_48_ram[1548] = 46;
    exp_48_ram[1549] = 32;
    exp_48_ram[1550] = 7;
    exp_48_ram[1551] = 133;
    exp_48_ram[1552] = 240;
    exp_48_ram[1553] = 40;
    exp_48_ram[1554] = 42;
    exp_48_ram[1555] = 39;
    exp_48_ram[1556] = 94;
    exp_48_ram[1557] = 38;
    exp_48_ram[1558] = 38;
    exp_48_ram[1559] = 245;
    exp_48_ram[1560] = 5;
    exp_48_ram[1561] = 5;
    exp_48_ram[1562] = 7;
    exp_48_ram[1563] = 8;
    exp_48_ram[1564] = 56;
    exp_48_ram[1565] = 135;
    exp_48_ram[1566] = 6;
    exp_48_ram[1567] = 135;
    exp_48_ram[1568] = 44;
    exp_48_ram[1569] = 46;
    exp_48_ram[1570] = 0;
    exp_48_ram[1571] = 39;
    exp_48_ram[1572] = 210;
    exp_48_ram[1573] = 35;
    exp_48_ram[1574] = 40;
    exp_48_ram[1575] = 40;
    exp_48_ram[1576] = 37;
    exp_48_ram[1577] = 37;
    exp_48_ram[1578] = 38;
    exp_48_ram[1579] = 38;
    exp_48_ram[1580] = 39;
    exp_48_ram[1581] = 39;
    exp_48_ram[1582] = 32;
    exp_48_ram[1583] = 34;
    exp_48_ram[1584] = 36;
    exp_48_ram[1585] = 38;
    exp_48_ram[1586] = 40;
    exp_48_ram[1587] = 42;
    exp_48_ram[1588] = 44;
    exp_48_ram[1589] = 46;
    exp_48_ram[1590] = 32;
    exp_48_ram[1591] = 7;
    exp_48_ram[1592] = 133;
    exp_48_ram[1593] = 240;
    exp_48_ram[1594] = 7;
    exp_48_ram[1595] = 138;
    exp_48_ram[1596] = 22;
    exp_48_ram[1597] = 6;
    exp_48_ram[1598] = 6;
    exp_48_ram[1599] = 0;
    exp_48_ram[1600] = 6;
    exp_48_ram[1601] = 6;
    exp_48_ram[1602] = 37;
    exp_48_ram[1603] = 37;
    exp_48_ram[1604] = 7;
    exp_48_ram[1605] = 8;
    exp_48_ram[1606] = 56;
    exp_48_ram[1607] = 135;
    exp_48_ram[1608] = 134;
    exp_48_ram[1609] = 135;
    exp_48_ram[1610] = 44;
    exp_48_ram[1611] = 46;
    exp_48_ram[1612] = 0;
    exp_48_ram[1613] = 39;
    exp_48_ram[1614] = 39;
    exp_48_ram[1615] = 44;
    exp_48_ram[1616] = 46;
    exp_48_ram[1617] = 71;
    exp_48_ram[1618] = 167;
    exp_48_ram[1619] = 137;
    exp_48_ram[1620] = 215;
    exp_48_ram[1621] = 137;
    exp_48_ram[1622] = 38;
    exp_48_ram[1623] = 38;
    exp_48_ram[1624] = 7;
    exp_48_ram[1625] = 5;
    exp_48_ram[1626] = 53;
    exp_48_ram[1627] = 135;
    exp_48_ram[1628] = 134;
    exp_48_ram[1629] = 135;
    exp_48_ram[1630] = 44;
    exp_48_ram[1631] = 46;
    exp_48_ram[1632] = 36;
    exp_48_ram[1633] = 7;
    exp_48_ram[1634] = 37;
    exp_48_ram[1635] = 38;
    exp_48_ram[1636] = 133;
    exp_48_ram[1637] = 0;
    exp_48_ram[1638] = 35;
    exp_48_ram[1639] = 40;
    exp_48_ram[1640] = 40;
    exp_48_ram[1641] = 37;
    exp_48_ram[1642] = 37;
    exp_48_ram[1643] = 38;
    exp_48_ram[1644] = 38;
    exp_48_ram[1645] = 39;
    exp_48_ram[1646] = 39;
    exp_48_ram[1647] = 160;
    exp_48_ram[1648] = 162;
    exp_48_ram[1649] = 164;
    exp_48_ram[1650] = 166;
    exp_48_ram[1651] = 168;
    exp_48_ram[1652] = 170;
    exp_48_ram[1653] = 172;
    exp_48_ram[1654] = 174;
    exp_48_ram[1655] = 160;
    exp_48_ram[1656] = 39;
    exp_48_ram[1657] = 90;
    exp_48_ram[1658] = 39;
    exp_48_ram[1659] = 7;
    exp_48_ram[1660] = 160;
    exp_48_ram[1661] = 0;
    exp_48_ram[1662] = 39;
    exp_48_ram[1663] = 212;
    exp_48_ram[1664] = 35;
    exp_48_ram[1665] = 40;
    exp_48_ram[1666] = 40;
    exp_48_ram[1667] = 37;
    exp_48_ram[1668] = 37;
    exp_48_ram[1669] = 38;
    exp_48_ram[1670] = 38;
    exp_48_ram[1671] = 39;
    exp_48_ram[1672] = 39;
    exp_48_ram[1673] = 32;
    exp_48_ram[1674] = 34;
    exp_48_ram[1675] = 36;
    exp_48_ram[1676] = 38;
    exp_48_ram[1677] = 40;
    exp_48_ram[1678] = 42;
    exp_48_ram[1679] = 44;
    exp_48_ram[1680] = 46;
    exp_48_ram[1681] = 32;
    exp_48_ram[1682] = 7;
    exp_48_ram[1683] = 133;
    exp_48_ram[1684] = 240;
    exp_48_ram[1685] = 7;
    exp_48_ram[1686] = 39;
    exp_48_ram[1687] = 160;
    exp_48_ram[1688] = 0;
    exp_48_ram[1689] = 39;
    exp_48_ram[1690] = 160;
    exp_48_ram[1691] = 39;
    exp_48_ram[1692] = 39;
    exp_48_ram[1693] = 5;
    exp_48_ram[1694] = 133;
    exp_48_ram[1695] = 32;
    exp_48_ram[1696] = 36;
    exp_48_ram[1697] = 36;
    exp_48_ram[1698] = 41;
    exp_48_ram[1699] = 41;
    exp_48_ram[1700] = 1;
    exp_48_ram[1701] = 128;
    exp_48_ram[1702] = 1;
    exp_48_ram[1703] = 46;
    exp_48_ram[1704] = 44;
    exp_48_ram[1705] = 42;
    exp_48_ram[1706] = 40;
    exp_48_ram[1707] = 38;
    exp_48_ram[1708] = 36;
    exp_48_ram[1709] = 34;
    exp_48_ram[1710] = 32;
    exp_48_ram[1711] = 4;
    exp_48_ram[1712] = 38;
    exp_48_ram[1713] = 240;
    exp_48_ram[1714] = 7;
    exp_48_ram[1715] = 135;
    exp_48_ram[1716] = 70;
    exp_48_ram[1717] = 166;
    exp_48_ram[1718] = 138;
    exp_48_ram[1719] = 10;
    exp_48_ram[1720] = 6;
    exp_48_ram[1721] = 134;
    exp_48_ram[1722] = 5;
    exp_48_ram[1723] = 133;
    exp_48_ram[1724] = 224;
    exp_48_ram[1725] = 7;
    exp_48_ram[1726] = 135;
    exp_48_ram[1727] = 46;
    exp_48_ram[1728] = 71;
    exp_48_ram[1729] = 167;
    exp_48_ram[1730] = 167;
    exp_48_ram[1731] = 39;
    exp_48_ram[1732] = 135;
    exp_48_ram[1733] = 46;
    exp_48_ram[1734] = 39;
    exp_48_ram[1735] = 142;
    exp_48_ram[1736] = 39;
    exp_48_ram[1737] = 137;
    exp_48_ram[1738] = 9;
    exp_48_ram[1739] = 39;
    exp_48_ram[1740] = 160;
    exp_48_ram[1741] = 162;
    exp_48_ram[1742] = 39;
    exp_48_ram[1743] = 139;
    exp_48_ram[1744] = 11;
    exp_48_ram[1745] = 7;
    exp_48_ram[1746] = 135;
    exp_48_ram[1747] = 5;
    exp_48_ram[1748] = 133;
    exp_48_ram[1749] = 32;
    exp_48_ram[1750] = 36;
    exp_48_ram[1751] = 41;
    exp_48_ram[1752] = 41;
    exp_48_ram[1753] = 42;
    exp_48_ram[1754] = 42;
    exp_48_ram[1755] = 43;
    exp_48_ram[1756] = 43;
    exp_48_ram[1757] = 1;
    exp_48_ram[1758] = 128;
    exp_48_ram[1759] = 1;
    exp_48_ram[1760] = 38;
    exp_48_ram[1761] = 36;
    exp_48_ram[1762] = 34;
    exp_48_ram[1763] = 32;
    exp_48_ram[1764] = 4;
    exp_48_ram[1765] = 44;
    exp_48_ram[1766] = 46;
    exp_48_ram[1767] = 240;
    exp_48_ram[1768] = 7;
    exp_48_ram[1769] = 135;
    exp_48_ram[1770] = 70;
    exp_48_ram[1771] = 166;
    exp_48_ram[1772] = 137;
    exp_48_ram[1773] = 9;
    exp_48_ram[1774] = 6;
    exp_48_ram[1775] = 134;
    exp_48_ram[1776] = 5;
    exp_48_ram[1777] = 133;
    exp_48_ram[1778] = 224;
    exp_48_ram[1779] = 7;
    exp_48_ram[1780] = 135;
    exp_48_ram[1781] = 36;
    exp_48_ram[1782] = 38;
    exp_48_ram[1783] = 39;
    exp_48_ram[1784] = 39;
    exp_48_ram[1785] = 37;
    exp_48_ram[1786] = 37;
    exp_48_ram[1787] = 6;
    exp_48_ram[1788] = 8;
    exp_48_ram[1789] = 56;
    exp_48_ram[1790] = 134;
    exp_48_ram[1791] = 135;
    exp_48_ram[1792] = 134;
    exp_48_ram[1793] = 7;
    exp_48_ram[1794] = 135;
    exp_48_ram[1795] = 70;
    exp_48_ram[1796] = 164;
    exp_48_ram[1797] = 166;
    exp_48_ram[1798] = 0;
    exp_48_ram[1799] = 32;
    exp_48_ram[1800] = 36;
    exp_48_ram[1801] = 41;
    exp_48_ram[1802] = 41;
    exp_48_ram[1803] = 1;
    exp_48_ram[1804] = 128;
    exp_48_ram[1805] = 1;
    exp_48_ram[1806] = 38;
    exp_48_ram[1807] = 36;
    exp_48_ram[1808] = 4;
    exp_48_ram[1809] = 46;
    exp_48_ram[1810] = 23;
    exp_48_ram[1811] = 135;
    exp_48_ram[1812] = 165;
    exp_48_ram[1813] = 165;
    exp_48_ram[1814] = 166;
    exp_48_ram[1815] = 166;
    exp_48_ram[1816] = 167;
    exp_48_ram[1817] = 42;
    exp_48_ram[1818] = 44;
    exp_48_ram[1819] = 46;
    exp_48_ram[1820] = 32;
    exp_48_ram[1821] = 34;
    exp_48_ram[1822] = 215;
    exp_48_ram[1823] = 20;
    exp_48_ram[1824] = 23;
    exp_48_ram[1825] = 135;
    exp_48_ram[1826] = 174;
    exp_48_ram[1827] = 163;
    exp_48_ram[1828] = 168;
    exp_48_ram[1829] = 168;
    exp_48_ram[1830] = 165;
    exp_48_ram[1831] = 165;
    exp_48_ram[1832] = 166;
    exp_48_ram[1833] = 166;
    exp_48_ram[1834] = 167;
    exp_48_ram[1835] = 38;
    exp_48_ram[1836] = 40;
    exp_48_ram[1837] = 42;
    exp_48_ram[1838] = 44;
    exp_48_ram[1839] = 46;
    exp_48_ram[1840] = 32;
    exp_48_ram[1841] = 34;
    exp_48_ram[1842] = 36;
    exp_48_ram[1843] = 38;
    exp_48_ram[1844] = 199;
    exp_48_ram[1845] = 8;
    exp_48_ram[1846] = 38;
    exp_48_ram[1847] = 0;
    exp_48_ram[1848] = 39;
    exp_48_ram[1849] = 167;
    exp_48_ram[1850] = 7;
    exp_48_ram[1851] = 151;
    exp_48_ram[1852] = 135;
    exp_48_ram[1853] = 39;
    exp_48_ram[1854] = 7;
    exp_48_ram[1855] = 7;
    exp_48_ram[1856] = 7;
    exp_48_ram[1857] = 199;
    exp_48_ram[1858] = 71;
    exp_48_ram[1859] = 134;
    exp_48_ram[1860] = 39;
    exp_48_ram[1861] = 135;
    exp_48_ram[1862] = 128;
    exp_48_ram[1863] = 39;
    exp_48_ram[1864] = 135;
    exp_48_ram[1865] = 38;
    exp_48_ram[1866] = 39;
    exp_48_ram[1867] = 7;
    exp_48_ram[1868] = 216;
    exp_48_ram[1869] = 71;
    exp_48_ram[1870] = 135;
    exp_48_ram[1871] = 7;
    exp_48_ram[1872] = 129;
    exp_48_ram[1873] = 38;
    exp_48_ram[1874] = 0;
    exp_48_ram[1875] = 39;
    exp_48_ram[1876] = 167;
    exp_48_ram[1877] = 7;
    exp_48_ram[1878] = 151;
    exp_48_ram[1879] = 135;
    exp_48_ram[1880] = 39;
    exp_48_ram[1881] = 7;
    exp_48_ram[1882] = 39;
    exp_48_ram[1883] = 135;
    exp_48_ram[1884] = 6;
    exp_48_ram[1885] = 135;
    exp_48_ram[1886] = 71;
    exp_48_ram[1887] = 70;
    exp_48_ram[1888] = 134;
    exp_48_ram[1889] = 135;
    exp_48_ram[1890] = 128;
    exp_48_ram[1891] = 39;
    exp_48_ram[1892] = 135;
    exp_48_ram[1893] = 38;
    exp_48_ram[1894] = 39;
    exp_48_ram[1895] = 7;
    exp_48_ram[1896] = 214;
    exp_48_ram[1897] = 71;
    exp_48_ram[1898] = 135;
    exp_48_ram[1899] = 7;
    exp_48_ram[1900] = 131;
    exp_48_ram[1901] = 39;
    exp_48_ram[1902] = 167;
    exp_48_ram[1903] = 5;
    exp_48_ram[1904] = 133;
    exp_48_ram[1905] = 32;
    exp_48_ram[1906] = 7;
    exp_48_ram[1907] = 135;
    exp_48_ram[1908] = 34;
    exp_48_ram[1909] = 36;
    exp_48_ram[1910] = 39;
    exp_48_ram[1911] = 247;
    exp_48_ram[1912] = 135;
    exp_48_ram[1913] = 247;
    exp_48_ram[1914] = 71;
    exp_48_ram[1915] = 135;
    exp_48_ram[1916] = 132;
    exp_48_ram[1917] = 39;
    exp_48_ram[1918] = 247;
    exp_48_ram[1919] = 135;
    exp_48_ram[1920] = 247;
    exp_48_ram[1921] = 71;
    exp_48_ram[1922] = 135;
    exp_48_ram[1923] = 132;
    exp_48_ram[1924] = 71;
    exp_48_ram[1925] = 135;
    exp_48_ram[1926] = 7;
    exp_48_ram[1927] = 133;
    exp_48_ram[1928] = 39;
    exp_48_ram[1929] = 167;
    exp_48_ram[1930] = 5;
    exp_48_ram[1931] = 133;
    exp_48_ram[1932] = 32;
    exp_48_ram[1933] = 7;
    exp_48_ram[1934] = 135;
    exp_48_ram[1935] = 34;
    exp_48_ram[1936] = 36;
    exp_48_ram[1937] = 39;
    exp_48_ram[1938] = 247;
    exp_48_ram[1939] = 135;
    exp_48_ram[1940] = 247;
    exp_48_ram[1941] = 71;
    exp_48_ram[1942] = 135;
    exp_48_ram[1943] = 133;
    exp_48_ram[1944] = 39;
    exp_48_ram[1945] = 247;
    exp_48_ram[1946] = 135;
    exp_48_ram[1947] = 247;
    exp_48_ram[1948] = 71;
    exp_48_ram[1949] = 135;
    exp_48_ram[1950] = 134;
    exp_48_ram[1951] = 71;
    exp_48_ram[1952] = 135;
    exp_48_ram[1953] = 7;
    exp_48_ram[1954] = 134;
    exp_48_ram[1955] = 39;
    exp_48_ram[1956] = 167;
    exp_48_ram[1957] = 5;
    exp_48_ram[1958] = 133;
    exp_48_ram[1959] = 32;
    exp_48_ram[1960] = 7;
    exp_48_ram[1961] = 135;
    exp_48_ram[1962] = 34;
    exp_48_ram[1963] = 36;
    exp_48_ram[1964] = 39;
    exp_48_ram[1965] = 247;
    exp_48_ram[1966] = 135;
    exp_48_ram[1967] = 247;
    exp_48_ram[1968] = 71;
    exp_48_ram[1969] = 135;
    exp_48_ram[1970] = 135;
    exp_48_ram[1971] = 39;
    exp_48_ram[1972] = 247;
    exp_48_ram[1973] = 135;
    exp_48_ram[1974] = 247;
    exp_48_ram[1975] = 71;
    exp_48_ram[1976] = 135;
    exp_48_ram[1977] = 135;
    exp_48_ram[1978] = 71;
    exp_48_ram[1979] = 135;
    exp_48_ram[1980] = 7;
    exp_48_ram[1981] = 136;
    exp_48_ram[1982] = 39;
    exp_48_ram[1983] = 167;
    exp_48_ram[1984] = 5;
    exp_48_ram[1985] = 133;
    exp_48_ram[1986] = 16;
    exp_48_ram[1987] = 7;
    exp_48_ram[1988] = 135;
    exp_48_ram[1989] = 34;
    exp_48_ram[1990] = 36;
    exp_48_ram[1991] = 39;
    exp_48_ram[1992] = 247;
    exp_48_ram[1993] = 135;
    exp_48_ram[1994] = 247;
    exp_48_ram[1995] = 71;
    exp_48_ram[1996] = 135;
    exp_48_ram[1997] = 136;
    exp_48_ram[1998] = 39;
    exp_48_ram[1999] = 247;
    exp_48_ram[2000] = 135;
    exp_48_ram[2001] = 247;
    exp_48_ram[2002] = 71;
    exp_48_ram[2003] = 135;
    exp_48_ram[2004] = 137;
    exp_48_ram[2005] = 71;
    exp_48_ram[2006] = 135;
    exp_48_ram[2007] = 7;
    exp_48_ram[2008] = 137;
    exp_48_ram[2009] = 39;
    exp_48_ram[2010] = 167;
    exp_48_ram[2011] = 135;
    exp_48_ram[2012] = 5;
    exp_48_ram[2013] = 133;
    exp_48_ram[2014] = 16;
    exp_48_ram[2015] = 7;
    exp_48_ram[2016] = 135;
    exp_48_ram[2017] = 34;
    exp_48_ram[2018] = 36;
    exp_48_ram[2019] = 39;
    exp_48_ram[2020] = 247;
    exp_48_ram[2021] = 135;
    exp_48_ram[2022] = 247;
    exp_48_ram[2023] = 71;
    exp_48_ram[2024] = 135;
    exp_48_ram[2025] = 138;
    exp_48_ram[2026] = 39;
    exp_48_ram[2027] = 5;
    exp_48_ram[2028] = 133;
    exp_48_ram[2029] = 16;
    exp_48_ram[2030] = 7;
    exp_48_ram[2031] = 135;
    exp_48_ram[2032] = 34;
    exp_48_ram[2033] = 36;
    exp_48_ram[2034] = 39;
    exp_48_ram[2035] = 247;
    exp_48_ram[2036] = 135;
    exp_48_ram[2037] = 247;
    exp_48_ram[2038] = 71;
    exp_48_ram[2039] = 135;
    exp_48_ram[2040] = 138;
    exp_48_ram[2041] = 39;
    exp_48_ram[2042] = 5;
    exp_48_ram[2043] = 133;
    exp_48_ram[2044] = 16;
    exp_48_ram[2045] = 7;
    exp_48_ram[2046] = 135;
    exp_48_ram[2047] = 34;
    exp_48_ram[2048] = 36;
    exp_48_ram[2049] = 39;
    exp_48_ram[2050] = 247;
    exp_48_ram[2051] = 135;
    exp_48_ram[2052] = 247;
    exp_48_ram[2053] = 71;
    exp_48_ram[2054] = 135;
    exp_48_ram[2055] = 139;
    exp_48_ram[2056] = 39;
    exp_48_ram[2057] = 247;
    exp_48_ram[2058] = 135;
    exp_48_ram[2059] = 247;
    exp_48_ram[2060] = 71;
    exp_48_ram[2061] = 135;
    exp_48_ram[2062] = 139;
    exp_48_ram[2063] = 71;
    exp_48_ram[2064] = 135;
    exp_48_ram[2065] = 7;
    exp_48_ram[2066] = 140;
    exp_48_ram[2067] = 71;
    exp_48_ram[2068] = 135;
    exp_48_ram[2069] = 140;
    exp_48_ram[2070] = 71;
    exp_48_ram[2071] = 135;
    exp_48_ram[2072] = 133;
    exp_48_ram[2073] = 32;
    exp_48_ram[2074] = 36;
    exp_48_ram[2075] = 1;
    exp_48_ram[2076] = 128;
    exp_48_ram[2077] = 1;
    exp_48_ram[2078] = 46;
    exp_48_ram[2079] = 44;
    exp_48_ram[2080] = 4;
    exp_48_ram[2081] = 38;
    exp_48_ram[2082] = 37;
    exp_48_ram[2083] = 0;
    exp_48_ram[2084] = 7;
    exp_48_ram[2085] = 133;
    exp_48_ram[2086] = 240;
    exp_48_ram[2087] = 7;
    exp_48_ram[2088] = 133;
    exp_48_ram[2089] = 32;
    exp_48_ram[2090] = 36;
    exp_48_ram[2091] = 1;
    exp_48_ram[2092] = 128;
    exp_48_ram[2093] = 1;
    exp_48_ram[2094] = 46;
    exp_48_ram[2095] = 44;
    exp_48_ram[2096] = 42;
    exp_48_ram[2097] = 40;
    exp_48_ram[2098] = 38;
    exp_48_ram[2099] = 36;
    exp_48_ram[2100] = 34;
    exp_48_ram[2101] = 32;
    exp_48_ram[2102] = 46;
    exp_48_ram[2103] = 44;
    exp_48_ram[2104] = 4;
    exp_48_ram[2105] = 38;
    exp_48_ram[2106] = 32;
    exp_48_ram[2107] = 34;
    exp_48_ram[2108] = 7;
    exp_48_ram[2109] = 44;
    exp_48_ram[2110] = 7;
    exp_48_ram[2111] = 46;
    exp_48_ram[2112] = 39;
    exp_48_ram[2113] = 133;
    exp_48_ram[2114] = 240;
    exp_48_ram[2115] = 38;
    exp_48_ram[2116] = 39;
    exp_48_ram[2117] = 87;
    exp_48_ram[2118] = 135;
    exp_48_ram[2119] = 7;
    exp_48_ram[2120] = 36;
    exp_48_ram[2121] = 39;
    exp_48_ram[2122] = 140;
    exp_48_ram[2123] = 12;
    exp_48_ram[2124] = 39;
    exp_48_ram[2125] = 135;
    exp_48_ram[2126] = 234;
    exp_48_ram[2127] = 39;
    exp_48_ram[2128] = 135;
    exp_48_ram[2129] = 152;
    exp_48_ram[2130] = 39;
    exp_48_ram[2131] = 7;
    exp_48_ram[2132] = 238;
    exp_48_ram[2133] = 39;
    exp_48_ram[2134] = 135;
    exp_48_ram[2135] = 44;
    exp_48_ram[2136] = 39;
    exp_48_ram[2137] = 135;
    exp_48_ram[2138] = 39;
    exp_48_ram[2139] = 7;
    exp_48_ram[2140] = 46;
    exp_48_ram[2141] = 39;
    exp_48_ram[2142] = 138;
    exp_48_ram[2143] = 10;
    exp_48_ram[2144] = 38;
    exp_48_ram[2145] = 38;
    exp_48_ram[2146] = 7;
    exp_48_ram[2147] = 5;
    exp_48_ram[2148] = 53;
    exp_48_ram[2149] = 135;
    exp_48_ram[2150] = 134;
    exp_48_ram[2151] = 135;
    exp_48_ram[2152] = 32;
    exp_48_ram[2153] = 34;
    exp_48_ram[2154] = 240;
    exp_48_ram[2155] = 0;
    exp_48_ram[2156] = 42;
    exp_48_ram[2157] = 32;
    exp_48_ram[2158] = 39;
    exp_48_ram[2159] = 135;
    exp_48_ram[2160] = 39;
    exp_48_ram[2161] = 133;
    exp_48_ram[2162] = 5;
    exp_48_ram[2163] = 240;
    exp_48_ram[2164] = 38;
    exp_48_ram[2165] = 39;
    exp_48_ram[2166] = 87;
    exp_48_ram[2167] = 135;
    exp_48_ram[2168] = 7;
    exp_48_ram[2169] = 36;
    exp_48_ram[2170] = 39;
    exp_48_ram[2171] = 139;
    exp_48_ram[2172] = 11;
    exp_48_ram[2173] = 39;
    exp_48_ram[2174] = 135;
    exp_48_ram[2175] = 228;
    exp_48_ram[2176] = 39;
    exp_48_ram[2177] = 135;
    exp_48_ram[2178] = 152;
    exp_48_ram[2179] = 39;
    exp_48_ram[2180] = 7;
    exp_48_ram[2181] = 232;
    exp_48_ram[2182] = 39;
    exp_48_ram[2183] = 135;
    exp_48_ram[2184] = 42;
    exp_48_ram[2185] = 39;
    exp_48_ram[2186] = 135;
    exp_48_ram[2187] = 39;
    exp_48_ram[2188] = 7;
    exp_48_ram[2189] = 46;
    exp_48_ram[2190] = 39;
    exp_48_ram[2191] = 135;
    exp_48_ram[2192] = 39;
    exp_48_ram[2193] = 7;
    exp_48_ram[2194] = 32;
    exp_48_ram[2195] = 39;
    exp_48_ram[2196] = 137;
    exp_48_ram[2197] = 9;
    exp_48_ram[2198] = 38;
    exp_48_ram[2199] = 38;
    exp_48_ram[2200] = 7;
    exp_48_ram[2201] = 5;
    exp_48_ram[2202] = 53;
    exp_48_ram[2203] = 135;
    exp_48_ram[2204] = 134;
    exp_48_ram[2205] = 135;
    exp_48_ram[2206] = 32;
    exp_48_ram[2207] = 34;
    exp_48_ram[2208] = 240;
    exp_48_ram[2209] = 0;
    exp_48_ram[2210] = 39;
    exp_48_ram[2211] = 135;
    exp_48_ram[2212] = 44;
    exp_48_ram[2213] = 39;
    exp_48_ram[2214] = 87;
    exp_48_ram[2215] = 133;
    exp_48_ram[2216] = 5;
    exp_48_ram[2217] = 16;
    exp_48_ram[2218] = 7;
    exp_48_ram[2219] = 135;
    exp_48_ram[2220] = 46;
    exp_48_ram[2221] = 32;
    exp_48_ram[2222] = 39;
    exp_48_ram[2223] = 135;
    exp_48_ram[2224] = 40;
    exp_48_ram[2225] = 39;
    exp_48_ram[2226] = 39;
    exp_48_ram[2227] = 7;
    exp_48_ram[2228] = 46;
    exp_48_ram[2229] = 39;
    exp_48_ram[2230] = 7;
    exp_48_ram[2231] = 103;
    exp_48_ram[2232] = 46;
    exp_48_ram[2233] = 39;
    exp_48_ram[2234] = 39;
    exp_48_ram[2235] = 7;
    exp_48_ram[2236] = 32;
    exp_48_ram[2237] = 39;
    exp_48_ram[2238] = 32;
    exp_48_ram[2239] = 215;
    exp_48_ram[2240] = 34;
    exp_48_ram[2241] = 39;
    exp_48_ram[2242] = 23;
    exp_48_ram[2243] = 133;
    exp_48_ram[2244] = 5;
    exp_48_ram[2245] = 16;
    exp_48_ram[2246] = 7;
    exp_48_ram[2247] = 135;
    exp_48_ram[2248] = 46;
    exp_48_ram[2249] = 32;
    exp_48_ram[2250] = 39;
    exp_48_ram[2251] = 38;
    exp_48_ram[2252] = 39;
    exp_48_ram[2253] = 32;
    exp_48_ram[2254] = 215;
    exp_48_ram[2255] = 34;
    exp_48_ram[2256] = 39;
    exp_48_ram[2257] = 5;
    exp_48_ram[2258] = 133;
    exp_48_ram[2259] = 16;
    exp_48_ram[2260] = 7;
    exp_48_ram[2261] = 135;
    exp_48_ram[2262] = 46;
    exp_48_ram[2263] = 32;
    exp_48_ram[2264] = 39;
    exp_48_ram[2265] = 36;
    exp_48_ram[2266] = 39;
    exp_48_ram[2267] = 32;
    exp_48_ram[2268] = 215;
    exp_48_ram[2269] = 34;
    exp_48_ram[2270] = 39;
    exp_48_ram[2271] = 34;
    exp_48_ram[2272] = 39;
    exp_48_ram[2273] = 46;
    exp_48_ram[2274] = 35;
    exp_48_ram[2275] = 40;
    exp_48_ram[2276] = 40;
    exp_48_ram[2277] = 37;
    exp_48_ram[2278] = 37;
    exp_48_ram[2279] = 38;
    exp_48_ram[2280] = 38;
    exp_48_ram[2281] = 39;
    exp_48_ram[2282] = 160;
    exp_48_ram[2283] = 162;
    exp_48_ram[2284] = 164;
    exp_48_ram[2285] = 166;
    exp_48_ram[2286] = 168;
    exp_48_ram[2287] = 170;
    exp_48_ram[2288] = 172;
    exp_48_ram[2289] = 174;
    exp_48_ram[2290] = 160;
    exp_48_ram[2291] = 37;
    exp_48_ram[2292] = 32;
    exp_48_ram[2293] = 36;
    exp_48_ram[2294] = 41;
    exp_48_ram[2295] = 41;
    exp_48_ram[2296] = 42;
    exp_48_ram[2297] = 42;
    exp_48_ram[2298] = 43;
    exp_48_ram[2299] = 43;
    exp_48_ram[2300] = 44;
    exp_48_ram[2301] = 44;
    exp_48_ram[2302] = 1;
    exp_48_ram[2303] = 128;
    exp_48_ram[2304] = 1;
    exp_48_ram[2305] = 46;
    exp_48_ram[2306] = 44;
    exp_48_ram[2307] = 42;
    exp_48_ram[2308] = 40;
    exp_48_ram[2309] = 38;
    exp_48_ram[2310] = 4;
    exp_48_ram[2311] = 46;
    exp_48_ram[2312] = 7;
    exp_48_ram[2313] = 8;
    exp_48_ram[2314] = 44;
    exp_48_ram[2315] = 46;
    exp_48_ram[2316] = 39;
    exp_48_ram[2317] = 167;
    exp_48_ram[2318] = 167;
    exp_48_ram[2319] = 40;
    exp_48_ram[2320] = 42;
    exp_48_ram[2321] = 37;
    exp_48_ram[2322] = 37;
    exp_48_ram[2323] = 224;
    exp_48_ram[2324] = 7;
    exp_48_ram[2325] = 140;
    exp_48_ram[2326] = 23;
    exp_48_ram[2327] = 7;
    exp_48_ram[2328] = 7;
    exp_48_ram[2329] = 44;
    exp_48_ram[2330] = 46;
    exp_48_ram[2331] = 71;
    exp_48_ram[2332] = 167;
    exp_48_ram[2333] = 137;
    exp_48_ram[2334] = 215;
    exp_48_ram[2335] = 137;
    exp_48_ram[2336] = 38;
    exp_48_ram[2337] = 38;
    exp_48_ram[2338] = 7;
    exp_48_ram[2339] = 5;
    exp_48_ram[2340] = 181;
    exp_48_ram[2341] = 135;
    exp_48_ram[2342] = 134;
    exp_48_ram[2343] = 135;
    exp_48_ram[2344] = 5;
    exp_48_ram[2345] = 133;
    exp_48_ram[2346] = 38;
    exp_48_ram[2347] = 38;
    exp_48_ram[2348] = 7;
    exp_48_ram[2349] = 8;
    exp_48_ram[2350] = 56;
    exp_48_ram[2351] = 135;
    exp_48_ram[2352] = 6;
    exp_48_ram[2353] = 135;
    exp_48_ram[2354] = 36;
    exp_48_ram[2355] = 38;
    exp_48_ram[2356] = 71;
    exp_48_ram[2357] = 132;
    exp_48_ram[2358] = 7;
    exp_48_ram[2359] = 37;
    exp_48_ram[2360] = 38;
    exp_48_ram[2361] = 133;
    exp_48_ram[2362] = 240;
    exp_48_ram[2363] = 35;
    exp_48_ram[2364] = 40;
    exp_48_ram[2365] = 40;
    exp_48_ram[2366] = 37;
    exp_48_ram[2367] = 37;
    exp_48_ram[2368] = 38;
    exp_48_ram[2369] = 38;
    exp_48_ram[2370] = 39;
    exp_48_ram[2371] = 39;
    exp_48_ram[2372] = 160;
    exp_48_ram[2373] = 162;
    exp_48_ram[2374] = 164;
    exp_48_ram[2375] = 166;
    exp_48_ram[2376] = 168;
    exp_48_ram[2377] = 170;
    exp_48_ram[2378] = 172;
    exp_48_ram[2379] = 174;
    exp_48_ram[2380] = 160;
    exp_48_ram[2381] = 37;
    exp_48_ram[2382] = 37;
    exp_48_ram[2383] = 224;
    exp_48_ram[2384] = 7;
    exp_48_ram[2385] = 71;
    exp_48_ram[2386] = 135;
    exp_48_ram[2387] = 160;
    exp_48_ram[2388] = 71;
    exp_48_ram[2389] = 135;
    exp_48_ram[2390] = 133;
    exp_48_ram[2391] = 32;
    exp_48_ram[2392] = 36;
    exp_48_ram[2393] = 36;
    exp_48_ram[2394] = 41;
    exp_48_ram[2395] = 41;
    exp_48_ram[2396] = 1;
    exp_48_ram[2397] = 128;
    exp_48_ram[2398] = 1;
    exp_48_ram[2399] = 38;
    exp_48_ram[2400] = 36;
    exp_48_ram[2401] = 4;
    exp_48_ram[2402] = 46;
    exp_48_ram[2403] = 38;
    exp_48_ram[2404] = 37;
    exp_48_ram[2405] = 224;
    exp_48_ram[2406] = 7;
    exp_48_ram[2407] = 5;
    exp_48_ram[2408] = 71;
    exp_48_ram[2409] = 135;
    exp_48_ram[2410] = 7;
    exp_48_ram[2411] = 234;
    exp_48_ram[2412] = 39;
    exp_48_ram[2413] = 7;
    exp_48_ram[2414] = 151;
    exp_48_ram[2415] = 135;
    exp_48_ram[2416] = 151;
    exp_48_ram[2417] = 38;
    exp_48_ram[2418] = 71;
    exp_48_ram[2419] = 39;
    exp_48_ram[2420] = 7;
    exp_48_ram[2421] = 135;
    exp_48_ram[2422] = 38;
    exp_48_ram[2423] = 240;
    exp_48_ram[2424] = 0;
    exp_48_ram[2425] = 39;
    exp_48_ram[2426] = 133;
    exp_48_ram[2427] = 32;
    exp_48_ram[2428] = 36;
    exp_48_ram[2429] = 1;
    exp_48_ram[2430] = 128;
    exp_48_ram[2431] = 1;
    exp_48_ram[2432] = 38;
    exp_48_ram[2433] = 36;
    exp_48_ram[2434] = 4;
    exp_48_ram[2435] = 71;
    exp_48_ram[2436] = 167;
    exp_48_ram[2437] = 133;
    exp_48_ram[2438] = 240;
    exp_48_ram[2439] = 7;
    exp_48_ram[2440] = 133;
    exp_48_ram[2441] = 32;
    exp_48_ram[2442] = 36;
    exp_48_ram[2443] = 1;
    exp_48_ram[2444] = 128;
    exp_48_ram[2445] = 1;
    exp_48_ram[2446] = 38;
    exp_48_ram[2447] = 36;
    exp_48_ram[2448] = 4;
    exp_48_ram[2449] = 46;
    exp_48_ram[2450] = 44;
    exp_48_ram[2451] = 42;
    exp_48_ram[2452] = 215;
    exp_48_ram[2453] = 135;
    exp_48_ram[2454] = 38;
    exp_48_ram[2455] = 7;
    exp_48_ram[2456] = 36;
    exp_48_ram[2457] = 34;
    exp_48_ram[2458] = 0;
    exp_48_ram[2459] = 39;
    exp_48_ram[2460] = 39;
    exp_48_ram[2461] = 87;
    exp_48_ram[2462] = 1;
    exp_48_ram[2463] = 71;
    exp_48_ram[2464] = 156;
    exp_48_ram[2465] = 39;
    exp_48_ram[2466] = 152;
    exp_48_ram[2467] = 39;
    exp_48_ram[2468] = 7;
    exp_48_ram[2469] = 18;
    exp_48_ram[2470] = 71;
    exp_48_ram[2471] = 135;
    exp_48_ram[2472] = 37;
    exp_48_ram[2473] = 133;
    exp_48_ram[2474] = 224;
    exp_48_ram[2475] = 7;
    exp_48_ram[2476] = 34;
    exp_48_ram[2477] = 0;
    exp_48_ram[2478] = 39;
    exp_48_ram[2479] = 39;
    exp_48_ram[2480] = 108;
    exp_48_ram[2481] = 71;
    exp_48_ram[2482] = 135;
    exp_48_ram[2483] = 37;
    exp_48_ram[2484] = 133;
    exp_48_ram[2485] = 224;
    exp_48_ram[2486] = 39;
    exp_48_ram[2487] = 39;
    exp_48_ram[2488] = 119;
    exp_48_ram[2489] = 46;
    exp_48_ram[2490] = 39;
    exp_48_ram[2491] = 7;
    exp_48_ram[2492] = 87;
    exp_48_ram[2493] = 38;
    exp_48_ram[2494] = 39;
    exp_48_ram[2495] = 135;
    exp_48_ram[2496] = 36;
    exp_48_ram[2497] = 39;
    exp_48_ram[2498] = 146;
    exp_48_ram[2499] = 0;
    exp_48_ram[2500] = 0;
    exp_48_ram[2501] = 32;
    exp_48_ram[2502] = 36;
    exp_48_ram[2503] = 1;
    exp_48_ram[2504] = 128;
    exp_48_ram[2505] = 1;
    exp_48_ram[2506] = 46;
    exp_48_ram[2507] = 44;
    exp_48_ram[2508] = 4;
    exp_48_ram[2509] = 38;
    exp_48_ram[2510] = 36;
    exp_48_ram[2511] = 39;
    exp_48_ram[2512] = 38;
    exp_48_ram[2513] = 71;
    exp_48_ram[2514] = 167;
    exp_48_ram[2515] = 134;
    exp_48_ram[2516] = 133;
    exp_48_ram[2517] = 5;
    exp_48_ram[2518] = 240;
    exp_48_ram[2519] = 0;
    exp_48_ram[2520] = 32;
    exp_48_ram[2521] = 36;
    exp_48_ram[2522] = 1;
    exp_48_ram[2523] = 128;
    exp_48_ram[2524] = 1;
    exp_48_ram[2525] = 38;
    exp_48_ram[2526] = 36;
    exp_48_ram[2527] = 34;
    exp_48_ram[2528] = 32;
    exp_48_ram[2529] = 4;
    exp_48_ram[2530] = 46;
    exp_48_ram[2531] = 224;
    exp_48_ram[2532] = 36;
    exp_48_ram[2533] = 38;
    exp_48_ram[2534] = 0;
    exp_48_ram[2535] = 224;
    exp_48_ram[2536] = 6;
    exp_48_ram[2537] = 134;
    exp_48_ram[2538] = 37;
    exp_48_ram[2539] = 37;
    exp_48_ram[2540] = 7;
    exp_48_ram[2541] = 8;
    exp_48_ram[2542] = 56;
    exp_48_ram[2543] = 135;
    exp_48_ram[2544] = 134;
    exp_48_ram[2545] = 135;
    exp_48_ram[2546] = 38;
    exp_48_ram[2547] = 137;
    exp_48_ram[2548] = 9;
    exp_48_ram[2549] = 134;
    exp_48_ram[2550] = 134;
    exp_48_ram[2551] = 224;
    exp_48_ram[2552] = 134;
    exp_48_ram[2553] = 134;
    exp_48_ram[2554] = 24;
    exp_48_ram[2555] = 6;
    exp_48_ram[2556] = 7;
    exp_48_ram[2557] = 228;
    exp_48_ram[2558] = 0;
    exp_48_ram[2559] = 133;
    exp_48_ram[2560] = 32;
    exp_48_ram[2561] = 36;
    exp_48_ram[2562] = 41;
    exp_48_ram[2563] = 41;
    exp_48_ram[2564] = 1;
    exp_48_ram[2565] = 128;
    exp_48_ram[2566] = 1;
    exp_48_ram[2567] = 38;
    exp_48_ram[2568] = 36;
    exp_48_ram[2569] = 4;
    exp_48_ram[2570] = 23;
    exp_48_ram[2571] = 133;
    exp_48_ram[2572] = 224;
    exp_48_ram[2573] = 0;
    exp_48_ram[2574] = 32;
    exp_48_ram[2575] = 36;
    exp_48_ram[2576] = 1;
    exp_48_ram[2577] = 128;
    exp_48_ram[2578] = 1;
    exp_48_ram[2579] = 46;
    exp_48_ram[2580] = 44;
    exp_48_ram[2581] = 4;
    exp_48_ram[2582] = 23;
    exp_48_ram[2583] = 133;
    exp_48_ram[2584] = 224;
    exp_48_ram[2585] = 7;
    exp_48_ram[2586] = 38;
    exp_48_ram[2587] = 36;
    exp_48_ram[2588] = 0;
    exp_48_ram[2589] = 5;
    exp_48_ram[2590] = 37;
    exp_48_ram[2591] = 240;
    exp_48_ram[2592] = 5;
    exp_48_ram[2593] = 224;
    exp_48_ram[2594] = 0;
    exp_48_ram[2595] = 39;
    exp_48_ram[2596] = 151;
    exp_48_ram[2597] = 38;
    exp_48_ram[2598] = 71;
    exp_48_ram[2599] = 167;
    exp_48_ram[2600] = 133;
    exp_48_ram[2601] = 37;
    exp_48_ram[2602] = 224;
    exp_48_ram[2603] = 71;
    exp_48_ram[2604] = 167;
    exp_48_ram[2605] = 7;
    exp_48_ram[2606] = 87;
    exp_48_ram[2607] = 133;
    exp_48_ram[2608] = 240;
    exp_48_ram[2609] = 39;
    exp_48_ram[2610] = 7;
    exp_48_ram[2611] = 208;
    exp_48_ram[2612] = 0;
    exp_48_ram[2613] = 39;
    exp_48_ram[2614] = 215;
    exp_48_ram[2615] = 38;
    exp_48_ram[2616] = 71;
    exp_48_ram[2617] = 167;
    exp_48_ram[2618] = 133;
    exp_48_ram[2619] = 37;
    exp_48_ram[2620] = 224;
    exp_48_ram[2621] = 71;
    exp_48_ram[2622] = 167;
    exp_48_ram[2623] = 7;
    exp_48_ram[2624] = 87;
    exp_48_ram[2625] = 133;
    exp_48_ram[2626] = 240;
    exp_48_ram[2627] = 39;
    exp_48_ram[2628] = 7;
    exp_48_ram[2629] = 192;
    exp_48_ram[2630] = 39;
    exp_48_ram[2631] = 135;
    exp_48_ram[2632] = 36;
    exp_48_ram[2633] = 39;
    exp_48_ram[2634] = 7;
    exp_48_ram[2635] = 212;
    exp_48_ram[2636] = 71;
    exp_48_ram[2637] = 167;
    exp_48_ram[2638] = 133;
    exp_48_ram[2639] = 5;
    exp_48_ram[2640] = 224;
    exp_48_ram[2641] = 0;
    exp_48_ram[2642] = 32;
    exp_48_ram[2643] = 36;
    exp_48_ram[2644] = 1;
    exp_48_ram[2645] = 128;
    exp_48_ram[2646] = 1;
    exp_48_ram[2647] = 46;
    exp_48_ram[2648] = 44;
    exp_48_ram[2649] = 4;
    exp_48_ram[2650] = 23;
    exp_48_ram[2651] = 133;
    exp_48_ram[2652] = 224;
    exp_48_ram[2653] = 36;
    exp_48_ram[2654] = 0;
    exp_48_ram[2655] = 5;
    exp_48_ram[2656] = 37;
    exp_48_ram[2657] = 240;
    exp_48_ram[2658] = 5;
    exp_48_ram[2659] = 224;
    exp_48_ram[2660] = 38;
    exp_48_ram[2661] = 0;
    exp_48_ram[2662] = 71;
    exp_48_ram[2663] = 167;
    exp_48_ram[2664] = 133;
    exp_48_ram[2665] = 37;
    exp_48_ram[2666] = 224;
    exp_48_ram[2667] = 71;
    exp_48_ram[2668] = 167;
    exp_48_ram[2669] = 7;
    exp_48_ram[2670] = 87;
    exp_48_ram[2671] = 133;
    exp_48_ram[2672] = 240;
    exp_48_ram[2673] = 39;
    exp_48_ram[2674] = 135;
    exp_48_ram[2675] = 38;
    exp_48_ram[2676] = 39;
    exp_48_ram[2677] = 7;
    exp_48_ram[2678] = 208;
    exp_48_ram[2679] = 7;
    exp_48_ram[2680] = 38;
    exp_48_ram[2681] = 0;
    exp_48_ram[2682] = 71;
    exp_48_ram[2683] = 167;
    exp_48_ram[2684] = 133;
    exp_48_ram[2685] = 37;
    exp_48_ram[2686] = 224;
    exp_48_ram[2687] = 71;
    exp_48_ram[2688] = 167;
    exp_48_ram[2689] = 7;
    exp_48_ram[2690] = 87;
    exp_48_ram[2691] = 133;
    exp_48_ram[2692] = 240;
    exp_48_ram[2693] = 39;
    exp_48_ram[2694] = 135;
    exp_48_ram[2695] = 38;
    exp_48_ram[2696] = 39;
    exp_48_ram[2697] = 210;
    exp_48_ram[2698] = 39;
    exp_48_ram[2699] = 135;
    exp_48_ram[2700] = 36;
    exp_48_ram[2701] = 39;
    exp_48_ram[2702] = 7;
    exp_48_ram[2703] = 208;
    exp_48_ram[2704] = 71;
    exp_48_ram[2705] = 167;
    exp_48_ram[2706] = 133;
    exp_48_ram[2707] = 5;
    exp_48_ram[2708] = 224;
    exp_48_ram[2709] = 0;
    exp_48_ram[2710] = 32;
    exp_48_ram[2711] = 36;
    exp_48_ram[2712] = 1;
    exp_48_ram[2713] = 128;
    exp_48_ram[2714] = 1;
    exp_48_ram[2715] = 38;
    exp_48_ram[2716] = 36;
    exp_48_ram[2717] = 34;
    exp_48_ram[2718] = 32;
    exp_48_ram[2719] = 46;
    exp_48_ram[2720] = 44;
    exp_48_ram[2721] = 42;
    exp_48_ram[2722] = 40;
    exp_48_ram[2723] = 38;
    exp_48_ram[2724] = 36;
    exp_48_ram[2725] = 34;
    exp_48_ram[2726] = 32;
    exp_48_ram[2727] = 4;
    exp_48_ram[2728] = 7;
    exp_48_ram[2729] = 46;
    exp_48_ram[2730] = 7;
    exp_48_ram[2731] = 7;
    exp_48_ram[2732] = 40;
    exp_48_ram[2733] = 42;
    exp_48_ram[2734] = 224;
    exp_48_ram[2735] = 32;
    exp_48_ram[2736] = 34;
    exp_48_ram[2737] = 38;
    exp_48_ram[2738] = 0;
    exp_48_ram[2739] = 39;
    exp_48_ram[2740] = 87;
    exp_48_ram[2741] = 135;
    exp_48_ram[2742] = 7;
    exp_48_ram[2743] = 46;
    exp_48_ram[2744] = 39;
    exp_48_ram[2745] = 87;
    exp_48_ram[2746] = 135;
    exp_48_ram[2747] = 7;
    exp_48_ram[2748] = 46;
    exp_48_ram[2749] = 39;
    exp_48_ram[2750] = 87;
    exp_48_ram[2751] = 135;
    exp_48_ram[2752] = 7;
    exp_48_ram[2753] = 46;
    exp_48_ram[2754] = 39;
    exp_48_ram[2755] = 87;
    exp_48_ram[2756] = 135;
    exp_48_ram[2757] = 7;
    exp_48_ram[2758] = 46;
    exp_48_ram[2759] = 39;
    exp_48_ram[2760] = 135;
    exp_48_ram[2761] = 38;
    exp_48_ram[2762] = 224;
    exp_48_ram[2763] = 6;
    exp_48_ram[2764] = 134;
    exp_48_ram[2765] = 37;
    exp_48_ram[2766] = 37;
    exp_48_ram[2767] = 7;
    exp_48_ram[2768] = 8;
    exp_48_ram[2769] = 56;
    exp_48_ram[2770] = 135;
    exp_48_ram[2771] = 134;
    exp_48_ram[2772] = 135;
    exp_48_ram[2773] = 70;
    exp_48_ram[2774] = 166;
    exp_48_ram[2775] = 36;
    exp_48_ram[2776] = 38;
    exp_48_ram[2777] = 37;
    exp_48_ram[2778] = 37;
    exp_48_ram[2779] = 134;
    exp_48_ram[2780] = 134;
    exp_48_ram[2781] = 236;
    exp_48_ram[2782] = 134;
    exp_48_ram[2783] = 134;
    exp_48_ram[2784] = 24;
    exp_48_ram[2785] = 6;
    exp_48_ram[2786] = 7;
    exp_48_ram[2787] = 224;
    exp_48_ram[2788] = 39;
    exp_48_ram[2789] = 5;
    exp_48_ram[2790] = 133;
    exp_48_ram[2791] = 240;
    exp_48_ram[2792] = 23;
    exp_48_ram[2793] = 133;
    exp_48_ram[2794] = 224;
    exp_48_ram[2795] = 224;
    exp_48_ram[2796] = 32;
    exp_48_ram[2797] = 34;
    exp_48_ram[2798] = 38;
    exp_48_ram[2799] = 0;
    exp_48_ram[2800] = 39;
    exp_48_ram[2801] = 39;
    exp_48_ram[2802] = 86;
    exp_48_ram[2803] = 134;
    exp_48_ram[2804] = 134;
    exp_48_ram[2805] = 6;
    exp_48_ram[2806] = 6;
    exp_48_ram[2807] = 6;
    exp_48_ram[2808] = 86;
    exp_48_ram[2809] = 134;
    exp_48_ram[2810] = 5;
    exp_48_ram[2811] = 57;
    exp_48_ram[2812] = 137;
    exp_48_ram[2813] = 7;
    exp_48_ram[2814] = 137;
    exp_48_ram[2815] = 40;
    exp_48_ram[2816] = 42;
    exp_48_ram[2817] = 39;
    exp_48_ram[2818] = 39;
    exp_48_ram[2819] = 86;
    exp_48_ram[2820] = 134;
    exp_48_ram[2821] = 134;
    exp_48_ram[2822] = 6;
    exp_48_ram[2823] = 6;
    exp_48_ram[2824] = 6;
    exp_48_ram[2825] = 86;
    exp_48_ram[2826] = 134;
    exp_48_ram[2827] = 5;
    exp_48_ram[2828] = 58;
    exp_48_ram[2829] = 138;
    exp_48_ram[2830] = 7;
    exp_48_ram[2831] = 138;
    exp_48_ram[2832] = 40;
    exp_48_ram[2833] = 42;
    exp_48_ram[2834] = 39;
    exp_48_ram[2835] = 39;
    exp_48_ram[2836] = 86;
    exp_48_ram[2837] = 134;
    exp_48_ram[2838] = 134;
    exp_48_ram[2839] = 6;
    exp_48_ram[2840] = 6;
    exp_48_ram[2841] = 6;
    exp_48_ram[2842] = 86;
    exp_48_ram[2843] = 134;
    exp_48_ram[2844] = 5;
    exp_48_ram[2845] = 59;
    exp_48_ram[2846] = 139;
    exp_48_ram[2847] = 7;
    exp_48_ram[2848] = 139;
    exp_48_ram[2849] = 40;
    exp_48_ram[2850] = 42;
    exp_48_ram[2851] = 39;
    exp_48_ram[2852] = 39;
    exp_48_ram[2853] = 86;
    exp_48_ram[2854] = 134;
    exp_48_ram[2855] = 134;
    exp_48_ram[2856] = 6;
    exp_48_ram[2857] = 6;
    exp_48_ram[2858] = 6;
    exp_48_ram[2859] = 86;
    exp_48_ram[2860] = 134;
    exp_48_ram[2861] = 5;
    exp_48_ram[2862] = 60;
    exp_48_ram[2863] = 140;
    exp_48_ram[2864] = 7;
    exp_48_ram[2865] = 140;
    exp_48_ram[2866] = 40;
    exp_48_ram[2867] = 42;
    exp_48_ram[2868] = 39;
    exp_48_ram[2869] = 135;
    exp_48_ram[2870] = 38;
    exp_48_ram[2871] = 224;
    exp_48_ram[2872] = 6;
    exp_48_ram[2873] = 134;
    exp_48_ram[2874] = 37;
    exp_48_ram[2875] = 37;
    exp_48_ram[2876] = 7;
    exp_48_ram[2877] = 8;
    exp_48_ram[2878] = 56;
    exp_48_ram[2879] = 135;
    exp_48_ram[2880] = 134;
    exp_48_ram[2881] = 135;
    exp_48_ram[2882] = 70;
    exp_48_ram[2883] = 166;
    exp_48_ram[2884] = 32;
    exp_48_ram[2885] = 34;
    exp_48_ram[2886] = 37;
    exp_48_ram[2887] = 37;
    exp_48_ram[2888] = 134;
    exp_48_ram[2889] = 134;
    exp_48_ram[2890] = 236;
    exp_48_ram[2891] = 134;
    exp_48_ram[2892] = 134;
    exp_48_ram[2893] = 24;
    exp_48_ram[2894] = 6;
    exp_48_ram[2895] = 7;
    exp_48_ram[2896] = 224;
    exp_48_ram[2897] = 39;
    exp_48_ram[2898] = 5;
    exp_48_ram[2899] = 133;
    exp_48_ram[2900] = 240;
    exp_48_ram[2901] = 23;
    exp_48_ram[2902] = 133;
    exp_48_ram[2903] = 224;
    exp_48_ram[2904] = 224;
    exp_48_ram[2905] = 32;
    exp_48_ram[2906] = 34;
    exp_48_ram[2907] = 38;
    exp_48_ram[2908] = 0;
    exp_48_ram[2909] = 39;
    exp_48_ram[2910] = 87;
    exp_48_ram[2911] = 135;
    exp_48_ram[2912] = 87;
    exp_48_ram[2913] = 46;
    exp_48_ram[2914] = 39;
    exp_48_ram[2915] = 87;
    exp_48_ram[2916] = 135;
    exp_48_ram[2917] = 87;
    exp_48_ram[2918] = 46;
    exp_48_ram[2919] = 39;
    exp_48_ram[2920] = 87;
    exp_48_ram[2921] = 135;
    exp_48_ram[2922] = 87;
    exp_48_ram[2923] = 46;
    exp_48_ram[2924] = 39;
    exp_48_ram[2925] = 87;
    exp_48_ram[2926] = 135;
    exp_48_ram[2927] = 87;
    exp_48_ram[2928] = 46;
    exp_48_ram[2929] = 39;
    exp_48_ram[2930] = 135;
    exp_48_ram[2931] = 38;
    exp_48_ram[2932] = 224;
    exp_48_ram[2933] = 6;
    exp_48_ram[2934] = 134;
    exp_48_ram[2935] = 37;
    exp_48_ram[2936] = 37;
    exp_48_ram[2937] = 7;
    exp_48_ram[2938] = 8;
    exp_48_ram[2939] = 56;
    exp_48_ram[2940] = 135;
    exp_48_ram[2941] = 134;
    exp_48_ram[2942] = 135;
    exp_48_ram[2943] = 70;
    exp_48_ram[2944] = 166;
    exp_48_ram[2945] = 44;
    exp_48_ram[2946] = 46;
    exp_48_ram[2947] = 37;
    exp_48_ram[2948] = 37;
    exp_48_ram[2949] = 134;
    exp_48_ram[2950] = 134;
    exp_48_ram[2951] = 236;
    exp_48_ram[2952] = 134;
    exp_48_ram[2953] = 134;
    exp_48_ram[2954] = 24;
    exp_48_ram[2955] = 6;
    exp_48_ram[2956] = 7;
    exp_48_ram[2957] = 224;
    exp_48_ram[2958] = 39;
    exp_48_ram[2959] = 5;
    exp_48_ram[2960] = 133;
    exp_48_ram[2961] = 240;
    exp_48_ram[2962] = 23;
    exp_48_ram[2963] = 133;
    exp_48_ram[2964] = 208;
    exp_48_ram[2965] = 224;
    exp_48_ram[2966] = 32;
    exp_48_ram[2967] = 34;
    exp_48_ram[2968] = 38;
    exp_48_ram[2969] = 0;
    exp_48_ram[2970] = 39;
    exp_48_ram[2971] = 39;
    exp_48_ram[2972] = 86;
    exp_48_ram[2973] = 6;
    exp_48_ram[2974] = 6;
    exp_48_ram[2975] = 5;
    exp_48_ram[2976] = 133;
    exp_48_ram[2977] = 208;
    exp_48_ram[2978] = 7;
    exp_48_ram[2979] = 135;
    exp_48_ram[2980] = 40;
    exp_48_ram[2981] = 42;
    exp_48_ram[2982] = 39;
    exp_48_ram[2983] = 39;
    exp_48_ram[2984] = 86;
    exp_48_ram[2985] = 6;
    exp_48_ram[2986] = 6;
    exp_48_ram[2987] = 5;
    exp_48_ram[2988] = 133;
    exp_48_ram[2989] = 208;
    exp_48_ram[2990] = 7;
    exp_48_ram[2991] = 135;
    exp_48_ram[2992] = 40;
    exp_48_ram[2993] = 42;
    exp_48_ram[2994] = 39;
    exp_48_ram[2995] = 39;
    exp_48_ram[2996] = 86;
    exp_48_ram[2997] = 6;
    exp_48_ram[2998] = 6;
    exp_48_ram[2999] = 5;
    exp_48_ram[3000] = 133;
    exp_48_ram[3001] = 208;
    exp_48_ram[3002] = 7;
    exp_48_ram[3003] = 135;
    exp_48_ram[3004] = 40;
    exp_48_ram[3005] = 42;
    exp_48_ram[3006] = 39;
    exp_48_ram[3007] = 39;
    exp_48_ram[3008] = 86;
    exp_48_ram[3009] = 6;
    exp_48_ram[3010] = 6;
    exp_48_ram[3011] = 5;
    exp_48_ram[3012] = 133;
    exp_48_ram[3013] = 208;
    exp_48_ram[3014] = 7;
    exp_48_ram[3015] = 135;
    exp_48_ram[3016] = 40;
    exp_48_ram[3017] = 42;
    exp_48_ram[3018] = 39;
    exp_48_ram[3019] = 135;
    exp_48_ram[3020] = 38;
    exp_48_ram[3021] = 224;
    exp_48_ram[3022] = 6;
    exp_48_ram[3023] = 134;
    exp_48_ram[3024] = 37;
    exp_48_ram[3025] = 37;
    exp_48_ram[3026] = 7;
    exp_48_ram[3027] = 8;
    exp_48_ram[3028] = 56;
    exp_48_ram[3029] = 135;
    exp_48_ram[3030] = 134;
    exp_48_ram[3031] = 135;
    exp_48_ram[3032] = 70;
    exp_48_ram[3033] = 166;
    exp_48_ram[3034] = 141;
    exp_48_ram[3035] = 13;
    exp_48_ram[3036] = 134;
    exp_48_ram[3037] = 134;
    exp_48_ram[3038] = 232;
    exp_48_ram[3039] = 134;
    exp_48_ram[3040] = 134;
    exp_48_ram[3041] = 24;
    exp_48_ram[3042] = 6;
    exp_48_ram[3043] = 7;
    exp_48_ram[3044] = 236;
    exp_48_ram[3045] = 39;
    exp_48_ram[3046] = 5;
    exp_48_ram[3047] = 133;
    exp_48_ram[3048] = 240;
    exp_48_ram[3049] = 23;
    exp_48_ram[3050] = 133;
    exp_48_ram[3051] = 208;
    exp_48_ram[3052] = 0;
    exp_48_ram[3053] = 32;
    exp_48_ram[3054] = 36;
    exp_48_ram[3055] = 41;
    exp_48_ram[3056] = 41;
    exp_48_ram[3057] = 42;
    exp_48_ram[3058] = 42;
    exp_48_ram[3059] = 43;
    exp_48_ram[3060] = 43;
    exp_48_ram[3061] = 44;
    exp_48_ram[3062] = 44;
    exp_48_ram[3063] = 45;
    exp_48_ram[3064] = 45;
    exp_48_ram[3065] = 1;
    exp_48_ram[3066] = 128;
    exp_48_ram[3067] = 1;
    exp_48_ram[3068] = 46;
    exp_48_ram[3069] = 44;
    exp_48_ram[3070] = 42;
    exp_48_ram[3071] = 40;
    exp_48_ram[3072] = 38;
    exp_48_ram[3073] = 36;
    exp_48_ram[3074] = 4;
    exp_48_ram[3075] = 23;
    exp_48_ram[3076] = 133;
    exp_48_ram[3077] = 208;
    exp_48_ram[3078] = 240;
    exp_48_ram[3079] = 7;
    exp_48_ram[3080] = 135;
    exp_48_ram[3081] = 34;
    exp_48_ram[3082] = 23;
    exp_48_ram[3083] = 133;
    exp_48_ram[3084] = 208;
    exp_48_ram[3085] = 240;
    exp_48_ram[3086] = 7;
    exp_48_ram[3087] = 135;
    exp_48_ram[3088] = 32;
    exp_48_ram[3089] = 23;
    exp_48_ram[3090] = 133;
    exp_48_ram[3091] = 208;
    exp_48_ram[3092] = 240;
    exp_48_ram[3093] = 7;
    exp_48_ram[3094] = 46;
    exp_48_ram[3095] = 23;
    exp_48_ram[3096] = 133;
    exp_48_ram[3097] = 208;
    exp_48_ram[3098] = 240;
    exp_48_ram[3099] = 7;
    exp_48_ram[3100] = 44;
    exp_48_ram[3101] = 23;
    exp_48_ram[3102] = 133;
    exp_48_ram[3103] = 208;
    exp_48_ram[3104] = 240;
    exp_48_ram[3105] = 7;
    exp_48_ram[3106] = 42;
    exp_48_ram[3107] = 7;
    exp_48_ram[3108] = 40;
    exp_48_ram[3109] = 7;
    exp_48_ram[3110] = 40;
    exp_48_ram[3111] = 7;
    exp_48_ram[3112] = 133;
    exp_48_ram[3113] = 224;
    exp_48_ram[3114] = 7;
    exp_48_ram[3115] = 135;
    exp_48_ram[3116] = 36;
    exp_48_ram[3117] = 38;
    exp_48_ram[3118] = 39;
    exp_48_ram[3119] = 39;
    exp_48_ram[3120] = 5;
    exp_48_ram[3121] = 133;
    exp_48_ram[3122] = 224;
    exp_48_ram[3123] = 224;
    exp_48_ram[3124] = 44;
    exp_48_ram[3125] = 46;
    exp_48_ram[3126] = 42;
    exp_48_ram[3127] = 0;
    exp_48_ram[3128] = 0;
    exp_48_ram[3129] = 224;
    exp_48_ram[3130] = 7;
    exp_48_ram[3131] = 135;
    exp_48_ram[3132] = 38;
    exp_48_ram[3133] = 38;
    exp_48_ram[3134] = 5;
    exp_48_ram[3135] = 133;
    exp_48_ram[3136] = 224;
    exp_48_ram[3137] = 10;
    exp_48_ram[3138] = 138;
    exp_48_ram[3139] = 71;
    exp_48_ram[3140] = 167;
    exp_48_ram[3141] = 133;
    exp_48_ram[3142] = 208;
    exp_48_ram[3143] = 7;
    exp_48_ram[3144] = 135;
    exp_48_ram[3145] = 6;
    exp_48_ram[3146] = 134;
    exp_48_ram[3147] = 5;
    exp_48_ram[3148] = 133;
    exp_48_ram[3149] = 208;
    exp_48_ram[3150] = 7;
    exp_48_ram[3151] = 196;
    exp_48_ram[3152] = 71;
    exp_48_ram[3153] = 167;
    exp_48_ram[3154] = 137;
    exp_48_ram[3155] = 9;
    exp_48_ram[3156] = 38;
    exp_48_ram[3157] = 38;
    exp_48_ram[3158] = 7;
    exp_48_ram[3159] = 5;
    exp_48_ram[3160] = 181;
    exp_48_ram[3161] = 135;
    exp_48_ram[3162] = 134;
    exp_48_ram[3163] = 135;
    exp_48_ram[3164] = 44;
    exp_48_ram[3165] = 46;
    exp_48_ram[3166] = 5;
    exp_48_ram[3167] = 224;
    exp_48_ram[3168] = 7;
    exp_48_ram[3169] = 135;
    exp_48_ram[3170] = 36;
    exp_48_ram[3171] = 38;
    exp_48_ram[3172] = 7;
    exp_48_ram[3173] = 133;
    exp_48_ram[3174] = 224;
    exp_48_ram[3175] = 7;
    exp_48_ram[3176] = 133;
    exp_48_ram[3177] = 208;
    exp_48_ram[3178] = 39;
    exp_48_ram[3179] = 135;
    exp_48_ram[3180] = 42;
    exp_48_ram[3181] = 39;
    exp_48_ram[3182] = 7;
    exp_48_ram[3183] = 210;
    exp_48_ram[3184] = 0;
    exp_48_ram[3185] = 0;
    exp_48_ram[3186] = 32;
    exp_48_ram[3187] = 36;
    exp_48_ram[3188] = 41;
    exp_48_ram[3189] = 41;
    exp_48_ram[3190] = 42;
    exp_48_ram[3191] = 42;
    exp_48_ram[3192] = 1;
    exp_48_ram[3193] = 128;
    exp_48_ram[3194] = 1;
    exp_48_ram[3195] = 46;
    exp_48_ram[3196] = 44;
    exp_48_ram[3197] = 4;
    exp_48_ram[3198] = 23;
    exp_48_ram[3199] = 133;
    exp_48_ram[3200] = 208;
    exp_48_ram[3201] = 23;
    exp_48_ram[3202] = 133;
    exp_48_ram[3203] = 208;
    exp_48_ram[3204] = 23;
    exp_48_ram[3205] = 133;
    exp_48_ram[3206] = 208;
    exp_48_ram[3207] = 23;
    exp_48_ram[3208] = 133;
    exp_48_ram[3209] = 208;
    exp_48_ram[3210] = 23;
    exp_48_ram[3211] = 133;
    exp_48_ram[3212] = 208;
    exp_48_ram[3213] = 23;
    exp_48_ram[3214] = 133;
    exp_48_ram[3215] = 208;
    exp_48_ram[3216] = 23;
    exp_48_ram[3217] = 133;
    exp_48_ram[3218] = 208;
    exp_48_ram[3219] = 208;
    exp_48_ram[3220] = 7;
    exp_48_ram[3221] = 7;
    exp_48_ram[3222] = 71;
    exp_48_ram[3223] = 135;
    exp_48_ram[3224] = 7;
    exp_48_ram[3225] = 106;
    exp_48_ram[3226] = 151;
    exp_48_ram[3227] = 71;
    exp_48_ram[3228] = 135;
    exp_48_ram[3229] = 7;
    exp_48_ram[3230] = 167;
    exp_48_ram[3231] = 128;
    exp_48_ram[3232] = 240;
    exp_48_ram[3233] = 0;
    exp_48_ram[3234] = 240;
    exp_48_ram[3235] = 0;
    exp_48_ram[3236] = 240;
    exp_48_ram[3237] = 0;
    exp_48_ram[3238] = 240;
    exp_48_ram[3239] = 0;
    exp_48_ram[3240] = 0;
    exp_48_ram[3241] = 0;
    exp_48_ram[3242] = 240;
    exp_48_ram[3243] = 0;
    exp_48_ram[3244] = 240;
    exp_48_ram[3245] = 1;
    exp_48_ram[3246] = 46;
    exp_48_ram[3247] = 4;
    exp_48_ram[3248] = 7;
    exp_48_ram[3249] = 7;
    exp_48_ram[3250] = 71;
    exp_48_ram[3251] = 135;
    exp_48_ram[3252] = 7;
    exp_48_ram[3253] = 103;
    exp_48_ram[3254] = 247;
    exp_48_ram[3255] = 133;
    exp_48_ram[3256] = 36;
    exp_48_ram[3257] = 1;
    exp_48_ram[3258] = 128;
    exp_48_ram[3259] = 1;
    exp_48_ram[3260] = 46;
    exp_48_ram[3261] = 44;
    exp_48_ram[3262] = 42;
    exp_48_ram[3263] = 4;
    exp_48_ram[3264] = 46;
    exp_48_ram[3265] = 44;
    exp_48_ram[3266] = 42;
    exp_48_ram[3267] = 40;
    exp_48_ram[3268] = 38;
    exp_48_ram[3269] = 6;
    exp_48_ram[3270] = 135;
    exp_48_ram[3271] = 5;
    exp_48_ram[3272] = 135;
    exp_48_ram[3273] = 5;
    exp_48_ram[3274] = 7;
    exp_48_ram[3275] = 4;
    exp_48_ram[3276] = 71;
    exp_48_ram[3277] = 135;
    exp_48_ram[3278] = 247;
    exp_48_ram[3279] = 39;
    exp_48_ram[3280] = 141;
    exp_48_ram[3281] = 71;
    exp_48_ram[3282] = 135;
    exp_48_ram[3283] = 247;
    exp_48_ram[3284] = 39;
    exp_48_ram[3285] = 142;
    exp_48_ram[3286] = 71;
    exp_48_ram[3287] = 135;
    exp_48_ram[3288] = 247;
    exp_48_ram[3289] = 39;
    exp_48_ram[3290] = 142;
    exp_48_ram[3291] = 39;
    exp_48_ram[3292] = 135;
    exp_48_ram[3293] = 199;
    exp_48_ram[3294] = 135;
    exp_48_ram[3295] = 247;
    exp_48_ram[3296] = 39;
    exp_48_ram[3297] = 140;
    exp_48_ram[3298] = 39;
    exp_48_ram[3299] = 135;
    exp_48_ram[3300] = 199;
    exp_48_ram[3301] = 135;
    exp_48_ram[3302] = 247;
    exp_48_ram[3303] = 39;
    exp_48_ram[3304] = 141;
    exp_48_ram[3305] = 71;
    exp_48_ram[3306] = 135;
    exp_48_ram[3307] = 247;
    exp_48_ram[3308] = 39;
    exp_48_ram[3309] = 139;
    exp_48_ram[3310] = 71;
    exp_48_ram[3311] = 135;
    exp_48_ram[3312] = 247;
    exp_48_ram[3313] = 39;
    exp_48_ram[3314] = 139;
    exp_48_ram[3315] = 71;
    exp_48_ram[3316] = 135;
    exp_48_ram[3317] = 247;
    exp_48_ram[3318] = 39;
    exp_48_ram[3319] = 140;
    exp_48_ram[3320] = 7;
    exp_48_ram[3321] = 0;
    exp_48_ram[3322] = 71;
    exp_48_ram[3323] = 39;
    exp_48_ram[3324] = 7;
    exp_48_ram[3325] = 199;
    exp_48_ram[3326] = 135;
    exp_48_ram[3327] = 7;
    exp_48_ram[3328] = 71;
    exp_48_ram[3329] = 39;
    exp_48_ram[3330] = 7;
    exp_48_ram[3331] = 199;
    exp_48_ram[3332] = 135;
    exp_48_ram[3333] = 6;
    exp_48_ram[3334] = 71;
    exp_48_ram[3335] = 39;
    exp_48_ram[3336] = 7;
    exp_48_ram[3337] = 199;
    exp_48_ram[3338] = 135;
    exp_48_ram[3339] = 6;
    exp_48_ram[3340] = 71;
    exp_48_ram[3341] = 39;
    exp_48_ram[3342] = 7;
    exp_48_ram[3343] = 199;
    exp_48_ram[3344] = 135;
    exp_48_ram[3345] = 5;
    exp_48_ram[3346] = 71;
    exp_48_ram[3347] = 133;
    exp_48_ram[3348] = 240;
    exp_48_ram[3349] = 7;
    exp_48_ram[3350] = 135;
    exp_48_ram[3351] = 39;
    exp_48_ram[3352] = 135;
    exp_48_ram[3353] = 71;
    exp_48_ram[3354] = 141;
    exp_48_ram[3355] = 71;
    exp_48_ram[3356] = 133;
    exp_48_ram[3357] = 240;
    exp_48_ram[3358] = 7;
    exp_48_ram[3359] = 135;
    exp_48_ram[3360] = 39;
    exp_48_ram[3361] = 135;
    exp_48_ram[3362] = 71;
    exp_48_ram[3363] = 135;
    exp_48_ram[3364] = 71;
    exp_48_ram[3365] = 133;
    exp_48_ram[3366] = 240;
    exp_48_ram[3367] = 7;
    exp_48_ram[3368] = 135;
    exp_48_ram[3369] = 39;
    exp_48_ram[3370] = 135;
    exp_48_ram[3371] = 71;
    exp_48_ram[3372] = 138;
    exp_48_ram[3373] = 71;
    exp_48_ram[3374] = 39;
    exp_48_ram[3375] = 7;
    exp_48_ram[3376] = 71;
    exp_48_ram[3377] = 128;
    exp_48_ram[3378] = 68;
    exp_48_ram[3379] = 71;
    exp_48_ram[3380] = 133;
    exp_48_ram[3381] = 240;
    exp_48_ram[3382] = 7;
    exp_48_ram[3383] = 135;
    exp_48_ram[3384] = 39;
    exp_48_ram[3385] = 135;
    exp_48_ram[3386] = 132;
    exp_48_ram[3387] = 68;
    exp_48_ram[3388] = 71;
    exp_48_ram[3389] = 133;
    exp_48_ram[3390] = 240;
    exp_48_ram[3391] = 7;
    exp_48_ram[3392] = 135;
    exp_48_ram[3393] = 39;
    exp_48_ram[3394] = 135;
    exp_48_ram[3395] = 142;
    exp_48_ram[3396] = 68;
    exp_48_ram[3397] = 71;
    exp_48_ram[3398] = 133;
    exp_48_ram[3399] = 240;
    exp_48_ram[3400] = 7;
    exp_48_ram[3401] = 135;
    exp_48_ram[3402] = 39;
    exp_48_ram[3403] = 135;
    exp_48_ram[3404] = 129;
    exp_48_ram[3405] = 71;
    exp_48_ram[3406] = 135;
    exp_48_ram[3407] = 7;
    exp_48_ram[3408] = 71;
    exp_48_ram[3409] = 7;
    exp_48_ram[3410] = 240;
    exp_48_ram[3411] = 0;
    exp_48_ram[3412] = 0;
    exp_48_ram[3413] = 32;
    exp_48_ram[3414] = 36;
    exp_48_ram[3415] = 36;
    exp_48_ram[3416] = 1;
    exp_48_ram[3417] = 128;
    exp_48_ram[3418] = 1;
    exp_48_ram[3419] = 38;
    exp_48_ram[3420] = 36;
    exp_48_ram[3421] = 4;
    exp_48_ram[3422] = 46;
    exp_48_ram[3423] = 135;
    exp_48_ram[3424] = 13;
    exp_48_ram[3425] = 39;
    exp_48_ram[3426] = 199;
    exp_48_ram[3427] = 39;
    exp_48_ram[3428] = 199;
    exp_48_ram[3429] = 22;
    exp_48_ram[3430] = 39;
    exp_48_ram[3431] = 199;
    exp_48_ram[3432] = 135;
    exp_48_ram[3433] = 247;
    exp_48_ram[3434] = 133;
    exp_48_ram[3435] = 240;
    exp_48_ram[3436] = 7;
    exp_48_ram[3437] = 135;
    exp_48_ram[3438] = 39;
    exp_48_ram[3439] = 141;
    exp_48_ram[3440] = 39;
    exp_48_ram[3441] = 199;
    exp_48_ram[3442] = 39;
    exp_48_ram[3443] = 199;
    exp_48_ram[3444] = 22;
    exp_48_ram[3445] = 39;
    exp_48_ram[3446] = 199;
    exp_48_ram[3447] = 135;
    exp_48_ram[3448] = 247;
    exp_48_ram[3449] = 133;
    exp_48_ram[3450] = 240;
    exp_48_ram[3451] = 7;
    exp_48_ram[3452] = 135;
    exp_48_ram[3453] = 39;
    exp_48_ram[3454] = 142;
    exp_48_ram[3455] = 39;
    exp_48_ram[3456] = 199;
    exp_48_ram[3457] = 135;
    exp_48_ram[3458] = 247;
    exp_48_ram[3459] = 133;
    exp_48_ram[3460] = 240;
    exp_48_ram[3461] = 7;
    exp_48_ram[3462] = 135;
    exp_48_ram[3463] = 39;
    exp_48_ram[3464] = 142;
    exp_48_ram[3465] = 71;
    exp_48_ram[3466] = 135;
    exp_48_ram[3467] = 7;
    exp_48_ram[3468] = 39;
    exp_48_ram[3469] = 199;
    exp_48_ram[3470] = 71;
    exp_48_ram[3471] = 7;
    exp_48_ram[3472] = 247;
    exp_48_ram[3473] = 39;
    exp_48_ram[3474] = 199;
    exp_48_ram[3475] = 7;
    exp_48_ram[3476] = 247;
    exp_48_ram[3477] = 133;
    exp_48_ram[3478] = 240;
    exp_48_ram[3479] = 7;
    exp_48_ram[3480] = 135;
    exp_48_ram[3481] = 39;
    exp_48_ram[3482] = 135;
    exp_48_ram[3483] = 199;
    exp_48_ram[3484] = 39;
    exp_48_ram[3485] = 199;
    exp_48_ram[3486] = 7;
    exp_48_ram[3487] = 247;
    exp_48_ram[3488] = 39;
    exp_48_ram[3489] = 199;
    exp_48_ram[3490] = 7;
    exp_48_ram[3491] = 247;
    exp_48_ram[3492] = 133;
    exp_48_ram[3493] = 240;
    exp_48_ram[3494] = 7;
    exp_48_ram[3495] = 7;
    exp_48_ram[3496] = 39;
    exp_48_ram[3497] = 199;
    exp_48_ram[3498] = 71;
    exp_48_ram[3499] = 7;
    exp_48_ram[3500] = 247;
    exp_48_ram[3501] = 39;
    exp_48_ram[3502] = 199;
    exp_48_ram[3503] = 7;
    exp_48_ram[3504] = 247;
    exp_48_ram[3505] = 133;
    exp_48_ram[3506] = 240;
    exp_48_ram[3507] = 7;
    exp_48_ram[3508] = 135;
    exp_48_ram[3509] = 39;
    exp_48_ram[3510] = 135;
    exp_48_ram[3511] = 199;
    exp_48_ram[3512] = 39;
    exp_48_ram[3513] = 199;
    exp_48_ram[3514] = 7;
    exp_48_ram[3515] = 247;
    exp_48_ram[3516] = 39;
    exp_48_ram[3517] = 199;
    exp_48_ram[3518] = 7;
    exp_48_ram[3519] = 247;
    exp_48_ram[3520] = 133;
    exp_48_ram[3521] = 240;
    exp_48_ram[3522] = 7;
    exp_48_ram[3523] = 7;
    exp_48_ram[3524] = 39;
    exp_48_ram[3525] = 199;
    exp_48_ram[3526] = 71;
    exp_48_ram[3527] = 7;
    exp_48_ram[3528] = 247;
    exp_48_ram[3529] = 39;
    exp_48_ram[3530] = 199;
    exp_48_ram[3531] = 7;
    exp_48_ram[3532] = 247;
    exp_48_ram[3533] = 133;
    exp_48_ram[3534] = 240;
    exp_48_ram[3535] = 7;
    exp_48_ram[3536] = 135;
    exp_48_ram[3537] = 39;
    exp_48_ram[3538] = 135;
    exp_48_ram[3539] = 199;
    exp_48_ram[3540] = 39;
    exp_48_ram[3541] = 199;
    exp_48_ram[3542] = 7;
    exp_48_ram[3543] = 247;
    exp_48_ram[3544] = 39;
    exp_48_ram[3545] = 199;
    exp_48_ram[3546] = 7;
    exp_48_ram[3547] = 247;
    exp_48_ram[3548] = 133;
    exp_48_ram[3549] = 240;
    exp_48_ram[3550] = 7;
    exp_48_ram[3551] = 7;
    exp_48_ram[3552] = 71;
    exp_48_ram[3553] = 39;
    exp_48_ram[3554] = 7;
    exp_48_ram[3555] = 199;
    exp_48_ram[3556] = 7;
    exp_48_ram[3557] = 39;
    exp_48_ram[3558] = 199;
    exp_48_ram[3559] = 71;
    exp_48_ram[3560] = 7;
    exp_48_ram[3561] = 247;
    exp_48_ram[3562] = 39;
    exp_48_ram[3563] = 199;
    exp_48_ram[3564] = 7;
    exp_48_ram[3565] = 247;
    exp_48_ram[3566] = 133;
    exp_48_ram[3567] = 240;
    exp_48_ram[3568] = 7;
    exp_48_ram[3569] = 135;
    exp_48_ram[3570] = 39;
    exp_48_ram[3571] = 135;
    exp_48_ram[3572] = 199;
    exp_48_ram[3573] = 39;
    exp_48_ram[3574] = 199;
    exp_48_ram[3575] = 7;
    exp_48_ram[3576] = 247;
    exp_48_ram[3577] = 39;
    exp_48_ram[3578] = 199;
    exp_48_ram[3579] = 7;
    exp_48_ram[3580] = 247;
    exp_48_ram[3581] = 133;
    exp_48_ram[3582] = 240;
    exp_48_ram[3583] = 7;
    exp_48_ram[3584] = 7;
    exp_48_ram[3585] = 39;
    exp_48_ram[3586] = 199;
    exp_48_ram[3587] = 71;
    exp_48_ram[3588] = 7;
    exp_48_ram[3589] = 247;
    exp_48_ram[3590] = 39;
    exp_48_ram[3591] = 199;
    exp_48_ram[3592] = 7;
    exp_48_ram[3593] = 247;
    exp_48_ram[3594] = 133;
    exp_48_ram[3595] = 240;
    exp_48_ram[3596] = 7;
    exp_48_ram[3597] = 135;
    exp_48_ram[3598] = 39;
    exp_48_ram[3599] = 135;
    exp_48_ram[3600] = 199;
    exp_48_ram[3601] = 39;
    exp_48_ram[3602] = 199;
    exp_48_ram[3603] = 7;
    exp_48_ram[3604] = 247;
    exp_48_ram[3605] = 39;
    exp_48_ram[3606] = 199;
    exp_48_ram[3607] = 7;
    exp_48_ram[3608] = 247;
    exp_48_ram[3609] = 133;
    exp_48_ram[3610] = 240;
    exp_48_ram[3611] = 7;
    exp_48_ram[3612] = 7;
    exp_48_ram[3613] = 39;
    exp_48_ram[3614] = 199;
    exp_48_ram[3615] = 71;
    exp_48_ram[3616] = 7;
    exp_48_ram[3617] = 247;
    exp_48_ram[3618] = 39;
    exp_48_ram[3619] = 199;
    exp_48_ram[3620] = 7;
    exp_48_ram[3621] = 247;
    exp_48_ram[3622] = 133;
    exp_48_ram[3623] = 240;
    exp_48_ram[3624] = 7;
    exp_48_ram[3625] = 135;
    exp_48_ram[3626] = 39;
    exp_48_ram[3627] = 135;
    exp_48_ram[3628] = 199;
    exp_48_ram[3629] = 39;
    exp_48_ram[3630] = 199;
    exp_48_ram[3631] = 7;
    exp_48_ram[3632] = 247;
    exp_48_ram[3633] = 39;
    exp_48_ram[3634] = 199;
    exp_48_ram[3635] = 7;
    exp_48_ram[3636] = 247;
    exp_48_ram[3637] = 133;
    exp_48_ram[3638] = 240;
    exp_48_ram[3639] = 7;
    exp_48_ram[3640] = 7;
    exp_48_ram[3641] = 71;
    exp_48_ram[3642] = 135;
    exp_48_ram[3643] = 247;
    exp_48_ram[3644] = 133;
    exp_48_ram[3645] = 32;
    exp_48_ram[3646] = 36;
    exp_48_ram[3647] = 1;
    exp_48_ram[3648] = 128;
    exp_48_ram[3649] = 1;
    exp_48_ram[3650] = 46;
    exp_48_ram[3651] = 44;
    exp_48_ram[3652] = 4;
    exp_48_ram[3653] = 208;
    exp_48_ram[3654] = 7;
    exp_48_ram[3655] = 7;
    exp_48_ram[3656] = 71;
    exp_48_ram[3657] = 7;
    exp_48_ram[3658] = 24;
    exp_48_ram[3659] = 71;
    exp_48_ram[3660] = 135;
    exp_48_ram[3661] = 0;
    exp_48_ram[3662] = 71;
    exp_48_ram[3663] = 7;
    exp_48_ram[3664] = 24;
    exp_48_ram[3665] = 71;
    exp_48_ram[3666] = 135;
    exp_48_ram[3667] = 0;
    exp_48_ram[3668] = 71;
    exp_48_ram[3669] = 7;
    exp_48_ram[3670] = 24;
    exp_48_ram[3671] = 71;
    exp_48_ram[3672] = 135;
    exp_48_ram[3673] = 0;
    exp_48_ram[3674] = 71;
    exp_48_ram[3675] = 7;
    exp_48_ram[3676] = 24;
    exp_48_ram[3677] = 71;
    exp_48_ram[3678] = 135;
    exp_48_ram[3679] = 0;
    exp_48_ram[3680] = 71;
    exp_48_ram[3681] = 7;
    exp_48_ram[3682] = 22;
    exp_48_ram[3683] = 71;
    exp_48_ram[3684] = 135;
    exp_48_ram[3685] = 133;
    exp_48_ram[3686] = 32;
    exp_48_ram[3687] = 36;
    exp_48_ram[3688] = 1;
    exp_48_ram[3689] = 128;
    exp_48_ram[3690] = 1;
    exp_48_ram[3691] = 46;
    exp_48_ram[3692] = 44;
    exp_48_ram[3693] = 4;
    exp_48_ram[3694] = 208;
    exp_48_ram[3695] = 7;
    exp_48_ram[3696] = 7;
    exp_48_ram[3697] = 71;
    exp_48_ram[3698] = 133;
    exp_48_ram[3699] = 208;
    exp_48_ram[3700] = 7;
    exp_48_ram[3701] = 7;
    exp_48_ram[3702] = 24;
    exp_48_ram[3703] = 71;
    exp_48_ram[3704] = 135;
    exp_48_ram[3705] = 0;
    exp_48_ram[3706] = 71;
    exp_48_ram[3707] = 133;
    exp_48_ram[3708] = 208;
    exp_48_ram[3709] = 7;
    exp_48_ram[3710] = 7;
    exp_48_ram[3711] = 24;
    exp_48_ram[3712] = 71;
    exp_48_ram[3713] = 135;
    exp_48_ram[3714] = 0;
    exp_48_ram[3715] = 71;
    exp_48_ram[3716] = 133;
    exp_48_ram[3717] = 208;
    exp_48_ram[3718] = 7;
    exp_48_ram[3719] = 7;
    exp_48_ram[3720] = 28;
    exp_48_ram[3721] = 71;
    exp_48_ram[3722] = 135;
    exp_48_ram[3723] = 133;
    exp_48_ram[3724] = 32;
    exp_48_ram[3725] = 36;
    exp_48_ram[3726] = 1;
    exp_48_ram[3727] = 128;
    exp_48_ram[3728] = 1;
    exp_48_ram[3729] = 46;
    exp_48_ram[3730] = 44;
    exp_48_ram[3731] = 4;
    exp_48_ram[3732] = 208;
    exp_48_ram[3733] = 7;
    exp_48_ram[3734] = 7;
    exp_48_ram[3735] = 71;
    exp_48_ram[3736] = 133;
    exp_48_ram[3737] = 208;
    exp_48_ram[3738] = 7;
    exp_48_ram[3739] = 130;
    exp_48_ram[3740] = 71;
    exp_48_ram[3741] = 133;
    exp_48_ram[3742] = 208;
    exp_48_ram[3743] = 7;
    exp_48_ram[3744] = 247;
    exp_48_ram[3745] = 133;
    exp_48_ram[3746] = 32;
    exp_48_ram[3747] = 36;
    exp_48_ram[3748] = 1;
    exp_48_ram[3749] = 128;
    exp_48_ram[3750] = 1;
    exp_48_ram[3751] = 46;
    exp_48_ram[3752] = 44;
    exp_48_ram[3753] = 4;
    exp_48_ram[3754] = 71;
    exp_48_ram[3755] = 165;
    exp_48_ram[3756] = 71;
    exp_48_ram[3757] = 166;
    exp_48_ram[3758] = 71;
    exp_48_ram[3759] = 165;
    exp_48_ram[3760] = 71;
    exp_48_ram[3761] = 163;
    exp_48_ram[3762] = 71;
    exp_48_ram[3763] = 206;
    exp_48_ram[3764] = 71;
    exp_48_ram[3765] = 200;
    exp_48_ram[3766] = 71;
    exp_48_ram[3767] = 200;
    exp_48_ram[3768] = 71;
    exp_48_ram[3769] = 199;
    exp_48_ram[3770] = 71;
    exp_48_ram[3771] = 71;
    exp_48_ram[3772] = 70;
    exp_48_ram[3773] = 198;
    exp_48_ram[3774] = 36;
    exp_48_ram[3775] = 34;
    exp_48_ram[3776] = 32;
    exp_48_ram[3777] = 7;
    exp_48_ram[3778] = 7;
    exp_48_ram[3779] = 6;
    exp_48_ram[3780] = 69;
    exp_48_ram[3781] = 5;
    exp_48_ram[3782] = 240;
    exp_48_ram[3783] = 23;
    exp_48_ram[3784] = 133;
    exp_48_ram[3785] = 208;
    exp_48_ram[3786] = 71;
    exp_48_ram[3787] = 199;
    exp_48_ram[3788] = 133;
    exp_48_ram[3789] = 208;
    exp_48_ram[3790] = 71;
    exp_48_ram[3791] = 199;
    exp_48_ram[3792] = 133;
    exp_48_ram[3793] = 208;
    exp_48_ram[3794] = 71;
    exp_48_ram[3795] = 199;
    exp_48_ram[3796] = 133;
    exp_48_ram[3797] = 208;
    exp_48_ram[3798] = 23;
    exp_48_ram[3799] = 133;
    exp_48_ram[3800] = 208;
    exp_48_ram[3801] = 0;
    exp_48_ram[3802] = 32;
    exp_48_ram[3803] = 36;
    exp_48_ram[3804] = 1;
    exp_48_ram[3805] = 128;
    exp_48_ram[3806] = 1;
    exp_48_ram[3807] = 46;
    exp_48_ram[3808] = 44;
    exp_48_ram[3809] = 4;
    exp_48_ram[3810] = 71;
    exp_48_ram[3811] = 71;
    exp_48_ram[3812] = 7;
    exp_48_ram[3813] = 168;
    exp_48_ram[3814] = 71;
    exp_48_ram[3815] = 71;
    exp_48_ram[3816] = 7;
    exp_48_ram[3817] = 170;
    exp_48_ram[3818] = 71;
    exp_48_ram[3819] = 71;
    exp_48_ram[3820] = 7;
    exp_48_ram[3821] = 172;
    exp_48_ram[3822] = 71;
    exp_48_ram[3823] = 71;
    exp_48_ram[3824] = 7;
    exp_48_ram[3825] = 174;
    exp_48_ram[3826] = 71;
    exp_48_ram[3827] = 7;
    exp_48_ram[3828] = 128;
    exp_48_ram[3829] = 71;
    exp_48_ram[3830] = 7;
    exp_48_ram[3831] = 128;
    exp_48_ram[3832] = 71;
    exp_48_ram[3833] = 7;
    exp_48_ram[3834] = 129;
    exp_48_ram[3835] = 71;
    exp_48_ram[3836] = 7;
    exp_48_ram[3837] = 129;
    exp_48_ram[3838] = 71;
    exp_48_ram[3839] = 7;
    exp_48_ram[3840] = 130;
    exp_48_ram[3841] = 71;
    exp_48_ram[3842] = 7;
    exp_48_ram[3843] = 130;
    exp_48_ram[3844] = 240;
    exp_48_ram[3845] = 23;
    exp_48_ram[3846] = 133;
    exp_48_ram[3847] = 208;
    exp_48_ram[3848] = 23;
    exp_48_ram[3849] = 133;
    exp_48_ram[3850] = 208;
    exp_48_ram[3851] = 23;
    exp_48_ram[3852] = 133;
    exp_48_ram[3853] = 208;
    exp_48_ram[3854] = 23;
    exp_48_ram[3855] = 133;
    exp_48_ram[3856] = 208;
    exp_48_ram[3857] = 23;
    exp_48_ram[3858] = 133;
    exp_48_ram[3859] = 208;
    exp_48_ram[3860] = 23;
    exp_48_ram[3861] = 133;
    exp_48_ram[3862] = 208;
    exp_48_ram[3863] = 23;
    exp_48_ram[3864] = 133;
    exp_48_ram[3865] = 208;
    exp_48_ram[3866] = 38;
    exp_48_ram[3867] = 208;
    exp_48_ram[3868] = 7;
    exp_48_ram[3869] = 5;
    exp_48_ram[3870] = 71;
    exp_48_ram[3871] = 133;
    exp_48_ram[3872] = 208;
    exp_48_ram[3873] = 7;
    exp_48_ram[3874] = 142;
    exp_48_ram[3875] = 39;
    exp_48_ram[3876] = 156;
    exp_48_ram[3877] = 71;
    exp_48_ram[3878] = 135;
    exp_48_ram[3879] = 199;
    exp_48_ram[3880] = 135;
    exp_48_ram[3881] = 133;
    exp_48_ram[3882] = 208;
    exp_48_ram[3883] = 71;
    exp_48_ram[3884] = 135;
    exp_48_ram[3885] = 199;
    exp_48_ram[3886] = 135;
    exp_48_ram[3887] = 133;
    exp_48_ram[3888] = 208;
    exp_48_ram[3889] = 71;
    exp_48_ram[3890] = 135;
    exp_48_ram[3891] = 199;
    exp_48_ram[3892] = 135;
    exp_48_ram[3893] = 133;
    exp_48_ram[3894] = 208;
    exp_48_ram[3895] = 23;
    exp_48_ram[3896] = 133;
    exp_48_ram[3897] = 208;
    exp_48_ram[3898] = 71;
    exp_48_ram[3899] = 133;
    exp_48_ram[3900] = 208;
    exp_48_ram[3901] = 7;
    exp_48_ram[3902] = 247;
    exp_48_ram[3903] = 133;
    exp_48_ram[3904] = 71;
    exp_48_ram[3905] = 133;
    exp_48_ram[3906] = 240;
    exp_48_ram[3907] = 7;
    exp_48_ram[3908] = 133;
    exp_48_ram[3909] = 192;
    exp_48_ram[3910] = 39;
    exp_48_ram[3911] = 7;
    exp_48_ram[3912] = 26;
    exp_48_ram[3913] = 38;
    exp_48_ram[3914] = 5;
    exp_48_ram[3915] = 192;
    exp_48_ram[3916] = 240;
    exp_48_ram[3917] = 39;
    exp_48_ram[3918] = 135;
    exp_48_ram[3919] = 38;
    exp_48_ram[3920] = 240;
    exp_48_ram[3921] = 71;
    exp_48_ram[3922] = 135;
    exp_48_ram[3923] = 7;
    exp_48_ram[3924] = 238;
    exp_48_ram[3925] = 71;
    exp_48_ram[3926] = 7;
    exp_48_ram[3927] = 22;
    exp_48_ram[3928] = 23;
    exp_48_ram[3929] = 133;
    exp_48_ram[3930] = 208;
    exp_48_ram[3931] = 240;
    exp_48_ram[3932] = 7;
    exp_48_ram[3933] = 71;
    exp_48_ram[3934] = 168;
    exp_48_ram[3935] = 240;
    exp_48_ram[3936] = 7;
    exp_48_ram[3937] = 71;
    exp_48_ram[3938] = 170;
    exp_48_ram[3939] = 240;
    exp_48_ram[3940] = 7;
    exp_48_ram[3941] = 71;
    exp_48_ram[3942] = 172;
    exp_48_ram[3943] = 240;
    exp_48_ram[3944] = 38;
    exp_48_ram[3945] = 240;
    exp_48_ram[3946] = 71;
    exp_48_ram[3947] = 7;
    exp_48_ram[3948] = 22;
    exp_48_ram[3949] = 23;
    exp_48_ram[3950] = 133;
    exp_48_ram[3951] = 208;
    exp_48_ram[3952] = 240;
    exp_48_ram[3953] = 7;
    exp_48_ram[3954] = 71;
    exp_48_ram[3955] = 174;
    exp_48_ram[3956] = 240;
    exp_48_ram[3957] = 38;
    exp_48_ram[3958] = 240;
    exp_48_ram[3959] = 71;
    exp_48_ram[3960] = 7;
    exp_48_ram[3961] = 28;
    exp_48_ram[3962] = 23;
    exp_48_ram[3963] = 133;
    exp_48_ram[3964] = 192;
    exp_48_ram[3965] = 240;
    exp_48_ram[3966] = 7;
    exp_48_ram[3967] = 135;
    exp_48_ram[3968] = 71;
    exp_48_ram[3969] = 128;
    exp_48_ram[3970] = 240;
    exp_48_ram[3971] = 7;
    exp_48_ram[3972] = 135;
    exp_48_ram[3973] = 71;
    exp_48_ram[3974] = 128;
    exp_48_ram[3975] = 240;
    exp_48_ram[3976] = 7;
    exp_48_ram[3977] = 135;
    exp_48_ram[3978] = 71;
    exp_48_ram[3979] = 129;
    exp_48_ram[3980] = 240;
    exp_48_ram[3981] = 38;
    exp_48_ram[3982] = 240;
    exp_48_ram[3983] = 71;
    exp_48_ram[3984] = 7;
    exp_48_ram[3985] = 20;
    exp_48_ram[3986] = 23;
    exp_48_ram[3987] = 133;
    exp_48_ram[3988] = 192;
    exp_48_ram[3989] = 240;
    exp_48_ram[3990] = 7;
    exp_48_ram[3991] = 135;
    exp_48_ram[3992] = 71;
    exp_48_ram[3993] = 129;
    exp_48_ram[3994] = 240;
    exp_48_ram[3995] = 7;
    exp_48_ram[3996] = 135;
    exp_48_ram[3997] = 71;
    exp_48_ram[3998] = 130;
    exp_48_ram[3999] = 240;
    exp_48_ram[4000] = 7;
    exp_48_ram[4001] = 135;
    exp_48_ram[4002] = 71;
    exp_48_ram[4003] = 130;
    exp_48_ram[4004] = 240;
    exp_48_ram[4005] = 38;
    exp_48_ram[4006] = 240;
    exp_48_ram[4007] = 7;
    exp_48_ram[4008] = 135;
    exp_48_ram[4009] = 69;
    exp_48_ram[4010] = 1;
    exp_48_ram[4011] = 101;
    exp_48_ram[4012] = 76;
    exp_48_ram[4013] = 214;
    exp_48_ram[4014] = 5;
    exp_48_ram[4015] = 133;
    exp_48_ram[4016] = 1;
    exp_48_ram[4017] = 128;
    exp_48_ram[4018] = 92;
    exp_48_ram[4019] = 5;
    exp_48_ram[4020] = 133;
    exp_48_ram[4021] = 240;
    exp_48_ram[4022] = 240;
    exp_48_ram[4023] = 0;
    exp_48_ram[4024] = 0;
    exp_48_ram[4025] = 0;
    exp_48_ram[4026] = 0;
    exp_48_ram[4027] = 50;
    exp_48_ram[4028] = 50;
    exp_48_ram[4029] = 50;
    exp_48_ram[4030] = 50;
    exp_48_ram[4031] = 50;
    exp_48_ram[4032] = 50;
    exp_48_ram[4033] = 75;
    exp_48_ram[4034] = 71;
    exp_48_ram[4035] = 90;
    exp_48_ram[4036] = 87;
    exp_48_ram[4037] = 85;
    exp_48_ram[4038] = 73;
    exp_48_ram[4039] = 74;
    exp_48_ram[4040] = 74;
    exp_48_ram[4041] = 73;
    exp_48_ram[4042] = 66;
    exp_48_ram[4043] = 84;
    exp_48_ram[4044] = 71;
    exp_48_ram[4045] = 89;
    exp_48_ram[4046] = 69;
    exp_48_ram[4047] = 68;
    exp_48_ram[4048] = 76;
    exp_48_ram[4049] = 84;
    exp_48_ram[4050] = 78;
    exp_48_ram[4051] = 87;
    exp_48_ram[4052] = 77;
    exp_48_ram[4053] = 79;
    exp_48_ram[4054] = 83;
    exp_48_ram[4055] = 90;
    exp_48_ram[4056] = 81;
    exp_48_ram[4057] = 72;
    exp_48_ram[4058] = 70;
    exp_48_ram[4059] = 68;
    exp_48_ram[4060] = 66;
    exp_48_ram[4061] = 90;
    exp_48_ram[4062] = 73;
    exp_48_ram[4063] = 80;
    exp_48_ram[4064] = 72;
    exp_48_ram[4065] = 87;
    exp_48_ram[4066] = 79;
    exp_48_ram[4067] = 75;
    exp_48_ram[4068] = 74;
    exp_48_ram[4069] = 76;
    exp_48_ram[4070] = 66;
    exp_48_ram[4071] = 82;
    exp_48_ram[4072] = 78;
    exp_48_ram[4073] = 73;
    exp_48_ram[4074] = 68;
    exp_48_ram[4075] = 82;
    exp_48_ram[4076] = 83;
    exp_48_ram[4077] = 88;
    exp_48_ram[4078] = 75;
    exp_48_ram[4079] = 66;
    exp_48_ram[4080] = 87;
    exp_48_ram[4081] = 84;
    exp_48_ram[4082] = 86;
    exp_48_ram[4083] = 65;
    exp_48_ram[4084] = 68;
    exp_48_ram[4085] = 87;
    exp_48_ram[4086] = 75;
    exp_48_ram[4087] = 66;
    exp_48_ram[4088] = 76;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_46) begin
      exp_48_ram[exp_42] <= exp_44;
    end
  end
  assign exp_48 = exp_48_ram[exp_43];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_74) begin
        exp_48_ram[exp_70] <= exp_72;
    end
  end
  assign exp_76 = exp_48_ram[exp_71];
  assign exp_75 = exp_98;
  assign exp_98 = 1;
  assign exp_71 = exp_97;
  assign exp_97 = exp_16[31:2];
  assign exp_74 = exp_92;
  assign exp_70 = exp_91;
  assign exp_72 = exp_91;
  assign exp_47 = exp_133;
  assign exp_133 = 1;
  assign exp_43 = exp_132;
  assign exp_132 = exp_18[31:2];
  assign exp_46 = exp_114;
  assign exp_114 = exp_112 & exp_113;
  assign exp_112 = exp_22 & exp_23;
  assign exp_113 = exp_24[1:1];
  assign exp_42 = exp_110;
  assign exp_110 = exp_18[31:2];
  assign exp_44 = exp_111;
  assign exp_111 = exp_19[15:8];

  //Create RAM
  reg [7:0] exp_41_ram [5119:0];


  //Initialise RAM contents
  initial
  begin
    exp_41_ram[0] = 147;
    exp_41_ram[1] = 19;
    exp_41_ram[2] = 147;
    exp_41_ram[3] = 19;
    exp_41_ram[4] = 147;
    exp_41_ram[5] = 19;
    exp_41_ram[6] = 147;
    exp_41_ram[7] = 19;
    exp_41_ram[8] = 147;
    exp_41_ram[9] = 19;
    exp_41_ram[10] = 147;
    exp_41_ram[11] = 19;
    exp_41_ram[12] = 147;
    exp_41_ram[13] = 19;
    exp_41_ram[14] = 147;
    exp_41_ram[15] = 19;
    exp_41_ram[16] = 147;
    exp_41_ram[17] = 19;
    exp_41_ram[18] = 147;
    exp_41_ram[19] = 19;
    exp_41_ram[20] = 147;
    exp_41_ram[21] = 19;
    exp_41_ram[22] = 147;
    exp_41_ram[23] = 19;
    exp_41_ram[24] = 147;
    exp_41_ram[25] = 19;
    exp_41_ram[26] = 147;
    exp_41_ram[27] = 19;
    exp_41_ram[28] = 147;
    exp_41_ram[29] = 19;
    exp_41_ram[30] = 147;
    exp_41_ram[31] = 55;
    exp_41_ram[32] = 19;
    exp_41_ram[33] = 239;
    exp_41_ram[34] = 111;
    exp_41_ram[35] = 147;
    exp_41_ram[36] = 147;
    exp_41_ram[37] = 19;
    exp_41_ram[38] = 19;
    exp_41_ram[39] = 19;
    exp_41_ram[40] = 99;
    exp_41_ram[41] = 183;
    exp_41_ram[42] = 147;
    exp_41_ram[43] = 99;
    exp_41_ram[44] = 55;
    exp_41_ram[45] = 99;
    exp_41_ram[46] = 19;
    exp_41_ram[47] = 51;
    exp_41_ram[48] = 19;
    exp_41_ram[49] = 51;
    exp_41_ram[50] = 179;
    exp_41_ram[51] = 131;
    exp_41_ram[52] = 19;
    exp_41_ram[53] = 51;
    exp_41_ram[54] = 179;
    exp_41_ram[55] = 99;
    exp_41_ram[56] = 179;
    exp_41_ram[57] = 51;
    exp_41_ram[58] = 51;
    exp_41_ram[59] = 179;
    exp_41_ram[60] = 51;
    exp_41_ram[61] = 147;
    exp_41_ram[62] = 179;
    exp_41_ram[63] = 19;
    exp_41_ram[64] = 19;
    exp_41_ram[65] = 147;
    exp_41_ram[66] = 51;
    exp_41_ram[67] = 19;
    exp_41_ram[68] = 179;
    exp_41_ram[69] = 19;
    exp_41_ram[70] = 179;
    exp_41_ram[71] = 99;
    exp_41_ram[72] = 179;
    exp_41_ram[73] = 19;
    exp_41_ram[74] = 99;
    exp_41_ram[75] = 99;
    exp_41_ram[76] = 19;
    exp_41_ram[77] = 179;
    exp_41_ram[78] = 179;
    exp_41_ram[79] = 51;
    exp_41_ram[80] = 19;
    exp_41_ram[81] = 19;
    exp_41_ram[82] = 179;
    exp_41_ram[83] = 19;
    exp_41_ram[84] = 51;
    exp_41_ram[85] = 179;
    exp_41_ram[86] = 19;
    exp_41_ram[87] = 99;
    exp_41_ram[88] = 51;
    exp_41_ram[89] = 19;
    exp_41_ram[90] = 99;
    exp_41_ram[91] = 99;
    exp_41_ram[92] = 19;
    exp_41_ram[93] = 19;
    exp_41_ram[94] = 51;
    exp_41_ram[95] = 147;
    exp_41_ram[96] = 111;
    exp_41_ram[97] = 55;
    exp_41_ram[98] = 19;
    exp_41_ram[99] = 227;
    exp_41_ram[100] = 19;
    exp_41_ram[101] = 111;
    exp_41_ram[102] = 99;
    exp_41_ram[103] = 19;
    exp_41_ram[104] = 51;
    exp_41_ram[105] = 55;
    exp_41_ram[106] = 99;
    exp_41_ram[107] = 19;
    exp_41_ram[108] = 99;
    exp_41_ram[109] = 19;
    exp_41_ram[110] = 51;
    exp_41_ram[111] = 179;
    exp_41_ram[112] = 3;
    exp_41_ram[113] = 19;
    exp_41_ram[114] = 51;
    exp_41_ram[115] = 179;
    exp_41_ram[116] = 99;
    exp_41_ram[117] = 179;
    exp_41_ram[118] = 147;
    exp_41_ram[119] = 147;
    exp_41_ram[120] = 19;
    exp_41_ram[121] = 19;
    exp_41_ram[122] = 19;
    exp_41_ram[123] = 179;
    exp_41_ram[124] = 179;
    exp_41_ram[125] = 147;
    exp_41_ram[126] = 51;
    exp_41_ram[127] = 51;
    exp_41_ram[128] = 19;
    exp_41_ram[129] = 99;
    exp_41_ram[130] = 51;
    exp_41_ram[131] = 19;
    exp_41_ram[132] = 99;
    exp_41_ram[133] = 99;
    exp_41_ram[134] = 19;
    exp_41_ram[135] = 51;
    exp_41_ram[136] = 51;
    exp_41_ram[137] = 179;
    exp_41_ram[138] = 19;
    exp_41_ram[139] = 19;
    exp_41_ram[140] = 51;
    exp_41_ram[141] = 147;
    exp_41_ram[142] = 51;
    exp_41_ram[143] = 179;
    exp_41_ram[144] = 19;
    exp_41_ram[145] = 99;
    exp_41_ram[146] = 51;
    exp_41_ram[147] = 19;
    exp_41_ram[148] = 99;
    exp_41_ram[149] = 99;
    exp_41_ram[150] = 19;
    exp_41_ram[151] = 19;
    exp_41_ram[152] = 51;
    exp_41_ram[153] = 103;
    exp_41_ram[154] = 55;
    exp_41_ram[155] = 19;
    exp_41_ram[156] = 227;
    exp_41_ram[157] = 19;
    exp_41_ram[158] = 111;
    exp_41_ram[159] = 51;
    exp_41_ram[160] = 51;
    exp_41_ram[161] = 51;
    exp_41_ram[162] = 179;
    exp_41_ram[163] = 51;
    exp_41_ram[164] = 147;
    exp_41_ram[165] = 51;
    exp_41_ram[166] = 51;
    exp_41_ram[167] = 147;
    exp_41_ram[168] = 147;
    exp_41_ram[169] = 147;
    exp_41_ram[170] = 51;
    exp_41_ram[171] = 19;
    exp_41_ram[172] = 51;
    exp_41_ram[173] = 179;
    exp_41_ram[174] = 147;
    exp_41_ram[175] = 99;
    exp_41_ram[176] = 51;
    exp_41_ram[177] = 147;
    exp_41_ram[178] = 99;
    exp_41_ram[179] = 99;
    exp_41_ram[180] = 147;
    exp_41_ram[181] = 51;
    exp_41_ram[182] = 179;
    exp_41_ram[183] = 51;
    exp_41_ram[184] = 19;
    exp_41_ram[185] = 19;
    exp_41_ram[186] = 179;
    exp_41_ram[187] = 19;
    exp_41_ram[188] = 51;
    exp_41_ram[189] = 179;
    exp_41_ram[190] = 19;
    exp_41_ram[191] = 99;
    exp_41_ram[192] = 179;
    exp_41_ram[193] = 19;
    exp_41_ram[194] = 99;
    exp_41_ram[195] = 99;
    exp_41_ram[196] = 19;
    exp_41_ram[197] = 179;
    exp_41_ram[198] = 147;
    exp_41_ram[199] = 179;
    exp_41_ram[200] = 179;
    exp_41_ram[201] = 111;
    exp_41_ram[202] = 99;
    exp_41_ram[203] = 55;
    exp_41_ram[204] = 99;
    exp_41_ram[205] = 19;
    exp_41_ram[206] = 179;
    exp_41_ram[207] = 147;
    exp_41_ram[208] = 55;
    exp_41_ram[209] = 51;
    exp_41_ram[210] = 19;
    exp_41_ram[211] = 51;
    exp_41_ram[212] = 3;
    exp_41_ram[213] = 19;
    exp_41_ram[214] = 51;
    exp_41_ram[215] = 179;
    exp_41_ram[216] = 99;
    exp_41_ram[217] = 19;
    exp_41_ram[218] = 227;
    exp_41_ram[219] = 51;
    exp_41_ram[220] = 19;
    exp_41_ram[221] = 111;
    exp_41_ram[222] = 55;
    exp_41_ram[223] = 147;
    exp_41_ram[224] = 227;
    exp_41_ram[225] = 147;
    exp_41_ram[226] = 111;
    exp_41_ram[227] = 51;
    exp_41_ram[228] = 179;
    exp_41_ram[229] = 51;
    exp_41_ram[230] = 51;
    exp_41_ram[231] = 147;
    exp_41_ram[232] = 179;
    exp_41_ram[233] = 179;
    exp_41_ram[234] = 51;
    exp_41_ram[235] = 51;
    exp_41_ram[236] = 51;
    exp_41_ram[237] = 147;
    exp_41_ram[238] = 147;
    exp_41_ram[239] = 19;
    exp_41_ram[240] = 51;
    exp_41_ram[241] = 147;
    exp_41_ram[242] = 51;
    exp_41_ram[243] = 51;
    exp_41_ram[244] = 19;
    exp_41_ram[245] = 99;
    exp_41_ram[246] = 51;
    exp_41_ram[247] = 19;
    exp_41_ram[248] = 99;
    exp_41_ram[249] = 99;
    exp_41_ram[250] = 19;
    exp_41_ram[251] = 51;
    exp_41_ram[252] = 51;
    exp_41_ram[253] = 179;
    exp_41_ram[254] = 51;
    exp_41_ram[255] = 147;
    exp_41_ram[256] = 51;
    exp_41_ram[257] = 147;
    exp_41_ram[258] = 147;
    exp_41_ram[259] = 179;
    exp_41_ram[260] = 19;
    exp_41_ram[261] = 99;
    exp_41_ram[262] = 179;
    exp_41_ram[263] = 19;
    exp_41_ram[264] = 99;
    exp_41_ram[265] = 99;
    exp_41_ram[266] = 19;
    exp_41_ram[267] = 179;
    exp_41_ram[268] = 19;
    exp_41_ram[269] = 183;
    exp_41_ram[270] = 51;
    exp_41_ram[271] = 147;
    exp_41_ram[272] = 51;
    exp_41_ram[273] = 19;
    exp_41_ram[274] = 179;
    exp_41_ram[275] = 19;
    exp_41_ram[276] = 179;
    exp_41_ram[277] = 51;
    exp_41_ram[278] = 179;
    exp_41_ram[279] = 19;
    exp_41_ram[280] = 51;
    exp_41_ram[281] = 51;
    exp_41_ram[282] = 51;
    exp_41_ram[283] = 51;
    exp_41_ram[284] = 99;
    exp_41_ram[285] = 51;
    exp_41_ram[286] = 147;
    exp_41_ram[287] = 51;
    exp_41_ram[288] = 99;
    exp_41_ram[289] = 227;
    exp_41_ram[290] = 183;
    exp_41_ram[291] = 147;
    exp_41_ram[292] = 51;
    exp_41_ram[293] = 19;
    exp_41_ram[294] = 51;
    exp_41_ram[295] = 179;
    exp_41_ram[296] = 51;
    exp_41_ram[297] = 147;
    exp_41_ram[298] = 227;
    exp_41_ram[299] = 19;
    exp_41_ram[300] = 111;
    exp_41_ram[301] = 147;
    exp_41_ram[302] = 19;
    exp_41_ram[303] = 111;
    exp_41_ram[304] = 55;
    exp_41_ram[305] = 19;
    exp_41_ram[306] = 19;
    exp_41_ram[307] = 179;
    exp_41_ram[308] = 147;
    exp_41_ram[309] = 19;
    exp_41_ram[310] = 19;
    exp_41_ram[311] = 19;
    exp_41_ram[312] = 147;
    exp_41_ram[313] = 147;
    exp_41_ram[314] = 51;
    exp_41_ram[315] = 19;
    exp_41_ram[316] = 147;
    exp_41_ram[317] = 147;
    exp_41_ram[318] = 99;
    exp_41_ram[319] = 179;
    exp_41_ram[320] = 99;
    exp_41_ram[321] = 19;
    exp_41_ram[322] = 103;
    exp_41_ram[323] = 99;
    exp_41_ram[324] = 179;
    exp_41_ram[325] = 227;
    exp_41_ram[326] = 99;
    exp_41_ram[327] = 179;
    exp_41_ram[328] = 147;
    exp_41_ram[329] = 99;
    exp_41_ram[330] = 51;
    exp_41_ram[331] = 99;
    exp_41_ram[332] = 99;
    exp_41_ram[333] = 99;
    exp_41_ram[334] = 99;
    exp_41_ram[335] = 99;
    exp_41_ram[336] = 19;
    exp_41_ram[337] = 103;
    exp_41_ram[338] = 19;
    exp_41_ram[339] = 99;
    exp_41_ram[340] = 19;
    exp_41_ram[341] = 103;
    exp_41_ram[342] = 99;
    exp_41_ram[343] = 227;
    exp_41_ram[344] = 103;
    exp_41_ram[345] = 227;
    exp_41_ram[346] = 99;
    exp_41_ram[347] = 227;
    exp_41_ram[348] = 227;
    exp_41_ram[349] = 19;
    exp_41_ram[350] = 103;
    exp_41_ram[351] = 19;
    exp_41_ram[352] = 103;
    exp_41_ram[353] = 227;
    exp_41_ram[354] = 111;
    exp_41_ram[355] = 227;
    exp_41_ram[356] = 111;
    exp_41_ram[357] = 227;
    exp_41_ram[358] = 227;
    exp_41_ram[359] = 147;
    exp_41_ram[360] = 111;
    exp_41_ram[361] = 19;
    exp_41_ram[362] = 35;
    exp_41_ram[363] = 35;
    exp_41_ram[364] = 19;
    exp_41_ram[365] = 99;
    exp_41_ram[366] = 239;
    exp_41_ram[367] = 19;
    exp_41_ram[368] = 147;
    exp_41_ram[369] = 51;
    exp_41_ram[370] = 99;
    exp_41_ram[371] = 147;
    exp_41_ram[372] = 179;
    exp_41_ram[373] = 19;
    exp_41_ram[374] = 179;
    exp_41_ram[375] = 51;
    exp_41_ram[376] = 131;
    exp_41_ram[377] = 19;
    exp_41_ram[378] = 147;
    exp_41_ram[379] = 3;
    exp_41_ram[380] = 19;
    exp_41_ram[381] = 147;
    exp_41_ram[382] = 179;
    exp_41_ram[383] = 147;
    exp_41_ram[384] = 19;
    exp_41_ram[385] = 103;
    exp_41_ram[386] = 147;
    exp_41_ram[387] = 179;
    exp_41_ram[388] = 19;
    exp_41_ram[389] = 111;
    exp_41_ram[390] = 147;
    exp_41_ram[391] = 19;
    exp_41_ram[392] = 111;
    exp_41_ram[393] = 19;
    exp_41_ram[394] = 35;
    exp_41_ram[395] = 35;
    exp_41_ram[396] = 35;
    exp_41_ram[397] = 35;
    exp_41_ram[398] = 35;
    exp_41_ram[399] = 35;
    exp_41_ram[400] = 179;
    exp_41_ram[401] = 99;
    exp_41_ram[402] = 19;
    exp_41_ram[403] = 19;
    exp_41_ram[404] = 147;
    exp_41_ram[405] = 99;
    exp_41_ram[406] = 19;
    exp_41_ram[407] = 239;
    exp_41_ram[408] = 147;
    exp_41_ram[409] = 19;
    exp_41_ram[410] = 51;
    exp_41_ram[411] = 147;
    exp_41_ram[412] = 99;
    exp_41_ram[413] = 19;
    exp_41_ram[414] = 147;
    exp_41_ram[415] = 99;
    exp_41_ram[416] = 19;
    exp_41_ram[417] = 99;
    exp_41_ram[418] = 147;
    exp_41_ram[419] = 19;
    exp_41_ram[420] = 179;
    exp_41_ram[421] = 179;
    exp_41_ram[422] = 179;
    exp_41_ram[423] = 179;
    exp_41_ram[424] = 179;
    exp_41_ram[425] = 131;
    exp_41_ram[426] = 3;
    exp_41_ram[427] = 147;
    exp_41_ram[428] = 19;
    exp_41_ram[429] = 147;
    exp_41_ram[430] = 51;
    exp_41_ram[431] = 131;
    exp_41_ram[432] = 3;
    exp_41_ram[433] = 131;
    exp_41_ram[434] = 3;
    exp_41_ram[435] = 19;
    exp_41_ram[436] = 147;
    exp_41_ram[437] = 19;
    exp_41_ram[438] = 103;
    exp_41_ram[439] = 239;
    exp_41_ram[440] = 147;
    exp_41_ram[441] = 111;
    exp_41_ram[442] = 147;
    exp_41_ram[443] = 179;
    exp_41_ram[444] = 147;
    exp_41_ram[445] = 111;
    exp_41_ram[446] = 147;
    exp_41_ram[447] = 99;
    exp_41_ram[448] = 19;
    exp_41_ram[449] = 19;
    exp_41_ram[450] = 147;
    exp_41_ram[451] = 239;
    exp_41_ram[452] = 51;
    exp_41_ram[453] = 19;
    exp_41_ram[454] = 179;
    exp_41_ram[455] = 147;
    exp_41_ram[456] = 19;
    exp_41_ram[457] = 51;
    exp_41_ram[458] = 239;
    exp_41_ram[459] = 51;
    exp_41_ram[460] = 19;
    exp_41_ram[461] = 19;
    exp_41_ram[462] = 147;
    exp_41_ram[463] = 147;
    exp_41_ram[464] = 99;
    exp_41_ram[465] = 19;
    exp_41_ram[466] = 99;
    exp_41_ram[467] = 19;
    exp_41_ram[468] = 179;
    exp_41_ram[469] = 19;
    exp_41_ram[470] = 51;
    exp_41_ram[471] = 51;
    exp_41_ram[472] = 179;
    exp_41_ram[473] = 179;
    exp_41_ram[474] = 55;
    exp_41_ram[475] = 19;
    exp_41_ram[476] = 179;
    exp_41_ram[477] = 19;
    exp_41_ram[478] = 99;
    exp_41_ram[479] = 19;
    exp_41_ram[480] = 147;
    exp_41_ram[481] = 99;
    exp_41_ram[482] = 19;
    exp_41_ram[483] = 179;
    exp_41_ram[484] = 179;
    exp_41_ram[485] = 147;
    exp_41_ram[486] = 55;
    exp_41_ram[487] = 51;
    exp_41_ram[488] = 99;
    exp_41_ram[489] = 55;
    exp_41_ram[490] = 19;
    exp_41_ram[491] = 19;
    exp_41_ram[492] = 179;
    exp_41_ram[493] = 51;
    exp_41_ram[494] = 147;
    exp_41_ram[495] = 19;
    exp_41_ram[496] = 179;
    exp_41_ram[497] = 147;
    exp_41_ram[498] = 111;
    exp_41_ram[499] = 147;
    exp_41_ram[500] = 179;
    exp_41_ram[501] = 147;
    exp_41_ram[502] = 111;
    exp_41_ram[503] = 147;
    exp_41_ram[504] = 147;
    exp_41_ram[505] = 19;
    exp_41_ram[506] = 111;
    exp_41_ram[507] = 99;
    exp_41_ram[508] = 147;
    exp_41_ram[509] = 179;
    exp_41_ram[510] = 99;
    exp_41_ram[511] = 19;
    exp_41_ram[512] = 19;
    exp_41_ram[513] = 51;
    exp_41_ram[514] = 147;
    exp_41_ram[515] = 103;
    exp_41_ram[516] = 51;
    exp_41_ram[517] = 51;
    exp_41_ram[518] = 179;
    exp_41_ram[519] = 51;
    exp_41_ram[520] = 111;
    exp_41_ram[521] = 99;
    exp_41_ram[522] = 147;
    exp_41_ram[523] = 179;
    exp_41_ram[524] = 99;
    exp_41_ram[525] = 147;
    exp_41_ram[526] = 19;
    exp_41_ram[527] = 179;
    exp_41_ram[528] = 19;
    exp_41_ram[529] = 103;
    exp_41_ram[530] = 51;
    exp_41_ram[531] = 179;
    exp_41_ram[532] = 51;
    exp_41_ram[533] = 179;
    exp_41_ram[534] = 111;
    exp_41_ram[535] = 183;
    exp_41_ram[536] = 99;
    exp_41_ram[537] = 147;
    exp_41_ram[538] = 179;
    exp_41_ram[539] = 147;
    exp_41_ram[540] = 55;
    exp_41_ram[541] = 147;
    exp_41_ram[542] = 179;
    exp_41_ram[543] = 51;
    exp_41_ram[544] = 147;
    exp_41_ram[545] = 51;
    exp_41_ram[546] = 3;
    exp_41_ram[547] = 51;
    exp_41_ram[548] = 103;
    exp_41_ram[549] = 55;
    exp_41_ram[550] = 147;
    exp_41_ram[551] = 227;
    exp_41_ram[552] = 147;
    exp_41_ram[553] = 111;
    exp_41_ram[554] = 83;
    exp_41_ram[555] = 111;
    exp_41_ram[556] = 101;
    exp_41_ram[557] = 84;
    exp_41_ram[558] = 114;
    exp_41_ram[559] = 116;
    exp_41_ram[560] = 74;
    exp_41_ram[561] = 101;
    exp_41_ram[562] = 114;
    exp_41_ram[563] = 77;
    exp_41_ram[564] = 117;
    exp_41_ram[565] = 108;
    exp_41_ram[566] = 83;
    exp_41_ram[567] = 99;
    exp_41_ram[568] = 118;
    exp_41_ram[569] = 0;
    exp_41_ram[570] = 72;
    exp_41_ram[571] = 111;
    exp_41_ram[572] = 114;
    exp_41_ram[573] = 0;
    exp_41_ram[574] = 114;
    exp_41_ram[575] = 105;
    exp_41_ram[576] = 107;
    exp_41_ram[577] = 104;
    exp_41_ram[578] = 105;
    exp_41_ram[579] = 32;
    exp_41_ram[580] = 111;
    exp_41_ram[581] = 0;
    exp_41_ram[582] = 114;
    exp_41_ram[583] = 105;
    exp_41_ram[584] = 80;
    exp_41_ram[585] = 100;
    exp_41_ram[586] = 46;
    exp_41_ram[587] = 32;
    exp_41_ram[588] = 98;
    exp_41_ram[589] = 105;
    exp_41_ram[590] = 103;
    exp_41_ram[591] = 109;
    exp_41_ram[592] = 105;
    exp_41_ram[593] = 101;
    exp_41_ram[594] = 110;
    exp_41_ram[595] = 115;
    exp_41_ram[596] = 110;
    exp_41_ram[597] = 32;
    exp_41_ram[598] = 98;
    exp_41_ram[599] = 105;
    exp_41_ram[600] = 103;
    exp_41_ram[601] = 109;
    exp_41_ram[602] = 105;
    exp_41_ram[603] = 101;
    exp_41_ram[604] = 110;
    exp_41_ram[605] = 115;
    exp_41_ram[606] = 110;
    exp_41_ram[607] = 32;
    exp_41_ram[608] = 98;
    exp_41_ram[609] = 105;
    exp_41_ram[610] = 103;
    exp_41_ram[611] = 100;
    exp_41_ram[612] = 100;
    exp_41_ram[613] = 105;
    exp_41_ram[614] = 32;
    exp_41_ram[615] = 111;
    exp_41_ram[616] = 32;
    exp_41_ram[617] = 98;
    exp_41_ram[618] = 105;
    exp_41_ram[619] = 103;
    exp_41_ram[620] = 100;
    exp_41_ram[621] = 100;
    exp_41_ram[622] = 105;
    exp_41_ram[623] = 32;
    exp_41_ram[624] = 111;
    exp_41_ram[625] = 89;
    exp_41_ram[626] = 58;
    exp_41_ram[627] = 77;
    exp_41_ram[628] = 104;
    exp_41_ram[629] = 68;
    exp_41_ram[630] = 0;
    exp_41_ram[631] = 72;
    exp_41_ram[632] = 58;
    exp_41_ram[633] = 77;
    exp_41_ram[634] = 116;
    exp_41_ram[635] = 10;
    exp_41_ram[636] = 112;
    exp_41_ram[637] = 32;
    exp_41_ram[638] = 111;
    exp_41_ram[639] = 10;
    exp_41_ram[640] = 72;
    exp_41_ram[641] = 111;
    exp_41_ram[642] = 114;
    exp_41_ram[643] = 98;
    exp_41_ram[644] = 110;
    exp_41_ram[645] = 116;
    exp_41_ram[646] = 100;
    exp_41_ram[647] = 99;
    exp_41_ram[648] = 101;
    exp_41_ram[649] = 77;
    exp_41_ram[650] = 105;
    exp_41_ram[651] = 99;
    exp_41_ram[652] = 111;
    exp_41_ram[653] = 100;
    exp_41_ram[654] = 97;
    exp_41_ram[655] = 67;
    exp_41_ram[656] = 107;
    exp_41_ram[657] = 101;
    exp_41_ram[658] = 110;
    exp_41_ram[659] = 97;
    exp_41_ram[660] = 99;
    exp_41_ram[661] = 101;
    exp_41_ram[662] = 102;
    exp_41_ram[663] = 87;
    exp_41_ram[664] = 101;
    exp_41_ram[665] = 82;
    exp_41_ram[666] = 114;
    exp_41_ram[667] = 115;
    exp_41_ram[668] = 111;
    exp_41_ram[669] = 32;
    exp_41_ram[670] = 10;
    exp_41_ram[671] = 69;
    exp_41_ram[672] = 109;
    exp_41_ram[673] = 97;
    exp_41_ram[674] = 110;
    exp_41_ram[675] = 61;
    exp_41_ram[676] = 61;
    exp_41_ram[677] = 61;
    exp_41_ram[678] = 61;
    exp_41_ram[679] = 0;
    exp_41_ram[680] = 49;
    exp_41_ram[681] = 104;
    exp_41_ram[682] = 32;
    exp_41_ram[683] = 116;
    exp_41_ram[684] = 115;
    exp_41_ram[685] = 97;
    exp_41_ram[686] = 110;
    exp_41_ram[687] = 101;
    exp_41_ram[688] = 49;
    exp_41_ram[689] = 41;
    exp_41_ram[690] = 102;
    exp_41_ram[691] = 109;
    exp_41_ram[692] = 108;
    exp_41_ram[693] = 114;
    exp_41_ram[694] = 116;
    exp_41_ram[695] = 103;
    exp_41_ram[696] = 50;
    exp_41_ram[697] = 50;
    exp_41_ram[698] = 101;
    exp_41_ram[699] = 99;
    exp_41_ram[700] = 32;
    exp_41_ram[701] = 62;
    exp_41_ram[702] = 101;
    exp_41_ram[703] = 32;
    exp_41_ram[704] = 51;
    exp_41_ram[705] = 105;
    exp_41_ram[706] = 115;
    exp_41_ram[707] = 105;
    exp_41_ram[708] = 32;
    exp_41_ram[709] = 110;
    exp_41_ram[710] = 101;
    exp_41_ram[711] = 110;
    exp_41_ram[712] = 40;
    exp_41_ram[713] = 122;
    exp_41_ram[714] = 101;
    exp_41_ram[715] = 32;
    exp_41_ram[716] = 100;
    exp_41_ram[717] = 32;
    exp_41_ram[718] = 104;
    exp_41_ram[719] = 46;
    exp_41_ram[720] = 97;
    exp_41_ram[721] = 0;
    exp_41_ram[722] = 52;
    exp_41_ram[723] = 111;
    exp_41_ram[724] = 32;
    exp_41_ram[725] = 105;
    exp_41_ram[726] = 110;
    exp_41_ram[727] = 97;
    exp_41_ram[728] = 41;
    exp_41_ram[729] = 102;
    exp_41_ram[730] = 109;
    exp_41_ram[731] = 108;
    exp_41_ram[732] = 114;
    exp_41_ram[733] = 116;
    exp_41_ram[734] = 103;
    exp_41_ram[735] = 97;
    exp_41_ram[736] = 114;
    exp_41_ram[737] = 121;
    exp_41_ram[738] = 46;
    exp_41_ram[739] = 58;
    exp_41_ram[740] = 10;
    exp_41_ram[741] = 0;
    exp_41_ram[742] = 3;
    exp_41_ram[743] = 4;
    exp_41_ram[744] = 4;
    exp_41_ram[745] = 5;
    exp_41_ram[746] = 5;
    exp_41_ram[747] = 5;
    exp_41_ram[748] = 5;
    exp_41_ram[749] = 6;
    exp_41_ram[750] = 6;
    exp_41_ram[751] = 6;
    exp_41_ram[752] = 6;
    exp_41_ram[753] = 6;
    exp_41_ram[754] = 6;
    exp_41_ram[755] = 6;
    exp_41_ram[756] = 6;
    exp_41_ram[757] = 7;
    exp_41_ram[758] = 7;
    exp_41_ram[759] = 7;
    exp_41_ram[760] = 7;
    exp_41_ram[761] = 7;
    exp_41_ram[762] = 7;
    exp_41_ram[763] = 7;
    exp_41_ram[764] = 7;
    exp_41_ram[765] = 7;
    exp_41_ram[766] = 7;
    exp_41_ram[767] = 7;
    exp_41_ram[768] = 7;
    exp_41_ram[769] = 7;
    exp_41_ram[770] = 7;
    exp_41_ram[771] = 7;
    exp_41_ram[772] = 7;
    exp_41_ram[773] = 8;
    exp_41_ram[774] = 8;
    exp_41_ram[775] = 8;
    exp_41_ram[776] = 8;
    exp_41_ram[777] = 8;
    exp_41_ram[778] = 8;
    exp_41_ram[779] = 8;
    exp_41_ram[780] = 8;
    exp_41_ram[781] = 8;
    exp_41_ram[782] = 8;
    exp_41_ram[783] = 8;
    exp_41_ram[784] = 8;
    exp_41_ram[785] = 8;
    exp_41_ram[786] = 8;
    exp_41_ram[787] = 8;
    exp_41_ram[788] = 8;
    exp_41_ram[789] = 8;
    exp_41_ram[790] = 8;
    exp_41_ram[791] = 8;
    exp_41_ram[792] = 8;
    exp_41_ram[793] = 8;
    exp_41_ram[794] = 8;
    exp_41_ram[795] = 8;
    exp_41_ram[796] = 8;
    exp_41_ram[797] = 8;
    exp_41_ram[798] = 8;
    exp_41_ram[799] = 8;
    exp_41_ram[800] = 8;
    exp_41_ram[801] = 8;
    exp_41_ram[802] = 8;
    exp_41_ram[803] = 8;
    exp_41_ram[804] = 8;
    exp_41_ram[805] = 19;
    exp_41_ram[806] = 35;
    exp_41_ram[807] = 19;
    exp_41_ram[808] = 35;
    exp_41_ram[809] = 131;
    exp_41_ram[810] = 35;
    exp_41_ram[811] = 131;
    exp_41_ram[812] = 131;
    exp_41_ram[813] = 19;
    exp_41_ram[814] = 3;
    exp_41_ram[815] = 19;
    exp_41_ram[816] = 103;
    exp_41_ram[817] = 19;
    exp_41_ram[818] = 35;
    exp_41_ram[819] = 19;
    exp_41_ram[820] = 35;
    exp_41_ram[821] = 35;
    exp_41_ram[822] = 131;
    exp_41_ram[823] = 35;
    exp_41_ram[824] = 3;
    exp_41_ram[825] = 131;
    exp_41_ram[826] = 35;
    exp_41_ram[827] = 131;
    exp_41_ram[828] = 19;
    exp_41_ram[829] = 3;
    exp_41_ram[830] = 19;
    exp_41_ram[831] = 103;
    exp_41_ram[832] = 19;
    exp_41_ram[833] = 35;
    exp_41_ram[834] = 35;
    exp_41_ram[835] = 19;
    exp_41_ram[836] = 35;
    exp_41_ram[837] = 183;
    exp_41_ram[838] = 131;
    exp_41_ram[839] = 147;
    exp_41_ram[840] = 3;
    exp_41_ram[841] = 239;
    exp_41_ram[842] = 147;
    exp_41_ram[843] = 19;
    exp_41_ram[844] = 131;
    exp_41_ram[845] = 3;
    exp_41_ram[846] = 19;
    exp_41_ram[847] = 103;
    exp_41_ram[848] = 19;
    exp_41_ram[849] = 35;
    exp_41_ram[850] = 35;
    exp_41_ram[851] = 19;
    exp_41_ram[852] = 183;
    exp_41_ram[853] = 131;
    exp_41_ram[854] = 19;
    exp_41_ram[855] = 239;
    exp_41_ram[856] = 147;
    exp_41_ram[857] = 19;
    exp_41_ram[858] = 131;
    exp_41_ram[859] = 3;
    exp_41_ram[860] = 19;
    exp_41_ram[861] = 103;
    exp_41_ram[862] = 19;
    exp_41_ram[863] = 35;
    exp_41_ram[864] = 35;
    exp_41_ram[865] = 19;
    exp_41_ram[866] = 35;
    exp_41_ram[867] = 35;
    exp_41_ram[868] = 35;
    exp_41_ram[869] = 111;
    exp_41_ram[870] = 131;
    exp_41_ram[871] = 19;
    exp_41_ram[872] = 35;
    exp_41_ram[873] = 3;
    exp_41_ram[874] = 179;
    exp_41_ram[875] = 131;
    exp_41_ram[876] = 131;
    exp_41_ram[877] = 19;
    exp_41_ram[878] = 239;
    exp_41_ram[879] = 3;
    exp_41_ram[880] = 131;
    exp_41_ram[881] = 179;
    exp_41_ram[882] = 131;
    exp_41_ram[883] = 227;
    exp_41_ram[884] = 131;
    exp_41_ram[885] = 19;
    exp_41_ram[886] = 131;
    exp_41_ram[887] = 3;
    exp_41_ram[888] = 19;
    exp_41_ram[889] = 103;
    exp_41_ram[890] = 19;
    exp_41_ram[891] = 35;
    exp_41_ram[892] = 35;
    exp_41_ram[893] = 19;
    exp_41_ram[894] = 35;
    exp_41_ram[895] = 183;
    exp_41_ram[896] = 131;
    exp_41_ram[897] = 147;
    exp_41_ram[898] = 3;
    exp_41_ram[899] = 239;
    exp_41_ram[900] = 183;
    exp_41_ram[901] = 131;
    exp_41_ram[902] = 147;
    exp_41_ram[903] = 19;
    exp_41_ram[904] = 239;
    exp_41_ram[905] = 147;
    exp_41_ram[906] = 19;
    exp_41_ram[907] = 131;
    exp_41_ram[908] = 3;
    exp_41_ram[909] = 19;
    exp_41_ram[910] = 103;
    exp_41_ram[911] = 19;
    exp_41_ram[912] = 35;
    exp_41_ram[913] = 19;
    exp_41_ram[914] = 35;
    exp_41_ram[915] = 3;
    exp_41_ram[916] = 147;
    exp_41_ram[917] = 99;
    exp_41_ram[918] = 3;
    exp_41_ram[919] = 147;
    exp_41_ram[920] = 99;
    exp_41_ram[921] = 3;
    exp_41_ram[922] = 147;
    exp_41_ram[923] = 99;
    exp_41_ram[924] = 3;
    exp_41_ram[925] = 147;
    exp_41_ram[926] = 99;
    exp_41_ram[927] = 147;
    exp_41_ram[928] = 111;
    exp_41_ram[929] = 147;
    exp_41_ram[930] = 19;
    exp_41_ram[931] = 3;
    exp_41_ram[932] = 19;
    exp_41_ram[933] = 103;
    exp_41_ram[934] = 19;
    exp_41_ram[935] = 35;
    exp_41_ram[936] = 19;
    exp_41_ram[937] = 35;
    exp_41_ram[938] = 3;
    exp_41_ram[939] = 147;
    exp_41_ram[940] = 99;
    exp_41_ram[941] = 3;
    exp_41_ram[942] = 147;
    exp_41_ram[943] = 99;
    exp_41_ram[944] = 147;
    exp_41_ram[945] = 111;
    exp_41_ram[946] = 147;
    exp_41_ram[947] = 19;
    exp_41_ram[948] = 3;
    exp_41_ram[949] = 19;
    exp_41_ram[950] = 103;
    exp_41_ram[951] = 19;
    exp_41_ram[952] = 35;
    exp_41_ram[953] = 35;
    exp_41_ram[954] = 19;
    exp_41_ram[955] = 35;
    exp_41_ram[956] = 3;
    exp_41_ram[957] = 239;
    exp_41_ram[958] = 147;
    exp_41_ram[959] = 99;
    exp_41_ram[960] = 131;
    exp_41_ram[961] = 147;
    exp_41_ram[962] = 111;
    exp_41_ram[963] = 131;
    exp_41_ram[964] = 19;
    exp_41_ram[965] = 131;
    exp_41_ram[966] = 3;
    exp_41_ram[967] = 19;
    exp_41_ram[968] = 103;
    exp_41_ram[969] = 19;
    exp_41_ram[970] = 35;
    exp_41_ram[971] = 35;
    exp_41_ram[972] = 35;
    exp_41_ram[973] = 19;
    exp_41_ram[974] = 147;
    exp_41_ram[975] = 131;
    exp_41_ram[976] = 35;
    exp_41_ram[977] = 147;
    exp_41_ram[978] = 35;
    exp_41_ram[979] = 147;
    exp_41_ram[980] = 35;
    exp_41_ram[981] = 147;
    exp_41_ram[982] = 35;
    exp_41_ram[983] = 35;
    exp_41_ram[984] = 35;
    exp_41_ram[985] = 35;
    exp_41_ram[986] = 3;
    exp_41_ram[987] = 131;
    exp_41_ram[988] = 3;
    exp_41_ram[989] = 3;
    exp_41_ram[990] = 131;
    exp_41_ram[991] = 3;
    exp_41_ram[992] = 131;
    exp_41_ram[993] = 3;
    exp_41_ram[994] = 131;
    exp_41_ram[995] = 35;
    exp_41_ram[996] = 35;
    exp_41_ram[997] = 35;
    exp_41_ram[998] = 35;
    exp_41_ram[999] = 35;
    exp_41_ram[1000] = 35;
    exp_41_ram[1001] = 35;
    exp_41_ram[1002] = 35;
    exp_41_ram[1003] = 35;
    exp_41_ram[1004] = 147;
    exp_41_ram[1005] = 19;
    exp_41_ram[1006] = 239;
    exp_41_ram[1007] = 35;
    exp_41_ram[1008] = 35;
    exp_41_ram[1009] = 147;
    exp_41_ram[1010] = 131;
    exp_41_ram[1011] = 3;
    exp_41_ram[1012] = 19;
    exp_41_ram[1013] = 239;
    exp_41_ram[1014] = 3;
    exp_41_ram[1015] = 131;
    exp_41_ram[1016] = 179;
    exp_41_ram[1017] = 35;
    exp_41_ram[1018] = 3;
    exp_41_ram[1019] = 131;
    exp_41_ram[1020] = 3;
    exp_41_ram[1021] = 3;
    exp_41_ram[1022] = 131;
    exp_41_ram[1023] = 3;
    exp_41_ram[1024] = 131;
    exp_41_ram[1025] = 3;
    exp_41_ram[1026] = 131;
    exp_41_ram[1027] = 35;
    exp_41_ram[1028] = 35;
    exp_41_ram[1029] = 35;
    exp_41_ram[1030] = 35;
    exp_41_ram[1031] = 35;
    exp_41_ram[1032] = 35;
    exp_41_ram[1033] = 35;
    exp_41_ram[1034] = 35;
    exp_41_ram[1035] = 35;
    exp_41_ram[1036] = 147;
    exp_41_ram[1037] = 19;
    exp_41_ram[1038] = 239;
    exp_41_ram[1039] = 35;
    exp_41_ram[1040] = 35;
    exp_41_ram[1041] = 131;
    exp_41_ram[1042] = 35;
    exp_41_ram[1043] = 147;
    exp_41_ram[1044] = 35;
    exp_41_ram[1045] = 147;
    exp_41_ram[1046] = 35;
    exp_41_ram[1047] = 147;
    exp_41_ram[1048] = 35;
    exp_41_ram[1049] = 35;
    exp_41_ram[1050] = 35;
    exp_41_ram[1051] = 35;
    exp_41_ram[1052] = 3;
    exp_41_ram[1053] = 131;
    exp_41_ram[1054] = 3;
    exp_41_ram[1055] = 3;
    exp_41_ram[1056] = 131;
    exp_41_ram[1057] = 3;
    exp_41_ram[1058] = 131;
    exp_41_ram[1059] = 3;
    exp_41_ram[1060] = 131;
    exp_41_ram[1061] = 35;
    exp_41_ram[1062] = 35;
    exp_41_ram[1063] = 35;
    exp_41_ram[1064] = 35;
    exp_41_ram[1065] = 35;
    exp_41_ram[1066] = 35;
    exp_41_ram[1067] = 35;
    exp_41_ram[1068] = 35;
    exp_41_ram[1069] = 35;
    exp_41_ram[1070] = 147;
    exp_41_ram[1071] = 19;
    exp_41_ram[1072] = 239;
    exp_41_ram[1073] = 35;
    exp_41_ram[1074] = 35;
    exp_41_ram[1075] = 147;
    exp_41_ram[1076] = 131;
    exp_41_ram[1077] = 3;
    exp_41_ram[1078] = 19;
    exp_41_ram[1079] = 239;
    exp_41_ram[1080] = 3;
    exp_41_ram[1081] = 131;
    exp_41_ram[1082] = 179;
    exp_41_ram[1083] = 35;
    exp_41_ram[1084] = 3;
    exp_41_ram[1085] = 131;
    exp_41_ram[1086] = 3;
    exp_41_ram[1087] = 3;
    exp_41_ram[1088] = 131;
    exp_41_ram[1089] = 3;
    exp_41_ram[1090] = 131;
    exp_41_ram[1091] = 3;
    exp_41_ram[1092] = 131;
    exp_41_ram[1093] = 35;
    exp_41_ram[1094] = 35;
    exp_41_ram[1095] = 35;
    exp_41_ram[1096] = 35;
    exp_41_ram[1097] = 35;
    exp_41_ram[1098] = 35;
    exp_41_ram[1099] = 35;
    exp_41_ram[1100] = 35;
    exp_41_ram[1101] = 35;
    exp_41_ram[1102] = 147;
    exp_41_ram[1103] = 19;
    exp_41_ram[1104] = 239;
    exp_41_ram[1105] = 35;
    exp_41_ram[1106] = 35;
    exp_41_ram[1107] = 3;
    exp_41_ram[1108] = 131;
    exp_41_ram[1109] = 3;
    exp_41_ram[1110] = 3;
    exp_41_ram[1111] = 131;
    exp_41_ram[1112] = 3;
    exp_41_ram[1113] = 131;
    exp_41_ram[1114] = 3;
    exp_41_ram[1115] = 131;
    exp_41_ram[1116] = 35;
    exp_41_ram[1117] = 35;
    exp_41_ram[1118] = 35;
    exp_41_ram[1119] = 35;
    exp_41_ram[1120] = 35;
    exp_41_ram[1121] = 35;
    exp_41_ram[1122] = 35;
    exp_41_ram[1123] = 35;
    exp_41_ram[1124] = 35;
    exp_41_ram[1125] = 147;
    exp_41_ram[1126] = 19;
    exp_41_ram[1127] = 239;
    exp_41_ram[1128] = 35;
    exp_41_ram[1129] = 35;
    exp_41_ram[1130] = 3;
    exp_41_ram[1131] = 131;
    exp_41_ram[1132] = 99;
    exp_41_ram[1133] = 3;
    exp_41_ram[1134] = 131;
    exp_41_ram[1135] = 99;
    exp_41_ram[1136] = 3;
    exp_41_ram[1137] = 131;
    exp_41_ram[1138] = 99;
    exp_41_ram[1139] = 3;
    exp_41_ram[1140] = 131;
    exp_41_ram[1141] = 99;
    exp_41_ram[1142] = 3;
    exp_41_ram[1143] = 131;
    exp_41_ram[1144] = 99;
    exp_41_ram[1145] = 3;
    exp_41_ram[1146] = 131;
    exp_41_ram[1147] = 99;
    exp_41_ram[1148] = 147;
    exp_41_ram[1149] = 111;
    exp_41_ram[1150] = 147;
    exp_41_ram[1151] = 19;
    exp_41_ram[1152] = 131;
    exp_41_ram[1153] = 3;
    exp_41_ram[1154] = 131;
    exp_41_ram[1155] = 19;
    exp_41_ram[1156] = 103;
    exp_41_ram[1157] = 19;
    exp_41_ram[1158] = 35;
    exp_41_ram[1159] = 35;
    exp_41_ram[1160] = 19;
    exp_41_ram[1161] = 35;
    exp_41_ram[1162] = 35;
    exp_41_ram[1163] = 147;
    exp_41_ram[1164] = 131;
    exp_41_ram[1165] = 3;
    exp_41_ram[1166] = 19;
    exp_41_ram[1167] = 239;
    exp_41_ram[1168] = 3;
    exp_41_ram[1169] = 131;
    exp_41_ram[1170] = 3;
    exp_41_ram[1171] = 3;
    exp_41_ram[1172] = 131;
    exp_41_ram[1173] = 3;
    exp_41_ram[1174] = 131;
    exp_41_ram[1175] = 3;
    exp_41_ram[1176] = 131;
    exp_41_ram[1177] = 35;
    exp_41_ram[1178] = 35;
    exp_41_ram[1179] = 35;
    exp_41_ram[1180] = 35;
    exp_41_ram[1181] = 35;
    exp_41_ram[1182] = 35;
    exp_41_ram[1183] = 35;
    exp_41_ram[1184] = 35;
    exp_41_ram[1185] = 35;
    exp_41_ram[1186] = 147;
    exp_41_ram[1187] = 19;
    exp_41_ram[1188] = 239;
    exp_41_ram[1189] = 147;
    exp_41_ram[1190] = 19;
    exp_41_ram[1191] = 131;
    exp_41_ram[1192] = 3;
    exp_41_ram[1193] = 19;
    exp_41_ram[1194] = 103;
    exp_41_ram[1195] = 19;
    exp_41_ram[1196] = 35;
    exp_41_ram[1197] = 19;
    exp_41_ram[1198] = 183;
    exp_41_ram[1199] = 35;
    exp_41_ram[1200] = 183;
    exp_41_ram[1201] = 147;
    exp_41_ram[1202] = 35;
    exp_41_ram[1203] = 131;
    exp_41_ram[1204] = 131;
    exp_41_ram[1205] = 35;
    exp_41_ram[1206] = 35;
    exp_41_ram[1207] = 131;
    exp_41_ram[1208] = 147;
    exp_41_ram[1209] = 35;
    exp_41_ram[1210] = 35;
    exp_41_ram[1211] = 131;
    exp_41_ram[1212] = 131;
    exp_41_ram[1213] = 19;
    exp_41_ram[1214] = 147;
    exp_41_ram[1215] = 131;
    exp_41_ram[1216] = 179;
    exp_41_ram[1217] = 35;
    exp_41_ram[1218] = 131;
    exp_41_ram[1219] = 179;
    exp_41_ram[1220] = 35;
    exp_41_ram[1221] = 3;
    exp_41_ram[1222] = 131;
    exp_41_ram[1223] = 19;
    exp_41_ram[1224] = 147;
    exp_41_ram[1225] = 3;
    exp_41_ram[1226] = 19;
    exp_41_ram[1227] = 103;
    exp_41_ram[1228] = 19;
    exp_41_ram[1229] = 35;
    exp_41_ram[1230] = 35;
    exp_41_ram[1231] = 19;
    exp_41_ram[1232] = 35;
    exp_41_ram[1233] = 35;
    exp_41_ram[1234] = 35;
    exp_41_ram[1235] = 35;
    exp_41_ram[1236] = 3;
    exp_41_ram[1237] = 131;
    exp_41_ram[1238] = 3;
    exp_41_ram[1239] = 131;
    exp_41_ram[1240] = 51;
    exp_41_ram[1241] = 19;
    exp_41_ram[1242] = 51;
    exp_41_ram[1243] = 179;
    exp_41_ram[1244] = 179;
    exp_41_ram[1245] = 147;
    exp_41_ram[1246] = 19;
    exp_41_ram[1247] = 147;
    exp_41_ram[1248] = 19;
    exp_41_ram[1249] = 147;
    exp_41_ram[1250] = 239;
    exp_41_ram[1251] = 19;
    exp_41_ram[1252] = 147;
    exp_41_ram[1253] = 19;
    exp_41_ram[1254] = 147;
    exp_41_ram[1255] = 131;
    exp_41_ram[1256] = 3;
    exp_41_ram[1257] = 19;
    exp_41_ram[1258] = 103;
    exp_41_ram[1259] = 19;
    exp_41_ram[1260] = 35;
    exp_41_ram[1261] = 19;
    exp_41_ram[1262] = 35;
    exp_41_ram[1263] = 131;
    exp_41_ram[1264] = 147;
    exp_41_ram[1265] = 99;
    exp_41_ram[1266] = 3;
    exp_41_ram[1267] = 147;
    exp_41_ram[1268] = 179;
    exp_41_ram[1269] = 99;
    exp_41_ram[1270] = 3;
    exp_41_ram[1271] = 147;
    exp_41_ram[1272] = 179;
    exp_41_ram[1273] = 99;
    exp_41_ram[1274] = 147;
    exp_41_ram[1275] = 111;
    exp_41_ram[1276] = 147;
    exp_41_ram[1277] = 19;
    exp_41_ram[1278] = 3;
    exp_41_ram[1279] = 19;
    exp_41_ram[1280] = 103;
    exp_41_ram[1281] = 19;
    exp_41_ram[1282] = 35;
    exp_41_ram[1283] = 35;
    exp_41_ram[1284] = 19;
    exp_41_ram[1285] = 35;
    exp_41_ram[1286] = 3;
    exp_41_ram[1287] = 239;
    exp_41_ram[1288] = 147;
    exp_41_ram[1289] = 99;
    exp_41_ram[1290] = 147;
    exp_41_ram[1291] = 111;
    exp_41_ram[1292] = 147;
    exp_41_ram[1293] = 19;
    exp_41_ram[1294] = 131;
    exp_41_ram[1295] = 3;
    exp_41_ram[1296] = 19;
    exp_41_ram[1297] = 103;
    exp_41_ram[1298] = 19;
    exp_41_ram[1299] = 35;
    exp_41_ram[1300] = 35;
    exp_41_ram[1301] = 19;
    exp_41_ram[1302] = 35;
    exp_41_ram[1303] = 35;
    exp_41_ram[1304] = 3;
    exp_41_ram[1305] = 147;
    exp_41_ram[1306] = 99;
    exp_41_ram[1307] = 3;
    exp_41_ram[1308] = 147;
    exp_41_ram[1309] = 99;
    exp_41_ram[1310] = 3;
    exp_41_ram[1311] = 147;
    exp_41_ram[1312] = 99;
    exp_41_ram[1313] = 3;
    exp_41_ram[1314] = 147;
    exp_41_ram[1315] = 99;
    exp_41_ram[1316] = 147;
    exp_41_ram[1317] = 111;
    exp_41_ram[1318] = 3;
    exp_41_ram[1319] = 147;
    exp_41_ram[1320] = 99;
    exp_41_ram[1321] = 3;
    exp_41_ram[1322] = 239;
    exp_41_ram[1323] = 147;
    exp_41_ram[1324] = 99;
    exp_41_ram[1325] = 147;
    exp_41_ram[1326] = 111;
    exp_41_ram[1327] = 147;
    exp_41_ram[1328] = 111;
    exp_41_ram[1329] = 147;
    exp_41_ram[1330] = 19;
    exp_41_ram[1331] = 131;
    exp_41_ram[1332] = 3;
    exp_41_ram[1333] = 19;
    exp_41_ram[1334] = 103;
    exp_41_ram[1335] = 19;
    exp_41_ram[1336] = 35;
    exp_41_ram[1337] = 35;
    exp_41_ram[1338] = 35;
    exp_41_ram[1339] = 35;
    exp_41_ram[1340] = 35;
    exp_41_ram[1341] = 35;
    exp_41_ram[1342] = 35;
    exp_41_ram[1343] = 35;
    exp_41_ram[1344] = 35;
    exp_41_ram[1345] = 35;
    exp_41_ram[1346] = 35;
    exp_41_ram[1347] = 35;
    exp_41_ram[1348] = 35;
    exp_41_ram[1349] = 19;
    exp_41_ram[1350] = 147;
    exp_41_ram[1351] = 147;
    exp_41_ram[1352] = 19;
    exp_41_ram[1353] = 35;
    exp_41_ram[1354] = 35;
    exp_41_ram[1355] = 147;
    exp_41_ram[1356] = 35;
    exp_41_ram[1357] = 131;
    exp_41_ram[1358] = 35;
    exp_41_ram[1359] = 131;
    exp_41_ram[1360] = 147;
    exp_41_ram[1361] = 3;
    exp_41_ram[1362] = 99;
    exp_41_ram[1363] = 3;
    exp_41_ram[1364] = 239;
    exp_41_ram[1365] = 19;
    exp_41_ram[1366] = 183;
    exp_41_ram[1367] = 147;
    exp_41_ram[1368] = 179;
    exp_41_ram[1369] = 35;
    exp_41_ram[1370] = 35;
    exp_41_ram[1371] = 3;
    exp_41_ram[1372] = 131;
    exp_41_ram[1373] = 3;
    exp_41_ram[1374] = 131;
    exp_41_ram[1375] = 147;
    exp_41_ram[1376] = 51;
    exp_41_ram[1377] = 147;
    exp_41_ram[1378] = 179;
    exp_41_ram[1379] = 19;
    exp_41_ram[1380] = 179;
    exp_41_ram[1381] = 179;
    exp_41_ram[1382] = 147;
    exp_41_ram[1383] = 35;
    exp_41_ram[1384] = 35;
    exp_41_ram[1385] = 131;
    exp_41_ram[1386] = 147;
    exp_41_ram[1387] = 35;
    exp_41_ram[1388] = 111;
    exp_41_ram[1389] = 19;
    exp_41_ram[1390] = 35;
    exp_41_ram[1391] = 131;
    exp_41_ram[1392] = 19;
    exp_41_ram[1393] = 131;
    exp_41_ram[1394] = 99;
    exp_41_ram[1395] = 131;
    exp_41_ram[1396] = 3;
    exp_41_ram[1397] = 239;
    exp_41_ram[1398] = 19;
    exp_41_ram[1399] = 183;
    exp_41_ram[1400] = 147;
    exp_41_ram[1401] = 179;
    exp_41_ram[1402] = 19;
    exp_41_ram[1403] = 147;
    exp_41_ram[1404] = 3;
    exp_41_ram[1405] = 131;
    exp_41_ram[1406] = 51;
    exp_41_ram[1407] = 147;
    exp_41_ram[1408] = 179;
    exp_41_ram[1409] = 179;
    exp_41_ram[1410] = 179;
    exp_41_ram[1411] = 147;
    exp_41_ram[1412] = 35;
    exp_41_ram[1413] = 35;
    exp_41_ram[1414] = 131;
    exp_41_ram[1415] = 147;
    exp_41_ram[1416] = 35;
    exp_41_ram[1417] = 111;
    exp_41_ram[1418] = 19;
    exp_41_ram[1419] = 131;
    exp_41_ram[1420] = 19;
    exp_41_ram[1421] = 183;
    exp_41_ram[1422] = 147;
    exp_41_ram[1423] = 179;
    exp_41_ram[1424] = 19;
    exp_41_ram[1425] = 147;
    exp_41_ram[1426] = 147;
    exp_41_ram[1427] = 3;
    exp_41_ram[1428] = 131;
    exp_41_ram[1429] = 51;
    exp_41_ram[1430] = 147;
    exp_41_ram[1431] = 179;
    exp_41_ram[1432] = 179;
    exp_41_ram[1433] = 179;
    exp_41_ram[1434] = 147;
    exp_41_ram[1435] = 35;
    exp_41_ram[1436] = 35;
    exp_41_ram[1437] = 3;
    exp_41_ram[1438] = 183;
    exp_41_ram[1439] = 147;
    exp_41_ram[1440] = 179;
    exp_41_ram[1441] = 19;
    exp_41_ram[1442] = 147;
    exp_41_ram[1443] = 147;
    exp_41_ram[1444] = 3;
    exp_41_ram[1445] = 131;
    exp_41_ram[1446] = 51;
    exp_41_ram[1447] = 147;
    exp_41_ram[1448] = 179;
    exp_41_ram[1449] = 179;
    exp_41_ram[1450] = 179;
    exp_41_ram[1451] = 147;
    exp_41_ram[1452] = 35;
    exp_41_ram[1453] = 35;
    exp_41_ram[1454] = 3;
    exp_41_ram[1455] = 147;
    exp_41_ram[1456] = 147;
    exp_41_ram[1457] = 179;
    exp_41_ram[1458] = 147;
    exp_41_ram[1459] = 19;
    exp_41_ram[1460] = 147;
    exp_41_ram[1461] = 147;
    exp_41_ram[1462] = 3;
    exp_41_ram[1463] = 131;
    exp_41_ram[1464] = 51;
    exp_41_ram[1465] = 147;
    exp_41_ram[1466] = 179;
    exp_41_ram[1467] = 179;
    exp_41_ram[1468] = 179;
    exp_41_ram[1469] = 147;
    exp_41_ram[1470] = 35;
    exp_41_ram[1471] = 35;
    exp_41_ram[1472] = 131;
    exp_41_ram[1473] = 19;
    exp_41_ram[1474] = 147;
    exp_41_ram[1475] = 147;
    exp_41_ram[1476] = 3;
    exp_41_ram[1477] = 131;
    exp_41_ram[1478] = 51;
    exp_41_ram[1479] = 147;
    exp_41_ram[1480] = 179;
    exp_41_ram[1481] = 179;
    exp_41_ram[1482] = 179;
    exp_41_ram[1483] = 147;
    exp_41_ram[1484] = 35;
    exp_41_ram[1485] = 35;
    exp_41_ram[1486] = 3;
    exp_41_ram[1487] = 131;
    exp_41_ram[1488] = 19;
    exp_41_ram[1489] = 147;
    exp_41_ram[1490] = 131;
    exp_41_ram[1491] = 3;
    exp_41_ram[1492] = 131;
    exp_41_ram[1493] = 3;
    exp_41_ram[1494] = 131;
    exp_41_ram[1495] = 3;
    exp_41_ram[1496] = 131;
    exp_41_ram[1497] = 3;
    exp_41_ram[1498] = 131;
    exp_41_ram[1499] = 3;
    exp_41_ram[1500] = 131;
    exp_41_ram[1501] = 3;
    exp_41_ram[1502] = 131;
    exp_41_ram[1503] = 19;
    exp_41_ram[1504] = 103;
    exp_41_ram[1505] = 19;
    exp_41_ram[1506] = 35;
    exp_41_ram[1507] = 35;
    exp_41_ram[1508] = 35;
    exp_41_ram[1509] = 35;
    exp_41_ram[1510] = 35;
    exp_41_ram[1511] = 19;
    exp_41_ram[1512] = 35;
    exp_41_ram[1513] = 131;
    exp_41_ram[1514] = 3;
    exp_41_ram[1515] = 131;
    exp_41_ram[1516] = 3;
    exp_41_ram[1517] = 3;
    exp_41_ram[1518] = 131;
    exp_41_ram[1519] = 3;
    exp_41_ram[1520] = 131;
    exp_41_ram[1521] = 3;
    exp_41_ram[1522] = 131;
    exp_41_ram[1523] = 35;
    exp_41_ram[1524] = 35;
    exp_41_ram[1525] = 35;
    exp_41_ram[1526] = 35;
    exp_41_ram[1527] = 35;
    exp_41_ram[1528] = 35;
    exp_41_ram[1529] = 35;
    exp_41_ram[1530] = 35;
    exp_41_ram[1531] = 35;
    exp_41_ram[1532] = 3;
    exp_41_ram[1533] = 131;
    exp_41_ram[1534] = 3;
    exp_41_ram[1535] = 3;
    exp_41_ram[1536] = 131;
    exp_41_ram[1537] = 3;
    exp_41_ram[1538] = 131;
    exp_41_ram[1539] = 3;
    exp_41_ram[1540] = 131;
    exp_41_ram[1541] = 35;
    exp_41_ram[1542] = 35;
    exp_41_ram[1543] = 35;
    exp_41_ram[1544] = 35;
    exp_41_ram[1545] = 35;
    exp_41_ram[1546] = 35;
    exp_41_ram[1547] = 35;
    exp_41_ram[1548] = 35;
    exp_41_ram[1549] = 35;
    exp_41_ram[1550] = 147;
    exp_41_ram[1551] = 19;
    exp_41_ram[1552] = 239;
    exp_41_ram[1553] = 35;
    exp_41_ram[1554] = 35;
    exp_41_ram[1555] = 131;
    exp_41_ram[1556] = 99;
    exp_41_ram[1557] = 3;
    exp_41_ram[1558] = 131;
    exp_41_ram[1559] = 55;
    exp_41_ram[1560] = 19;
    exp_41_ram[1561] = 147;
    exp_41_ram[1562] = 51;
    exp_41_ram[1563] = 19;
    exp_41_ram[1564] = 51;
    exp_41_ram[1565] = 179;
    exp_41_ram[1566] = 179;
    exp_41_ram[1567] = 147;
    exp_41_ram[1568] = 35;
    exp_41_ram[1569] = 35;
    exp_41_ram[1570] = 111;
    exp_41_ram[1571] = 131;
    exp_41_ram[1572] = 99;
    exp_41_ram[1573] = 3;
    exp_41_ram[1574] = 131;
    exp_41_ram[1575] = 3;
    exp_41_ram[1576] = 3;
    exp_41_ram[1577] = 131;
    exp_41_ram[1578] = 3;
    exp_41_ram[1579] = 131;
    exp_41_ram[1580] = 3;
    exp_41_ram[1581] = 131;
    exp_41_ram[1582] = 35;
    exp_41_ram[1583] = 35;
    exp_41_ram[1584] = 35;
    exp_41_ram[1585] = 35;
    exp_41_ram[1586] = 35;
    exp_41_ram[1587] = 35;
    exp_41_ram[1588] = 35;
    exp_41_ram[1589] = 35;
    exp_41_ram[1590] = 35;
    exp_41_ram[1591] = 147;
    exp_41_ram[1592] = 19;
    exp_41_ram[1593] = 239;
    exp_41_ram[1594] = 147;
    exp_41_ram[1595] = 99;
    exp_41_ram[1596] = 55;
    exp_41_ram[1597] = 19;
    exp_41_ram[1598] = 147;
    exp_41_ram[1599] = 111;
    exp_41_ram[1600] = 19;
    exp_41_ram[1601] = 147;
    exp_41_ram[1602] = 3;
    exp_41_ram[1603] = 131;
    exp_41_ram[1604] = 51;
    exp_41_ram[1605] = 19;
    exp_41_ram[1606] = 51;
    exp_41_ram[1607] = 179;
    exp_41_ram[1608] = 179;
    exp_41_ram[1609] = 147;
    exp_41_ram[1610] = 35;
    exp_41_ram[1611] = 35;
    exp_41_ram[1612] = 111;
    exp_41_ram[1613] = 3;
    exp_41_ram[1614] = 131;
    exp_41_ram[1615] = 35;
    exp_41_ram[1616] = 35;
    exp_41_ram[1617] = 183;
    exp_41_ram[1618] = 131;
    exp_41_ram[1619] = 19;
    exp_41_ram[1620] = 147;
    exp_41_ram[1621] = 147;
    exp_41_ram[1622] = 3;
    exp_41_ram[1623] = 131;
    exp_41_ram[1624] = 51;
    exp_41_ram[1625] = 147;
    exp_41_ram[1626] = 179;
    exp_41_ram[1627] = 179;
    exp_41_ram[1628] = 179;
    exp_41_ram[1629] = 147;
    exp_41_ram[1630] = 35;
    exp_41_ram[1631] = 35;
    exp_41_ram[1632] = 131;
    exp_41_ram[1633] = 147;
    exp_41_ram[1634] = 131;
    exp_41_ram[1635] = 3;
    exp_41_ram[1636] = 19;
    exp_41_ram[1637] = 239;
    exp_41_ram[1638] = 3;
    exp_41_ram[1639] = 131;
    exp_41_ram[1640] = 3;
    exp_41_ram[1641] = 3;
    exp_41_ram[1642] = 131;
    exp_41_ram[1643] = 3;
    exp_41_ram[1644] = 131;
    exp_41_ram[1645] = 3;
    exp_41_ram[1646] = 131;
    exp_41_ram[1647] = 35;
    exp_41_ram[1648] = 35;
    exp_41_ram[1649] = 35;
    exp_41_ram[1650] = 35;
    exp_41_ram[1651] = 35;
    exp_41_ram[1652] = 35;
    exp_41_ram[1653] = 35;
    exp_41_ram[1654] = 35;
    exp_41_ram[1655] = 35;
    exp_41_ram[1656] = 131;
    exp_41_ram[1657] = 99;
    exp_41_ram[1658] = 131;
    exp_41_ram[1659] = 19;
    exp_41_ram[1660] = 35;
    exp_41_ram[1661] = 111;
    exp_41_ram[1662] = 131;
    exp_41_ram[1663] = 99;
    exp_41_ram[1664] = 3;
    exp_41_ram[1665] = 131;
    exp_41_ram[1666] = 3;
    exp_41_ram[1667] = 3;
    exp_41_ram[1668] = 131;
    exp_41_ram[1669] = 3;
    exp_41_ram[1670] = 131;
    exp_41_ram[1671] = 3;
    exp_41_ram[1672] = 131;
    exp_41_ram[1673] = 35;
    exp_41_ram[1674] = 35;
    exp_41_ram[1675] = 35;
    exp_41_ram[1676] = 35;
    exp_41_ram[1677] = 35;
    exp_41_ram[1678] = 35;
    exp_41_ram[1679] = 35;
    exp_41_ram[1680] = 35;
    exp_41_ram[1681] = 35;
    exp_41_ram[1682] = 147;
    exp_41_ram[1683] = 19;
    exp_41_ram[1684] = 239;
    exp_41_ram[1685] = 19;
    exp_41_ram[1686] = 131;
    exp_41_ram[1687] = 35;
    exp_41_ram[1688] = 111;
    exp_41_ram[1689] = 131;
    exp_41_ram[1690] = 35;
    exp_41_ram[1691] = 3;
    exp_41_ram[1692] = 131;
    exp_41_ram[1693] = 19;
    exp_41_ram[1694] = 147;
    exp_41_ram[1695] = 131;
    exp_41_ram[1696] = 3;
    exp_41_ram[1697] = 131;
    exp_41_ram[1698] = 3;
    exp_41_ram[1699] = 131;
    exp_41_ram[1700] = 19;
    exp_41_ram[1701] = 103;
    exp_41_ram[1702] = 19;
    exp_41_ram[1703] = 35;
    exp_41_ram[1704] = 35;
    exp_41_ram[1705] = 35;
    exp_41_ram[1706] = 35;
    exp_41_ram[1707] = 35;
    exp_41_ram[1708] = 35;
    exp_41_ram[1709] = 35;
    exp_41_ram[1710] = 35;
    exp_41_ram[1711] = 19;
    exp_41_ram[1712] = 35;
    exp_41_ram[1713] = 239;
    exp_41_ram[1714] = 19;
    exp_41_ram[1715] = 147;
    exp_41_ram[1716] = 183;
    exp_41_ram[1717] = 131;
    exp_41_ram[1718] = 19;
    exp_41_ram[1719] = 147;
    exp_41_ram[1720] = 19;
    exp_41_ram[1721] = 147;
    exp_41_ram[1722] = 19;
    exp_41_ram[1723] = 147;
    exp_41_ram[1724] = 239;
    exp_41_ram[1725] = 19;
    exp_41_ram[1726] = 147;
    exp_41_ram[1727] = 35;
    exp_41_ram[1728] = 183;
    exp_41_ram[1729] = 3;
    exp_41_ram[1730] = 131;
    exp_41_ram[1731] = 131;
    exp_41_ram[1732] = 179;
    exp_41_ram[1733] = 35;
    exp_41_ram[1734] = 131;
    exp_41_ram[1735] = 99;
    exp_41_ram[1736] = 131;
    exp_41_ram[1737] = 19;
    exp_41_ram[1738] = 147;
    exp_41_ram[1739] = 131;
    exp_41_ram[1740] = 35;
    exp_41_ram[1741] = 35;
    exp_41_ram[1742] = 131;
    exp_41_ram[1743] = 19;
    exp_41_ram[1744] = 147;
    exp_41_ram[1745] = 19;
    exp_41_ram[1746] = 147;
    exp_41_ram[1747] = 19;
    exp_41_ram[1748] = 147;
    exp_41_ram[1749] = 131;
    exp_41_ram[1750] = 3;
    exp_41_ram[1751] = 3;
    exp_41_ram[1752] = 131;
    exp_41_ram[1753] = 3;
    exp_41_ram[1754] = 131;
    exp_41_ram[1755] = 3;
    exp_41_ram[1756] = 131;
    exp_41_ram[1757] = 19;
    exp_41_ram[1758] = 103;
    exp_41_ram[1759] = 19;
    exp_41_ram[1760] = 35;
    exp_41_ram[1761] = 35;
    exp_41_ram[1762] = 35;
    exp_41_ram[1763] = 35;
    exp_41_ram[1764] = 19;
    exp_41_ram[1765] = 35;
    exp_41_ram[1766] = 35;
    exp_41_ram[1767] = 239;
    exp_41_ram[1768] = 19;
    exp_41_ram[1769] = 147;
    exp_41_ram[1770] = 183;
    exp_41_ram[1771] = 131;
    exp_41_ram[1772] = 19;
    exp_41_ram[1773] = 147;
    exp_41_ram[1774] = 19;
    exp_41_ram[1775] = 147;
    exp_41_ram[1776] = 19;
    exp_41_ram[1777] = 147;
    exp_41_ram[1778] = 239;
    exp_41_ram[1779] = 19;
    exp_41_ram[1780] = 147;
    exp_41_ram[1781] = 35;
    exp_41_ram[1782] = 35;
    exp_41_ram[1783] = 3;
    exp_41_ram[1784] = 131;
    exp_41_ram[1785] = 3;
    exp_41_ram[1786] = 131;
    exp_41_ram[1787] = 51;
    exp_41_ram[1788] = 19;
    exp_41_ram[1789] = 51;
    exp_41_ram[1790] = 179;
    exp_41_ram[1791] = 179;
    exp_41_ram[1792] = 147;
    exp_41_ram[1793] = 19;
    exp_41_ram[1794] = 147;
    exp_41_ram[1795] = 183;
    exp_41_ram[1796] = 35;
    exp_41_ram[1797] = 35;
    exp_41_ram[1798] = 19;
    exp_41_ram[1799] = 131;
    exp_41_ram[1800] = 3;
    exp_41_ram[1801] = 3;
    exp_41_ram[1802] = 131;
    exp_41_ram[1803] = 19;
    exp_41_ram[1804] = 103;
    exp_41_ram[1805] = 19;
    exp_41_ram[1806] = 35;
    exp_41_ram[1807] = 35;
    exp_41_ram[1808] = 19;
    exp_41_ram[1809] = 35;
    exp_41_ram[1810] = 183;
    exp_41_ram[1811] = 147;
    exp_41_ram[1812] = 3;
    exp_41_ram[1813] = 131;
    exp_41_ram[1814] = 3;
    exp_41_ram[1815] = 131;
    exp_41_ram[1816] = 3;
    exp_41_ram[1817] = 35;
    exp_41_ram[1818] = 35;
    exp_41_ram[1819] = 35;
    exp_41_ram[1820] = 35;
    exp_41_ram[1821] = 35;
    exp_41_ram[1822] = 131;
    exp_41_ram[1823] = 35;
    exp_41_ram[1824] = 183;
    exp_41_ram[1825] = 147;
    exp_41_ram[1826] = 3;
    exp_41_ram[1827] = 3;
    exp_41_ram[1828] = 131;
    exp_41_ram[1829] = 3;
    exp_41_ram[1830] = 3;
    exp_41_ram[1831] = 131;
    exp_41_ram[1832] = 3;
    exp_41_ram[1833] = 131;
    exp_41_ram[1834] = 3;
    exp_41_ram[1835] = 35;
    exp_41_ram[1836] = 35;
    exp_41_ram[1837] = 35;
    exp_41_ram[1838] = 35;
    exp_41_ram[1839] = 35;
    exp_41_ram[1840] = 35;
    exp_41_ram[1841] = 35;
    exp_41_ram[1842] = 35;
    exp_41_ram[1843] = 35;
    exp_41_ram[1844] = 131;
    exp_41_ram[1845] = 35;
    exp_41_ram[1846] = 35;
    exp_41_ram[1847] = 111;
    exp_41_ram[1848] = 131;
    exp_41_ram[1849] = 3;
    exp_41_ram[1850] = 147;
    exp_41_ram[1851] = 147;
    exp_41_ram[1852] = 51;
    exp_41_ram[1853] = 131;
    exp_41_ram[1854] = 179;
    exp_41_ram[1855] = 19;
    exp_41_ram[1856] = 179;
    exp_41_ram[1857] = 3;
    exp_41_ram[1858] = 183;
    exp_41_ram[1859] = 147;
    exp_41_ram[1860] = 131;
    exp_41_ram[1861] = 179;
    exp_41_ram[1862] = 35;
    exp_41_ram[1863] = 131;
    exp_41_ram[1864] = 147;
    exp_41_ram[1865] = 35;
    exp_41_ram[1866] = 3;
    exp_41_ram[1867] = 147;
    exp_41_ram[1868] = 227;
    exp_41_ram[1869] = 183;
    exp_41_ram[1870] = 147;
    exp_41_ram[1871] = 19;
    exp_41_ram[1872] = 163;
    exp_41_ram[1873] = 35;
    exp_41_ram[1874] = 111;
    exp_41_ram[1875] = 131;
    exp_41_ram[1876] = 3;
    exp_41_ram[1877] = 147;
    exp_41_ram[1878] = 147;
    exp_41_ram[1879] = 51;
    exp_41_ram[1880] = 131;
    exp_41_ram[1881] = 51;
    exp_41_ram[1882] = 131;
    exp_41_ram[1883] = 147;
    exp_41_ram[1884] = 147;
    exp_41_ram[1885] = 51;
    exp_41_ram[1886] = 3;
    exp_41_ram[1887] = 183;
    exp_41_ram[1888] = 147;
    exp_41_ram[1889] = 179;
    exp_41_ram[1890] = 35;
    exp_41_ram[1891] = 131;
    exp_41_ram[1892] = 147;
    exp_41_ram[1893] = 35;
    exp_41_ram[1894] = 3;
    exp_41_ram[1895] = 147;
    exp_41_ram[1896] = 227;
    exp_41_ram[1897] = 183;
    exp_41_ram[1898] = 147;
    exp_41_ram[1899] = 19;
    exp_41_ram[1900] = 163;
    exp_41_ram[1901] = 131;
    exp_41_ram[1902] = 131;
    exp_41_ram[1903] = 147;
    exp_41_ram[1904] = 19;
    exp_41_ram[1905] = 239;
    exp_41_ram[1906] = 19;
    exp_41_ram[1907] = 147;
    exp_41_ram[1908] = 35;
    exp_41_ram[1909] = 35;
    exp_41_ram[1910] = 131;
    exp_41_ram[1911] = 147;
    exp_41_ram[1912] = 147;
    exp_41_ram[1913] = 19;
    exp_41_ram[1914] = 183;
    exp_41_ram[1915] = 147;
    exp_41_ram[1916] = 35;
    exp_41_ram[1917] = 131;
    exp_41_ram[1918] = 147;
    exp_41_ram[1919] = 147;
    exp_41_ram[1920] = 19;
    exp_41_ram[1921] = 183;
    exp_41_ram[1922] = 147;
    exp_41_ram[1923] = 163;
    exp_41_ram[1924] = 183;
    exp_41_ram[1925] = 147;
    exp_41_ram[1926] = 19;
    exp_41_ram[1927] = 35;
    exp_41_ram[1928] = 131;
    exp_41_ram[1929] = 131;
    exp_41_ram[1930] = 147;
    exp_41_ram[1931] = 19;
    exp_41_ram[1932] = 239;
    exp_41_ram[1933] = 19;
    exp_41_ram[1934] = 147;
    exp_41_ram[1935] = 35;
    exp_41_ram[1936] = 35;
    exp_41_ram[1937] = 131;
    exp_41_ram[1938] = 147;
    exp_41_ram[1939] = 147;
    exp_41_ram[1940] = 19;
    exp_41_ram[1941] = 183;
    exp_41_ram[1942] = 147;
    exp_41_ram[1943] = 163;
    exp_41_ram[1944] = 131;
    exp_41_ram[1945] = 147;
    exp_41_ram[1946] = 147;
    exp_41_ram[1947] = 19;
    exp_41_ram[1948] = 183;
    exp_41_ram[1949] = 147;
    exp_41_ram[1950] = 35;
    exp_41_ram[1951] = 183;
    exp_41_ram[1952] = 147;
    exp_41_ram[1953] = 19;
    exp_41_ram[1954] = 163;
    exp_41_ram[1955] = 131;
    exp_41_ram[1956] = 131;
    exp_41_ram[1957] = 147;
    exp_41_ram[1958] = 19;
    exp_41_ram[1959] = 239;
    exp_41_ram[1960] = 19;
    exp_41_ram[1961] = 147;
    exp_41_ram[1962] = 35;
    exp_41_ram[1963] = 35;
    exp_41_ram[1964] = 131;
    exp_41_ram[1965] = 147;
    exp_41_ram[1966] = 147;
    exp_41_ram[1967] = 19;
    exp_41_ram[1968] = 183;
    exp_41_ram[1969] = 147;
    exp_41_ram[1970] = 35;
    exp_41_ram[1971] = 131;
    exp_41_ram[1972] = 147;
    exp_41_ram[1973] = 147;
    exp_41_ram[1974] = 19;
    exp_41_ram[1975] = 183;
    exp_41_ram[1976] = 147;
    exp_41_ram[1977] = 163;
    exp_41_ram[1978] = 183;
    exp_41_ram[1979] = 147;
    exp_41_ram[1980] = 19;
    exp_41_ram[1981] = 35;
    exp_41_ram[1982] = 131;
    exp_41_ram[1983] = 131;
    exp_41_ram[1984] = 147;
    exp_41_ram[1985] = 19;
    exp_41_ram[1986] = 239;
    exp_41_ram[1987] = 19;
    exp_41_ram[1988] = 147;
    exp_41_ram[1989] = 35;
    exp_41_ram[1990] = 35;
    exp_41_ram[1991] = 131;
    exp_41_ram[1992] = 147;
    exp_41_ram[1993] = 147;
    exp_41_ram[1994] = 19;
    exp_41_ram[1995] = 183;
    exp_41_ram[1996] = 147;
    exp_41_ram[1997] = 163;
    exp_41_ram[1998] = 131;
    exp_41_ram[1999] = 147;
    exp_41_ram[2000] = 147;
    exp_41_ram[2001] = 19;
    exp_41_ram[2002] = 183;
    exp_41_ram[2003] = 147;
    exp_41_ram[2004] = 35;
    exp_41_ram[2005] = 183;
    exp_41_ram[2006] = 147;
    exp_41_ram[2007] = 19;
    exp_41_ram[2008] = 163;
    exp_41_ram[2009] = 131;
    exp_41_ram[2010] = 131;
    exp_41_ram[2011] = 147;
    exp_41_ram[2012] = 147;
    exp_41_ram[2013] = 19;
    exp_41_ram[2014] = 239;
    exp_41_ram[2015] = 19;
    exp_41_ram[2016] = 147;
    exp_41_ram[2017] = 35;
    exp_41_ram[2018] = 35;
    exp_41_ram[2019] = 131;
    exp_41_ram[2020] = 147;
    exp_41_ram[2021] = 147;
    exp_41_ram[2022] = 19;
    exp_41_ram[2023] = 183;
    exp_41_ram[2024] = 147;
    exp_41_ram[2025] = 35;
    exp_41_ram[2026] = 131;
    exp_41_ram[2027] = 147;
    exp_41_ram[2028] = 19;
    exp_41_ram[2029] = 239;
    exp_41_ram[2030] = 19;
    exp_41_ram[2031] = 147;
    exp_41_ram[2032] = 35;
    exp_41_ram[2033] = 35;
    exp_41_ram[2034] = 131;
    exp_41_ram[2035] = 147;
    exp_41_ram[2036] = 147;
    exp_41_ram[2037] = 19;
    exp_41_ram[2038] = 183;
    exp_41_ram[2039] = 147;
    exp_41_ram[2040] = 163;
    exp_41_ram[2041] = 131;
    exp_41_ram[2042] = 147;
    exp_41_ram[2043] = 19;
    exp_41_ram[2044] = 239;
    exp_41_ram[2045] = 19;
    exp_41_ram[2046] = 147;
    exp_41_ram[2047] = 35;
    exp_41_ram[2048] = 35;
    exp_41_ram[2049] = 131;
    exp_41_ram[2050] = 147;
    exp_41_ram[2051] = 147;
    exp_41_ram[2052] = 19;
    exp_41_ram[2053] = 183;
    exp_41_ram[2054] = 147;
    exp_41_ram[2055] = 35;
    exp_41_ram[2056] = 131;
    exp_41_ram[2057] = 147;
    exp_41_ram[2058] = 147;
    exp_41_ram[2059] = 19;
    exp_41_ram[2060] = 183;
    exp_41_ram[2061] = 147;
    exp_41_ram[2062] = 163;
    exp_41_ram[2063] = 183;
    exp_41_ram[2064] = 147;
    exp_41_ram[2065] = 19;
    exp_41_ram[2066] = 35;
    exp_41_ram[2067] = 183;
    exp_41_ram[2068] = 147;
    exp_41_ram[2069] = 163;
    exp_41_ram[2070] = 183;
    exp_41_ram[2071] = 147;
    exp_41_ram[2072] = 19;
    exp_41_ram[2073] = 131;
    exp_41_ram[2074] = 3;
    exp_41_ram[2075] = 19;
    exp_41_ram[2076] = 103;
    exp_41_ram[2077] = 19;
    exp_41_ram[2078] = 35;
    exp_41_ram[2079] = 35;
    exp_41_ram[2080] = 19;
    exp_41_ram[2081] = 35;
    exp_41_ram[2082] = 3;
    exp_41_ram[2083] = 239;
    exp_41_ram[2084] = 147;
    exp_41_ram[2085] = 19;
    exp_41_ram[2086] = 239;
    exp_41_ram[2087] = 147;
    exp_41_ram[2088] = 19;
    exp_41_ram[2089] = 131;
    exp_41_ram[2090] = 3;
    exp_41_ram[2091] = 19;
    exp_41_ram[2092] = 103;
    exp_41_ram[2093] = 19;
    exp_41_ram[2094] = 35;
    exp_41_ram[2095] = 35;
    exp_41_ram[2096] = 35;
    exp_41_ram[2097] = 35;
    exp_41_ram[2098] = 35;
    exp_41_ram[2099] = 35;
    exp_41_ram[2100] = 35;
    exp_41_ram[2101] = 35;
    exp_41_ram[2102] = 35;
    exp_41_ram[2103] = 35;
    exp_41_ram[2104] = 19;
    exp_41_ram[2105] = 35;
    exp_41_ram[2106] = 35;
    exp_41_ram[2107] = 35;
    exp_41_ram[2108] = 147;
    exp_41_ram[2109] = 35;
    exp_41_ram[2110] = 147;
    exp_41_ram[2111] = 35;
    exp_41_ram[2112] = 131;
    exp_41_ram[2113] = 19;
    exp_41_ram[2114] = 239;
    exp_41_ram[2115] = 35;
    exp_41_ram[2116] = 3;
    exp_41_ram[2117] = 183;
    exp_41_ram[2118] = 147;
    exp_41_ram[2119] = 179;
    exp_41_ram[2120] = 35;
    exp_41_ram[2121] = 131;
    exp_41_ram[2122] = 19;
    exp_41_ram[2123] = 147;
    exp_41_ram[2124] = 131;
    exp_41_ram[2125] = 19;
    exp_41_ram[2126] = 99;
    exp_41_ram[2127] = 131;
    exp_41_ram[2128] = 19;
    exp_41_ram[2129] = 99;
    exp_41_ram[2130] = 131;
    exp_41_ram[2131] = 19;
    exp_41_ram[2132] = 99;
    exp_41_ram[2133] = 131;
    exp_41_ram[2134] = 147;
    exp_41_ram[2135] = 35;
    exp_41_ram[2136] = 131;
    exp_41_ram[2137] = 19;
    exp_41_ram[2138] = 131;
    exp_41_ram[2139] = 179;
    exp_41_ram[2140] = 35;
    exp_41_ram[2141] = 131;
    exp_41_ram[2142] = 19;
    exp_41_ram[2143] = 147;
    exp_41_ram[2144] = 3;
    exp_41_ram[2145] = 131;
    exp_41_ram[2146] = 51;
    exp_41_ram[2147] = 147;
    exp_41_ram[2148] = 179;
    exp_41_ram[2149] = 179;
    exp_41_ram[2150] = 179;
    exp_41_ram[2151] = 147;
    exp_41_ram[2152] = 35;
    exp_41_ram[2153] = 35;
    exp_41_ram[2154] = 111;
    exp_41_ram[2155] = 19;
    exp_41_ram[2156] = 35;
    exp_41_ram[2157] = 35;
    exp_41_ram[2158] = 131;
    exp_41_ram[2159] = 19;
    exp_41_ram[2160] = 131;
    exp_41_ram[2161] = 147;
    exp_41_ram[2162] = 19;
    exp_41_ram[2163] = 239;
    exp_41_ram[2164] = 35;
    exp_41_ram[2165] = 3;
    exp_41_ram[2166] = 183;
    exp_41_ram[2167] = 147;
    exp_41_ram[2168] = 179;
    exp_41_ram[2169] = 35;
    exp_41_ram[2170] = 131;
    exp_41_ram[2171] = 19;
    exp_41_ram[2172] = 147;
    exp_41_ram[2173] = 131;
    exp_41_ram[2174] = 19;
    exp_41_ram[2175] = 99;
    exp_41_ram[2176] = 131;
    exp_41_ram[2177] = 19;
    exp_41_ram[2178] = 99;
    exp_41_ram[2179] = 131;
    exp_41_ram[2180] = 19;
    exp_41_ram[2181] = 99;
    exp_41_ram[2182] = 131;
    exp_41_ram[2183] = 147;
    exp_41_ram[2184] = 35;
    exp_41_ram[2185] = 131;
    exp_41_ram[2186] = 19;
    exp_41_ram[2187] = 131;
    exp_41_ram[2188] = 179;
    exp_41_ram[2189] = 35;
    exp_41_ram[2190] = 131;
    exp_41_ram[2191] = 19;
    exp_41_ram[2192] = 131;
    exp_41_ram[2193] = 179;
    exp_41_ram[2194] = 35;
    exp_41_ram[2195] = 131;
    exp_41_ram[2196] = 19;
    exp_41_ram[2197] = 147;
    exp_41_ram[2198] = 3;
    exp_41_ram[2199] = 131;
    exp_41_ram[2200] = 51;
    exp_41_ram[2201] = 147;
    exp_41_ram[2202] = 179;
    exp_41_ram[2203] = 179;
    exp_41_ram[2204] = 179;
    exp_41_ram[2205] = 147;
    exp_41_ram[2206] = 35;
    exp_41_ram[2207] = 35;
    exp_41_ram[2208] = 111;
    exp_41_ram[2209] = 19;
    exp_41_ram[2210] = 131;
    exp_41_ram[2211] = 147;
    exp_41_ram[2212] = 35;
    exp_41_ram[2213] = 3;
    exp_41_ram[2214] = 183;
    exp_41_ram[2215] = 147;
    exp_41_ram[2216] = 19;
    exp_41_ram[2217] = 239;
    exp_41_ram[2218] = 19;
    exp_41_ram[2219] = 147;
    exp_41_ram[2220] = 35;
    exp_41_ram[2221] = 35;
    exp_41_ram[2222] = 131;
    exp_41_ram[2223] = 147;
    exp_41_ram[2224] = 35;
    exp_41_ram[2225] = 3;
    exp_41_ram[2226] = 131;
    exp_41_ram[2227] = 179;
    exp_41_ram[2228] = 35;
    exp_41_ram[2229] = 3;
    exp_41_ram[2230] = 147;
    exp_41_ram[2231] = 179;
    exp_41_ram[2232] = 35;
    exp_41_ram[2233] = 3;
    exp_41_ram[2234] = 131;
    exp_41_ram[2235] = 179;
    exp_41_ram[2236] = 35;
    exp_41_ram[2237] = 131;
    exp_41_ram[2238] = 35;
    exp_41_ram[2239] = 147;
    exp_41_ram[2240] = 35;
    exp_41_ram[2241] = 3;
    exp_41_ram[2242] = 183;
    exp_41_ram[2243] = 147;
    exp_41_ram[2244] = 19;
    exp_41_ram[2245] = 239;
    exp_41_ram[2246] = 19;
    exp_41_ram[2247] = 147;
    exp_41_ram[2248] = 35;
    exp_41_ram[2249] = 35;
    exp_41_ram[2250] = 131;
    exp_41_ram[2251] = 35;
    exp_41_ram[2252] = 131;
    exp_41_ram[2253] = 35;
    exp_41_ram[2254] = 147;
    exp_41_ram[2255] = 35;
    exp_41_ram[2256] = 131;
    exp_41_ram[2257] = 147;
    exp_41_ram[2258] = 19;
    exp_41_ram[2259] = 239;
    exp_41_ram[2260] = 19;
    exp_41_ram[2261] = 147;
    exp_41_ram[2262] = 35;
    exp_41_ram[2263] = 35;
    exp_41_ram[2264] = 131;
    exp_41_ram[2265] = 35;
    exp_41_ram[2266] = 131;
    exp_41_ram[2267] = 35;
    exp_41_ram[2268] = 147;
    exp_41_ram[2269] = 35;
    exp_41_ram[2270] = 131;
    exp_41_ram[2271] = 35;
    exp_41_ram[2272] = 131;
    exp_41_ram[2273] = 3;
    exp_41_ram[2274] = 3;
    exp_41_ram[2275] = 131;
    exp_41_ram[2276] = 3;
    exp_41_ram[2277] = 3;
    exp_41_ram[2278] = 131;
    exp_41_ram[2279] = 3;
    exp_41_ram[2280] = 131;
    exp_41_ram[2281] = 3;
    exp_41_ram[2282] = 35;
    exp_41_ram[2283] = 35;
    exp_41_ram[2284] = 35;
    exp_41_ram[2285] = 35;
    exp_41_ram[2286] = 35;
    exp_41_ram[2287] = 35;
    exp_41_ram[2288] = 35;
    exp_41_ram[2289] = 35;
    exp_41_ram[2290] = 35;
    exp_41_ram[2291] = 3;
    exp_41_ram[2292] = 131;
    exp_41_ram[2293] = 3;
    exp_41_ram[2294] = 3;
    exp_41_ram[2295] = 131;
    exp_41_ram[2296] = 3;
    exp_41_ram[2297] = 131;
    exp_41_ram[2298] = 3;
    exp_41_ram[2299] = 131;
    exp_41_ram[2300] = 3;
    exp_41_ram[2301] = 131;
    exp_41_ram[2302] = 19;
    exp_41_ram[2303] = 103;
    exp_41_ram[2304] = 19;
    exp_41_ram[2305] = 35;
    exp_41_ram[2306] = 35;
    exp_41_ram[2307] = 35;
    exp_41_ram[2308] = 35;
    exp_41_ram[2309] = 35;
    exp_41_ram[2310] = 19;
    exp_41_ram[2311] = 35;
    exp_41_ram[2312] = 147;
    exp_41_ram[2313] = 19;
    exp_41_ram[2314] = 35;
    exp_41_ram[2315] = 35;
    exp_41_ram[2316] = 131;
    exp_41_ram[2317] = 3;
    exp_41_ram[2318] = 131;
    exp_41_ram[2319] = 35;
    exp_41_ram[2320] = 35;
    exp_41_ram[2321] = 3;
    exp_41_ram[2322] = 131;
    exp_41_ram[2323] = 239;
    exp_41_ram[2324] = 147;
    exp_41_ram[2325] = 99;
    exp_41_ram[2326] = 55;
    exp_41_ram[2327] = 19;
    exp_41_ram[2328] = 147;
    exp_41_ram[2329] = 35;
    exp_41_ram[2330] = 35;
    exp_41_ram[2331] = 183;
    exp_41_ram[2332] = 131;
    exp_41_ram[2333] = 19;
    exp_41_ram[2334] = 147;
    exp_41_ram[2335] = 147;
    exp_41_ram[2336] = 3;
    exp_41_ram[2337] = 131;
    exp_41_ram[2338] = 51;
    exp_41_ram[2339] = 147;
    exp_41_ram[2340] = 179;
    exp_41_ram[2341] = 179;
    exp_41_ram[2342] = 179;
    exp_41_ram[2343] = 147;
    exp_41_ram[2344] = 19;
    exp_41_ram[2345] = 147;
    exp_41_ram[2346] = 3;
    exp_41_ram[2347] = 131;
    exp_41_ram[2348] = 51;
    exp_41_ram[2349] = 19;
    exp_41_ram[2350] = 51;
    exp_41_ram[2351] = 179;
    exp_41_ram[2352] = 179;
    exp_41_ram[2353] = 147;
    exp_41_ram[2354] = 35;
    exp_41_ram[2355] = 35;
    exp_41_ram[2356] = 183;
    exp_41_ram[2357] = 147;
    exp_41_ram[2358] = 147;
    exp_41_ram[2359] = 131;
    exp_41_ram[2360] = 3;
    exp_41_ram[2361] = 19;
    exp_41_ram[2362] = 239;
    exp_41_ram[2363] = 3;
    exp_41_ram[2364] = 131;
    exp_41_ram[2365] = 3;
    exp_41_ram[2366] = 3;
    exp_41_ram[2367] = 131;
    exp_41_ram[2368] = 3;
    exp_41_ram[2369] = 131;
    exp_41_ram[2370] = 3;
    exp_41_ram[2371] = 131;
    exp_41_ram[2372] = 35;
    exp_41_ram[2373] = 35;
    exp_41_ram[2374] = 35;
    exp_41_ram[2375] = 35;
    exp_41_ram[2376] = 35;
    exp_41_ram[2377] = 35;
    exp_41_ram[2378] = 35;
    exp_41_ram[2379] = 35;
    exp_41_ram[2380] = 35;
    exp_41_ram[2381] = 3;
    exp_41_ram[2382] = 131;
    exp_41_ram[2383] = 239;
    exp_41_ram[2384] = 19;
    exp_41_ram[2385] = 183;
    exp_41_ram[2386] = 147;
    exp_41_ram[2387] = 35;
    exp_41_ram[2388] = 183;
    exp_41_ram[2389] = 147;
    exp_41_ram[2390] = 19;
    exp_41_ram[2391] = 131;
    exp_41_ram[2392] = 3;
    exp_41_ram[2393] = 131;
    exp_41_ram[2394] = 3;
    exp_41_ram[2395] = 131;
    exp_41_ram[2396] = 19;
    exp_41_ram[2397] = 103;
    exp_41_ram[2398] = 19;
    exp_41_ram[2399] = 35;
    exp_41_ram[2400] = 35;
    exp_41_ram[2401] = 19;
    exp_41_ram[2402] = 35;
    exp_41_ram[2403] = 35;
    exp_41_ram[2404] = 3;
    exp_41_ram[2405] = 239;
    exp_41_ram[2406] = 147;
    exp_41_ram[2407] = 163;
    exp_41_ram[2408] = 131;
    exp_41_ram[2409] = 19;
    exp_41_ram[2410] = 147;
    exp_41_ram[2411] = 99;
    exp_41_ram[2412] = 3;
    exp_41_ram[2413] = 147;
    exp_41_ram[2414] = 147;
    exp_41_ram[2415] = 179;
    exp_41_ram[2416] = 147;
    exp_41_ram[2417] = 35;
    exp_41_ram[2418] = 3;
    exp_41_ram[2419] = 131;
    exp_41_ram[2420] = 179;
    exp_41_ram[2421] = 147;
    exp_41_ram[2422] = 35;
    exp_41_ram[2423] = 111;
    exp_41_ram[2424] = 19;
    exp_41_ram[2425] = 131;
    exp_41_ram[2426] = 19;
    exp_41_ram[2427] = 131;
    exp_41_ram[2428] = 3;
    exp_41_ram[2429] = 19;
    exp_41_ram[2430] = 103;
    exp_41_ram[2431] = 19;
    exp_41_ram[2432] = 35;
    exp_41_ram[2433] = 35;
    exp_41_ram[2434] = 19;
    exp_41_ram[2435] = 183;
    exp_41_ram[2436] = 131;
    exp_41_ram[2437] = 19;
    exp_41_ram[2438] = 239;
    exp_41_ram[2439] = 147;
    exp_41_ram[2440] = 19;
    exp_41_ram[2441] = 131;
    exp_41_ram[2442] = 3;
    exp_41_ram[2443] = 19;
    exp_41_ram[2444] = 103;
    exp_41_ram[2445] = 19;
    exp_41_ram[2446] = 35;
    exp_41_ram[2447] = 35;
    exp_41_ram[2448] = 19;
    exp_41_ram[2449] = 35;
    exp_41_ram[2450] = 35;
    exp_41_ram[2451] = 35;
    exp_41_ram[2452] = 183;
    exp_41_ram[2453] = 147;
    exp_41_ram[2454] = 35;
    exp_41_ram[2455] = 147;
    exp_41_ram[2456] = 35;
    exp_41_ram[2457] = 35;
    exp_41_ram[2458] = 111;
    exp_41_ram[2459] = 3;
    exp_41_ram[2460] = 131;
    exp_41_ram[2461] = 179;
    exp_41_ram[2462] = 163;
    exp_41_ram[2463] = 131;
    exp_41_ram[2464] = 99;
    exp_41_ram[2465] = 131;
    exp_41_ram[2466] = 99;
    exp_41_ram[2467] = 3;
    exp_41_ram[2468] = 147;
    exp_41_ram[2469] = 99;
    exp_41_ram[2470] = 131;
    exp_41_ram[2471] = 147;
    exp_41_ram[2472] = 131;
    exp_41_ram[2473] = 19;
    exp_41_ram[2474] = 239;
    exp_41_ram[2475] = 147;
    exp_41_ram[2476] = 35;
    exp_41_ram[2477] = 111;
    exp_41_ram[2478] = 131;
    exp_41_ram[2479] = 3;
    exp_41_ram[2480] = 99;
    exp_41_ram[2481] = 131;
    exp_41_ram[2482] = 147;
    exp_41_ram[2483] = 131;
    exp_41_ram[2484] = 19;
    exp_41_ram[2485] = 239;
    exp_41_ram[2486] = 3;
    exp_41_ram[2487] = 131;
    exp_41_ram[2488] = 179;
    exp_41_ram[2489] = 35;
    exp_41_ram[2490] = 3;
    exp_41_ram[2491] = 147;
    exp_41_ram[2492] = 179;
    exp_41_ram[2493] = 35;
    exp_41_ram[2494] = 131;
    exp_41_ram[2495] = 147;
    exp_41_ram[2496] = 35;
    exp_41_ram[2497] = 131;
    exp_41_ram[2498] = 227;
    exp_41_ram[2499] = 19;
    exp_41_ram[2500] = 19;
    exp_41_ram[2501] = 131;
    exp_41_ram[2502] = 3;
    exp_41_ram[2503] = 19;
    exp_41_ram[2504] = 103;
    exp_41_ram[2505] = 19;
    exp_41_ram[2506] = 35;
    exp_41_ram[2507] = 35;
    exp_41_ram[2508] = 19;
    exp_41_ram[2509] = 35;
    exp_41_ram[2510] = 35;
    exp_41_ram[2511] = 3;
    exp_41_ram[2512] = 131;
    exp_41_ram[2513] = 183;
    exp_41_ram[2514] = 131;
    exp_41_ram[2515] = 19;
    exp_41_ram[2516] = 147;
    exp_41_ram[2517] = 19;
    exp_41_ram[2518] = 239;
    exp_41_ram[2519] = 19;
    exp_41_ram[2520] = 131;
    exp_41_ram[2521] = 3;
    exp_41_ram[2522] = 19;
    exp_41_ram[2523] = 103;
    exp_41_ram[2524] = 19;
    exp_41_ram[2525] = 35;
    exp_41_ram[2526] = 35;
    exp_41_ram[2527] = 35;
    exp_41_ram[2528] = 35;
    exp_41_ram[2529] = 19;
    exp_41_ram[2530] = 35;
    exp_41_ram[2531] = 239;
    exp_41_ram[2532] = 35;
    exp_41_ram[2533] = 35;
    exp_41_ram[2534] = 19;
    exp_41_ram[2535] = 239;
    exp_41_ram[2536] = 19;
    exp_41_ram[2537] = 147;
    exp_41_ram[2538] = 3;
    exp_41_ram[2539] = 131;
    exp_41_ram[2540] = 51;
    exp_41_ram[2541] = 19;
    exp_41_ram[2542] = 51;
    exp_41_ram[2543] = 179;
    exp_41_ram[2544] = 179;
    exp_41_ram[2545] = 147;
    exp_41_ram[2546] = 131;
    exp_41_ram[2547] = 19;
    exp_41_ram[2548] = 147;
    exp_41_ram[2549] = 19;
    exp_41_ram[2550] = 147;
    exp_41_ram[2551] = 227;
    exp_41_ram[2552] = 19;
    exp_41_ram[2553] = 147;
    exp_41_ram[2554] = 99;
    exp_41_ram[2555] = 147;
    exp_41_ram[2556] = 147;
    exp_41_ram[2557] = 227;
    exp_41_ram[2558] = 19;
    exp_41_ram[2559] = 19;
    exp_41_ram[2560] = 131;
    exp_41_ram[2561] = 3;
    exp_41_ram[2562] = 3;
    exp_41_ram[2563] = 131;
    exp_41_ram[2564] = 19;
    exp_41_ram[2565] = 103;
    exp_41_ram[2566] = 19;
    exp_41_ram[2567] = 35;
    exp_41_ram[2568] = 35;
    exp_41_ram[2569] = 19;
    exp_41_ram[2570] = 183;
    exp_41_ram[2571] = 19;
    exp_41_ram[2572] = 239;
    exp_41_ram[2573] = 19;
    exp_41_ram[2574] = 131;
    exp_41_ram[2575] = 3;
    exp_41_ram[2576] = 19;
    exp_41_ram[2577] = 103;
    exp_41_ram[2578] = 19;
    exp_41_ram[2579] = 35;
    exp_41_ram[2580] = 35;
    exp_41_ram[2581] = 19;
    exp_41_ram[2582] = 183;
    exp_41_ram[2583] = 19;
    exp_41_ram[2584] = 239;
    exp_41_ram[2585] = 147;
    exp_41_ram[2586] = 35;
    exp_41_ram[2587] = 35;
    exp_41_ram[2588] = 111;
    exp_41_ram[2589] = 147;
    exp_41_ram[2590] = 3;
    exp_41_ram[2591] = 239;
    exp_41_ram[2592] = 19;
    exp_41_ram[2593] = 239;
    exp_41_ram[2594] = 111;
    exp_41_ram[2595] = 131;
    exp_41_ram[2596] = 147;
    exp_41_ram[2597] = 35;
    exp_41_ram[2598] = 183;
    exp_41_ram[2599] = 131;
    exp_41_ram[2600] = 147;
    exp_41_ram[2601] = 3;
    exp_41_ram[2602] = 239;
    exp_41_ram[2603] = 183;
    exp_41_ram[2604] = 3;
    exp_41_ram[2605] = 147;
    exp_41_ram[2606] = 179;
    exp_41_ram[2607] = 19;
    exp_41_ram[2608] = 239;
    exp_41_ram[2609] = 3;
    exp_41_ram[2610] = 147;
    exp_41_ram[2611] = 227;
    exp_41_ram[2612] = 111;
    exp_41_ram[2613] = 131;
    exp_41_ram[2614] = 147;
    exp_41_ram[2615] = 35;
    exp_41_ram[2616] = 183;
    exp_41_ram[2617] = 131;
    exp_41_ram[2618] = 147;
    exp_41_ram[2619] = 3;
    exp_41_ram[2620] = 239;
    exp_41_ram[2621] = 183;
    exp_41_ram[2622] = 3;
    exp_41_ram[2623] = 147;
    exp_41_ram[2624] = 179;
    exp_41_ram[2625] = 19;
    exp_41_ram[2626] = 239;
    exp_41_ram[2627] = 3;
    exp_41_ram[2628] = 147;
    exp_41_ram[2629] = 227;
    exp_41_ram[2630] = 131;
    exp_41_ram[2631] = 147;
    exp_41_ram[2632] = 35;
    exp_41_ram[2633] = 3;
    exp_41_ram[2634] = 147;
    exp_41_ram[2635] = 227;
    exp_41_ram[2636] = 183;
    exp_41_ram[2637] = 131;
    exp_41_ram[2638] = 147;
    exp_41_ram[2639] = 19;
    exp_41_ram[2640] = 239;
    exp_41_ram[2641] = 19;
    exp_41_ram[2642] = 131;
    exp_41_ram[2643] = 3;
    exp_41_ram[2644] = 19;
    exp_41_ram[2645] = 103;
    exp_41_ram[2646] = 19;
    exp_41_ram[2647] = 35;
    exp_41_ram[2648] = 35;
    exp_41_ram[2649] = 19;
    exp_41_ram[2650] = 183;
    exp_41_ram[2651] = 19;
    exp_41_ram[2652] = 239;
    exp_41_ram[2653] = 35;
    exp_41_ram[2654] = 111;
    exp_41_ram[2655] = 147;
    exp_41_ram[2656] = 3;
    exp_41_ram[2657] = 239;
    exp_41_ram[2658] = 19;
    exp_41_ram[2659] = 239;
    exp_41_ram[2660] = 35;
    exp_41_ram[2661] = 111;
    exp_41_ram[2662] = 183;
    exp_41_ram[2663] = 131;
    exp_41_ram[2664] = 147;
    exp_41_ram[2665] = 3;
    exp_41_ram[2666] = 239;
    exp_41_ram[2667] = 183;
    exp_41_ram[2668] = 3;
    exp_41_ram[2669] = 147;
    exp_41_ram[2670] = 179;
    exp_41_ram[2671] = 19;
    exp_41_ram[2672] = 239;
    exp_41_ram[2673] = 131;
    exp_41_ram[2674] = 147;
    exp_41_ram[2675] = 35;
    exp_41_ram[2676] = 3;
    exp_41_ram[2677] = 147;
    exp_41_ram[2678] = 227;
    exp_41_ram[2679] = 147;
    exp_41_ram[2680] = 35;
    exp_41_ram[2681] = 111;
    exp_41_ram[2682] = 183;
    exp_41_ram[2683] = 131;
    exp_41_ram[2684] = 147;
    exp_41_ram[2685] = 3;
    exp_41_ram[2686] = 239;
    exp_41_ram[2687] = 183;
    exp_41_ram[2688] = 3;
    exp_41_ram[2689] = 147;
    exp_41_ram[2690] = 179;
    exp_41_ram[2691] = 19;
    exp_41_ram[2692] = 239;
    exp_41_ram[2693] = 131;
    exp_41_ram[2694] = 147;
    exp_41_ram[2695] = 35;
    exp_41_ram[2696] = 131;
    exp_41_ram[2697] = 227;
    exp_41_ram[2698] = 131;
    exp_41_ram[2699] = 147;
    exp_41_ram[2700] = 35;
    exp_41_ram[2701] = 3;
    exp_41_ram[2702] = 147;
    exp_41_ram[2703] = 227;
    exp_41_ram[2704] = 183;
    exp_41_ram[2705] = 131;
    exp_41_ram[2706] = 147;
    exp_41_ram[2707] = 19;
    exp_41_ram[2708] = 239;
    exp_41_ram[2709] = 19;
    exp_41_ram[2710] = 131;
    exp_41_ram[2711] = 3;
    exp_41_ram[2712] = 19;
    exp_41_ram[2713] = 103;
    exp_41_ram[2714] = 19;
    exp_41_ram[2715] = 35;
    exp_41_ram[2716] = 35;
    exp_41_ram[2717] = 35;
    exp_41_ram[2718] = 35;
    exp_41_ram[2719] = 35;
    exp_41_ram[2720] = 35;
    exp_41_ram[2721] = 35;
    exp_41_ram[2722] = 35;
    exp_41_ram[2723] = 35;
    exp_41_ram[2724] = 35;
    exp_41_ram[2725] = 35;
    exp_41_ram[2726] = 35;
    exp_41_ram[2727] = 19;
    exp_41_ram[2728] = 147;
    exp_41_ram[2729] = 35;
    exp_41_ram[2730] = 19;
    exp_41_ram[2731] = 147;
    exp_41_ram[2732] = 35;
    exp_41_ram[2733] = 35;
    exp_41_ram[2734] = 239;
    exp_41_ram[2735] = 35;
    exp_41_ram[2736] = 35;
    exp_41_ram[2737] = 35;
    exp_41_ram[2738] = 111;
    exp_41_ram[2739] = 3;
    exp_41_ram[2740] = 183;
    exp_41_ram[2741] = 147;
    exp_41_ram[2742] = 179;
    exp_41_ram[2743] = 35;
    exp_41_ram[2744] = 3;
    exp_41_ram[2745] = 183;
    exp_41_ram[2746] = 147;
    exp_41_ram[2747] = 179;
    exp_41_ram[2748] = 35;
    exp_41_ram[2749] = 3;
    exp_41_ram[2750] = 183;
    exp_41_ram[2751] = 147;
    exp_41_ram[2752] = 179;
    exp_41_ram[2753] = 35;
    exp_41_ram[2754] = 3;
    exp_41_ram[2755] = 183;
    exp_41_ram[2756] = 147;
    exp_41_ram[2757] = 179;
    exp_41_ram[2758] = 35;
    exp_41_ram[2759] = 131;
    exp_41_ram[2760] = 147;
    exp_41_ram[2761] = 35;
    exp_41_ram[2762] = 239;
    exp_41_ram[2763] = 19;
    exp_41_ram[2764] = 147;
    exp_41_ram[2765] = 3;
    exp_41_ram[2766] = 131;
    exp_41_ram[2767] = 51;
    exp_41_ram[2768] = 19;
    exp_41_ram[2769] = 51;
    exp_41_ram[2770] = 179;
    exp_41_ram[2771] = 179;
    exp_41_ram[2772] = 147;
    exp_41_ram[2773] = 183;
    exp_41_ram[2774] = 131;
    exp_41_ram[2775] = 35;
    exp_41_ram[2776] = 35;
    exp_41_ram[2777] = 3;
    exp_41_ram[2778] = 131;
    exp_41_ram[2779] = 19;
    exp_41_ram[2780] = 147;
    exp_41_ram[2781] = 227;
    exp_41_ram[2782] = 19;
    exp_41_ram[2783] = 147;
    exp_41_ram[2784] = 99;
    exp_41_ram[2785] = 147;
    exp_41_ram[2786] = 147;
    exp_41_ram[2787] = 227;
    exp_41_ram[2788] = 131;
    exp_41_ram[2789] = 147;
    exp_41_ram[2790] = 19;
    exp_41_ram[2791] = 239;
    exp_41_ram[2792] = 183;
    exp_41_ram[2793] = 19;
    exp_41_ram[2794] = 239;
    exp_41_ram[2795] = 239;
    exp_41_ram[2796] = 35;
    exp_41_ram[2797] = 35;
    exp_41_ram[2798] = 35;
    exp_41_ram[2799] = 111;
    exp_41_ram[2800] = 3;
    exp_41_ram[2801] = 131;
    exp_41_ram[2802] = 183;
    exp_41_ram[2803] = 147;
    exp_41_ram[2804] = 51;
    exp_41_ram[2805] = 147;
    exp_41_ram[2806] = 179;
    exp_41_ram[2807] = 51;
    exp_41_ram[2808] = 183;
    exp_41_ram[2809] = 147;
    exp_41_ram[2810] = 179;
    exp_41_ram[2811] = 179;
    exp_41_ram[2812] = 19;
    exp_41_ram[2813] = 179;
    exp_41_ram[2814] = 147;
    exp_41_ram[2815] = 35;
    exp_41_ram[2816] = 35;
    exp_41_ram[2817] = 3;
    exp_41_ram[2818] = 131;
    exp_41_ram[2819] = 183;
    exp_41_ram[2820] = 147;
    exp_41_ram[2821] = 51;
    exp_41_ram[2822] = 147;
    exp_41_ram[2823] = 179;
    exp_41_ram[2824] = 51;
    exp_41_ram[2825] = 183;
    exp_41_ram[2826] = 147;
    exp_41_ram[2827] = 179;
    exp_41_ram[2828] = 179;
    exp_41_ram[2829] = 19;
    exp_41_ram[2830] = 179;
    exp_41_ram[2831] = 147;
    exp_41_ram[2832] = 35;
    exp_41_ram[2833] = 35;
    exp_41_ram[2834] = 3;
    exp_41_ram[2835] = 131;
    exp_41_ram[2836] = 183;
    exp_41_ram[2837] = 147;
    exp_41_ram[2838] = 51;
    exp_41_ram[2839] = 147;
    exp_41_ram[2840] = 179;
    exp_41_ram[2841] = 51;
    exp_41_ram[2842] = 183;
    exp_41_ram[2843] = 147;
    exp_41_ram[2844] = 179;
    exp_41_ram[2845] = 179;
    exp_41_ram[2846] = 19;
    exp_41_ram[2847] = 179;
    exp_41_ram[2848] = 147;
    exp_41_ram[2849] = 35;
    exp_41_ram[2850] = 35;
    exp_41_ram[2851] = 3;
    exp_41_ram[2852] = 131;
    exp_41_ram[2853] = 183;
    exp_41_ram[2854] = 147;
    exp_41_ram[2855] = 51;
    exp_41_ram[2856] = 147;
    exp_41_ram[2857] = 179;
    exp_41_ram[2858] = 51;
    exp_41_ram[2859] = 183;
    exp_41_ram[2860] = 147;
    exp_41_ram[2861] = 179;
    exp_41_ram[2862] = 179;
    exp_41_ram[2863] = 19;
    exp_41_ram[2864] = 179;
    exp_41_ram[2865] = 147;
    exp_41_ram[2866] = 35;
    exp_41_ram[2867] = 35;
    exp_41_ram[2868] = 131;
    exp_41_ram[2869] = 147;
    exp_41_ram[2870] = 35;
    exp_41_ram[2871] = 239;
    exp_41_ram[2872] = 19;
    exp_41_ram[2873] = 147;
    exp_41_ram[2874] = 3;
    exp_41_ram[2875] = 131;
    exp_41_ram[2876] = 51;
    exp_41_ram[2877] = 19;
    exp_41_ram[2878] = 51;
    exp_41_ram[2879] = 179;
    exp_41_ram[2880] = 179;
    exp_41_ram[2881] = 147;
    exp_41_ram[2882] = 183;
    exp_41_ram[2883] = 131;
    exp_41_ram[2884] = 35;
    exp_41_ram[2885] = 35;
    exp_41_ram[2886] = 3;
    exp_41_ram[2887] = 131;
    exp_41_ram[2888] = 19;
    exp_41_ram[2889] = 147;
    exp_41_ram[2890] = 227;
    exp_41_ram[2891] = 19;
    exp_41_ram[2892] = 147;
    exp_41_ram[2893] = 99;
    exp_41_ram[2894] = 147;
    exp_41_ram[2895] = 147;
    exp_41_ram[2896] = 227;
    exp_41_ram[2897] = 131;
    exp_41_ram[2898] = 147;
    exp_41_ram[2899] = 19;
    exp_41_ram[2900] = 239;
    exp_41_ram[2901] = 183;
    exp_41_ram[2902] = 19;
    exp_41_ram[2903] = 239;
    exp_41_ram[2904] = 239;
    exp_41_ram[2905] = 35;
    exp_41_ram[2906] = 35;
    exp_41_ram[2907] = 35;
    exp_41_ram[2908] = 111;
    exp_41_ram[2909] = 3;
    exp_41_ram[2910] = 183;
    exp_41_ram[2911] = 147;
    exp_41_ram[2912] = 179;
    exp_41_ram[2913] = 35;
    exp_41_ram[2914] = 3;
    exp_41_ram[2915] = 183;
    exp_41_ram[2916] = 147;
    exp_41_ram[2917] = 179;
    exp_41_ram[2918] = 35;
    exp_41_ram[2919] = 3;
    exp_41_ram[2920] = 183;
    exp_41_ram[2921] = 147;
    exp_41_ram[2922] = 179;
    exp_41_ram[2923] = 35;
    exp_41_ram[2924] = 3;
    exp_41_ram[2925] = 183;
    exp_41_ram[2926] = 147;
    exp_41_ram[2927] = 179;
    exp_41_ram[2928] = 35;
    exp_41_ram[2929] = 131;
    exp_41_ram[2930] = 147;
    exp_41_ram[2931] = 35;
    exp_41_ram[2932] = 239;
    exp_41_ram[2933] = 19;
    exp_41_ram[2934] = 147;
    exp_41_ram[2935] = 3;
    exp_41_ram[2936] = 131;
    exp_41_ram[2937] = 51;
    exp_41_ram[2938] = 19;
    exp_41_ram[2939] = 51;
    exp_41_ram[2940] = 179;
    exp_41_ram[2941] = 179;
    exp_41_ram[2942] = 147;
    exp_41_ram[2943] = 183;
    exp_41_ram[2944] = 131;
    exp_41_ram[2945] = 35;
    exp_41_ram[2946] = 35;
    exp_41_ram[2947] = 3;
    exp_41_ram[2948] = 131;
    exp_41_ram[2949] = 19;
    exp_41_ram[2950] = 147;
    exp_41_ram[2951] = 227;
    exp_41_ram[2952] = 19;
    exp_41_ram[2953] = 147;
    exp_41_ram[2954] = 99;
    exp_41_ram[2955] = 147;
    exp_41_ram[2956] = 147;
    exp_41_ram[2957] = 227;
    exp_41_ram[2958] = 131;
    exp_41_ram[2959] = 147;
    exp_41_ram[2960] = 19;
    exp_41_ram[2961] = 239;
    exp_41_ram[2962] = 183;
    exp_41_ram[2963] = 19;
    exp_41_ram[2964] = 239;
    exp_41_ram[2965] = 239;
    exp_41_ram[2966] = 35;
    exp_41_ram[2967] = 35;
    exp_41_ram[2968] = 35;
    exp_41_ram[2969] = 111;
    exp_41_ram[2970] = 3;
    exp_41_ram[2971] = 131;
    exp_41_ram[2972] = 55;
    exp_41_ram[2973] = 19;
    exp_41_ram[2974] = 147;
    exp_41_ram[2975] = 19;
    exp_41_ram[2976] = 147;
    exp_41_ram[2977] = 239;
    exp_41_ram[2978] = 19;
    exp_41_ram[2979] = 147;
    exp_41_ram[2980] = 35;
    exp_41_ram[2981] = 35;
    exp_41_ram[2982] = 3;
    exp_41_ram[2983] = 131;
    exp_41_ram[2984] = 55;
    exp_41_ram[2985] = 19;
    exp_41_ram[2986] = 147;
    exp_41_ram[2987] = 19;
    exp_41_ram[2988] = 147;
    exp_41_ram[2989] = 239;
    exp_41_ram[2990] = 19;
    exp_41_ram[2991] = 147;
    exp_41_ram[2992] = 35;
    exp_41_ram[2993] = 35;
    exp_41_ram[2994] = 3;
    exp_41_ram[2995] = 131;
    exp_41_ram[2996] = 55;
    exp_41_ram[2997] = 19;
    exp_41_ram[2998] = 147;
    exp_41_ram[2999] = 19;
    exp_41_ram[3000] = 147;
    exp_41_ram[3001] = 239;
    exp_41_ram[3002] = 19;
    exp_41_ram[3003] = 147;
    exp_41_ram[3004] = 35;
    exp_41_ram[3005] = 35;
    exp_41_ram[3006] = 3;
    exp_41_ram[3007] = 131;
    exp_41_ram[3008] = 55;
    exp_41_ram[3009] = 19;
    exp_41_ram[3010] = 147;
    exp_41_ram[3011] = 19;
    exp_41_ram[3012] = 147;
    exp_41_ram[3013] = 239;
    exp_41_ram[3014] = 19;
    exp_41_ram[3015] = 147;
    exp_41_ram[3016] = 35;
    exp_41_ram[3017] = 35;
    exp_41_ram[3018] = 131;
    exp_41_ram[3019] = 147;
    exp_41_ram[3020] = 35;
    exp_41_ram[3021] = 239;
    exp_41_ram[3022] = 19;
    exp_41_ram[3023] = 147;
    exp_41_ram[3024] = 3;
    exp_41_ram[3025] = 131;
    exp_41_ram[3026] = 51;
    exp_41_ram[3027] = 19;
    exp_41_ram[3028] = 51;
    exp_41_ram[3029] = 179;
    exp_41_ram[3030] = 179;
    exp_41_ram[3031] = 147;
    exp_41_ram[3032] = 183;
    exp_41_ram[3033] = 131;
    exp_41_ram[3034] = 19;
    exp_41_ram[3035] = 147;
    exp_41_ram[3036] = 19;
    exp_41_ram[3037] = 147;
    exp_41_ram[3038] = 227;
    exp_41_ram[3039] = 19;
    exp_41_ram[3040] = 147;
    exp_41_ram[3041] = 99;
    exp_41_ram[3042] = 147;
    exp_41_ram[3043] = 147;
    exp_41_ram[3044] = 227;
    exp_41_ram[3045] = 131;
    exp_41_ram[3046] = 147;
    exp_41_ram[3047] = 19;
    exp_41_ram[3048] = 239;
    exp_41_ram[3049] = 183;
    exp_41_ram[3050] = 19;
    exp_41_ram[3051] = 239;
    exp_41_ram[3052] = 19;
    exp_41_ram[3053] = 131;
    exp_41_ram[3054] = 3;
    exp_41_ram[3055] = 3;
    exp_41_ram[3056] = 131;
    exp_41_ram[3057] = 3;
    exp_41_ram[3058] = 131;
    exp_41_ram[3059] = 3;
    exp_41_ram[3060] = 131;
    exp_41_ram[3061] = 3;
    exp_41_ram[3062] = 131;
    exp_41_ram[3063] = 3;
    exp_41_ram[3064] = 131;
    exp_41_ram[3065] = 19;
    exp_41_ram[3066] = 103;
    exp_41_ram[3067] = 19;
    exp_41_ram[3068] = 35;
    exp_41_ram[3069] = 35;
    exp_41_ram[3070] = 35;
    exp_41_ram[3071] = 35;
    exp_41_ram[3072] = 35;
    exp_41_ram[3073] = 35;
    exp_41_ram[3074] = 19;
    exp_41_ram[3075] = 183;
    exp_41_ram[3076] = 19;
    exp_41_ram[3077] = 239;
    exp_41_ram[3078] = 239;
    exp_41_ram[3079] = 147;
    exp_41_ram[3080] = 147;
    exp_41_ram[3081] = 35;
    exp_41_ram[3082] = 183;
    exp_41_ram[3083] = 19;
    exp_41_ram[3084] = 239;
    exp_41_ram[3085] = 239;
    exp_41_ram[3086] = 147;
    exp_41_ram[3087] = 147;
    exp_41_ram[3088] = 35;
    exp_41_ram[3089] = 183;
    exp_41_ram[3090] = 19;
    exp_41_ram[3091] = 239;
    exp_41_ram[3092] = 239;
    exp_41_ram[3093] = 147;
    exp_41_ram[3094] = 35;
    exp_41_ram[3095] = 183;
    exp_41_ram[3096] = 19;
    exp_41_ram[3097] = 239;
    exp_41_ram[3098] = 239;
    exp_41_ram[3099] = 147;
    exp_41_ram[3100] = 35;
    exp_41_ram[3101] = 183;
    exp_41_ram[3102] = 19;
    exp_41_ram[3103] = 239;
    exp_41_ram[3104] = 239;
    exp_41_ram[3105] = 147;
    exp_41_ram[3106] = 35;
    exp_41_ram[3107] = 147;
    exp_41_ram[3108] = 35;
    exp_41_ram[3109] = 147;
    exp_41_ram[3110] = 35;
    exp_41_ram[3111] = 147;
    exp_41_ram[3112] = 19;
    exp_41_ram[3113] = 239;
    exp_41_ram[3114] = 19;
    exp_41_ram[3115] = 147;
    exp_41_ram[3116] = 35;
    exp_41_ram[3117] = 35;
    exp_41_ram[3118] = 3;
    exp_41_ram[3119] = 131;
    exp_41_ram[3120] = 19;
    exp_41_ram[3121] = 147;
    exp_41_ram[3122] = 239;
    exp_41_ram[3123] = 239;
    exp_41_ram[3124] = 35;
    exp_41_ram[3125] = 35;
    exp_41_ram[3126] = 35;
    exp_41_ram[3127] = 111;
    exp_41_ram[3128] = 19;
    exp_41_ram[3129] = 239;
    exp_41_ram[3130] = 19;
    exp_41_ram[3131] = 147;
    exp_41_ram[3132] = 3;
    exp_41_ram[3133] = 131;
    exp_41_ram[3134] = 19;
    exp_41_ram[3135] = 147;
    exp_41_ram[3136] = 239;
    exp_41_ram[3137] = 19;
    exp_41_ram[3138] = 147;
    exp_41_ram[3139] = 183;
    exp_41_ram[3140] = 131;
    exp_41_ram[3141] = 19;
    exp_41_ram[3142] = 239;
    exp_41_ram[3143] = 19;
    exp_41_ram[3144] = 147;
    exp_41_ram[3145] = 19;
    exp_41_ram[3146] = 147;
    exp_41_ram[3147] = 19;
    exp_41_ram[3148] = 147;
    exp_41_ram[3149] = 239;
    exp_41_ram[3150] = 147;
    exp_41_ram[3151] = 227;
    exp_41_ram[3152] = 183;
    exp_41_ram[3153] = 131;
    exp_41_ram[3154] = 19;
    exp_41_ram[3155] = 147;
    exp_41_ram[3156] = 3;
    exp_41_ram[3157] = 131;
    exp_41_ram[3158] = 51;
    exp_41_ram[3159] = 147;
    exp_41_ram[3160] = 179;
    exp_41_ram[3161] = 179;
    exp_41_ram[3162] = 179;
    exp_41_ram[3163] = 147;
    exp_41_ram[3164] = 35;
    exp_41_ram[3165] = 35;
    exp_41_ram[3166] = 19;
    exp_41_ram[3167] = 239;
    exp_41_ram[3168] = 19;
    exp_41_ram[3169] = 147;
    exp_41_ram[3170] = 35;
    exp_41_ram[3171] = 35;
    exp_41_ram[3172] = 147;
    exp_41_ram[3173] = 19;
    exp_41_ram[3174] = 239;
    exp_41_ram[3175] = 147;
    exp_41_ram[3176] = 19;
    exp_41_ram[3177] = 239;
    exp_41_ram[3178] = 131;
    exp_41_ram[3179] = 147;
    exp_41_ram[3180] = 35;
    exp_41_ram[3181] = 3;
    exp_41_ram[3182] = 147;
    exp_41_ram[3183] = 227;
    exp_41_ram[3184] = 19;
    exp_41_ram[3185] = 19;
    exp_41_ram[3186] = 131;
    exp_41_ram[3187] = 3;
    exp_41_ram[3188] = 3;
    exp_41_ram[3189] = 131;
    exp_41_ram[3190] = 3;
    exp_41_ram[3191] = 131;
    exp_41_ram[3192] = 19;
    exp_41_ram[3193] = 103;
    exp_41_ram[3194] = 19;
    exp_41_ram[3195] = 35;
    exp_41_ram[3196] = 35;
    exp_41_ram[3197] = 19;
    exp_41_ram[3198] = 183;
    exp_41_ram[3199] = 19;
    exp_41_ram[3200] = 239;
    exp_41_ram[3201] = 183;
    exp_41_ram[3202] = 19;
    exp_41_ram[3203] = 239;
    exp_41_ram[3204] = 183;
    exp_41_ram[3205] = 19;
    exp_41_ram[3206] = 239;
    exp_41_ram[3207] = 183;
    exp_41_ram[3208] = 19;
    exp_41_ram[3209] = 239;
    exp_41_ram[3210] = 183;
    exp_41_ram[3211] = 19;
    exp_41_ram[3212] = 239;
    exp_41_ram[3213] = 183;
    exp_41_ram[3214] = 19;
    exp_41_ram[3215] = 239;
    exp_41_ram[3216] = 183;
    exp_41_ram[3217] = 19;
    exp_41_ram[3218] = 239;
    exp_41_ram[3219] = 239;
    exp_41_ram[3220] = 147;
    exp_41_ram[3221] = 163;
    exp_41_ram[3222] = 131;
    exp_41_ram[3223] = 147;
    exp_41_ram[3224] = 19;
    exp_41_ram[3225] = 227;
    exp_41_ram[3226] = 19;
    exp_41_ram[3227] = 183;
    exp_41_ram[3228] = 147;
    exp_41_ram[3229] = 179;
    exp_41_ram[3230] = 131;
    exp_41_ram[3231] = 103;
    exp_41_ram[3232] = 239;
    exp_41_ram[3233] = 111;
    exp_41_ram[3234] = 239;
    exp_41_ram[3235] = 111;
    exp_41_ram[3236] = 239;
    exp_41_ram[3237] = 111;
    exp_41_ram[3238] = 239;
    exp_41_ram[3239] = 111;
    exp_41_ram[3240] = 239;
    exp_41_ram[3241] = 111;
    exp_41_ram[3242] = 239;
    exp_41_ram[3243] = 19;
    exp_41_ram[3244] = 111;
    exp_41_ram[3245] = 19;
    exp_41_ram[3246] = 35;
    exp_41_ram[3247] = 19;
    exp_41_ram[3248] = 147;
    exp_41_ram[3249] = 163;
    exp_41_ram[3250] = 131;
    exp_41_ram[3251] = 19;
    exp_41_ram[3252] = 147;
    exp_41_ram[3253] = 179;
    exp_41_ram[3254] = 147;
    exp_41_ram[3255] = 19;
    exp_41_ram[3256] = 3;
    exp_41_ram[3257] = 19;
    exp_41_ram[3258] = 103;
    exp_41_ram[3259] = 19;
    exp_41_ram[3260] = 35;
    exp_41_ram[3261] = 35;
    exp_41_ram[3262] = 35;
    exp_41_ram[3263] = 19;
    exp_41_ram[3264] = 35;
    exp_41_ram[3265] = 35;
    exp_41_ram[3266] = 35;
    exp_41_ram[3267] = 35;
    exp_41_ram[3268] = 35;
    exp_41_ram[3269] = 147;
    exp_41_ram[3270] = 19;
    exp_41_ram[3271] = 163;
    exp_41_ram[3272] = 147;
    exp_41_ram[3273] = 35;
    exp_41_ram[3274] = 147;
    exp_41_ram[3275] = 163;
    exp_41_ram[3276] = 131;
    exp_41_ram[3277] = 147;
    exp_41_ram[3278] = 19;
    exp_41_ram[3279] = 131;
    exp_41_ram[3280] = 163;
    exp_41_ram[3281] = 131;
    exp_41_ram[3282] = 147;
    exp_41_ram[3283] = 19;
    exp_41_ram[3284] = 131;
    exp_41_ram[3285] = 35;
    exp_41_ram[3286] = 131;
    exp_41_ram[3287] = 147;
    exp_41_ram[3288] = 19;
    exp_41_ram[3289] = 131;
    exp_41_ram[3290] = 163;
    exp_41_ram[3291] = 131;
    exp_41_ram[3292] = 147;
    exp_41_ram[3293] = 131;
    exp_41_ram[3294] = 147;
    exp_41_ram[3295] = 19;
    exp_41_ram[3296] = 131;
    exp_41_ram[3297] = 163;
    exp_41_ram[3298] = 131;
    exp_41_ram[3299] = 147;
    exp_41_ram[3300] = 131;
    exp_41_ram[3301] = 147;
    exp_41_ram[3302] = 19;
    exp_41_ram[3303] = 131;
    exp_41_ram[3304] = 35;
    exp_41_ram[3305] = 131;
    exp_41_ram[3306] = 147;
    exp_41_ram[3307] = 19;
    exp_41_ram[3308] = 131;
    exp_41_ram[3309] = 35;
    exp_41_ram[3310] = 131;
    exp_41_ram[3311] = 147;
    exp_41_ram[3312] = 19;
    exp_41_ram[3313] = 131;
    exp_41_ram[3314] = 163;
    exp_41_ram[3315] = 131;
    exp_41_ram[3316] = 147;
    exp_41_ram[3317] = 19;
    exp_41_ram[3318] = 131;
    exp_41_ram[3319] = 35;
    exp_41_ram[3320] = 163;
    exp_41_ram[3321] = 111;
    exp_41_ram[3322] = 131;
    exp_41_ram[3323] = 3;
    exp_41_ram[3324] = 179;
    exp_41_ram[3325] = 131;
    exp_41_ram[3326] = 147;
    exp_41_ram[3327] = 35;
    exp_41_ram[3328] = 131;
    exp_41_ram[3329] = 3;
    exp_41_ram[3330] = 179;
    exp_41_ram[3331] = 131;
    exp_41_ram[3332] = 147;
    exp_41_ram[3333] = 163;
    exp_41_ram[3334] = 131;
    exp_41_ram[3335] = 3;
    exp_41_ram[3336] = 179;
    exp_41_ram[3337] = 131;
    exp_41_ram[3338] = 147;
    exp_41_ram[3339] = 35;
    exp_41_ram[3340] = 131;
    exp_41_ram[3341] = 3;
    exp_41_ram[3342] = 179;
    exp_41_ram[3343] = 131;
    exp_41_ram[3344] = 147;
    exp_41_ram[3345] = 163;
    exp_41_ram[3346] = 131;
    exp_41_ram[3347] = 19;
    exp_41_ram[3348] = 239;
    exp_41_ram[3349] = 147;
    exp_41_ram[3350] = 19;
    exp_41_ram[3351] = 131;
    exp_41_ram[3352] = 179;
    exp_41_ram[3353] = 3;
    exp_41_ram[3354] = 35;
    exp_41_ram[3355] = 131;
    exp_41_ram[3356] = 19;
    exp_41_ram[3357] = 239;
    exp_41_ram[3358] = 147;
    exp_41_ram[3359] = 19;
    exp_41_ram[3360] = 131;
    exp_41_ram[3361] = 179;
    exp_41_ram[3362] = 3;
    exp_41_ram[3363] = 35;
    exp_41_ram[3364] = 131;
    exp_41_ram[3365] = 19;
    exp_41_ram[3366] = 239;
    exp_41_ram[3367] = 147;
    exp_41_ram[3368] = 19;
    exp_41_ram[3369] = 131;
    exp_41_ram[3370] = 179;
    exp_41_ram[3371] = 3;
    exp_41_ram[3372] = 35;
    exp_41_ram[3373] = 131;
    exp_41_ram[3374] = 3;
    exp_41_ram[3375] = 179;
    exp_41_ram[3376] = 3;
    exp_41_ram[3377] = 35;
    exp_41_ram[3378] = 131;
    exp_41_ram[3379] = 131;
    exp_41_ram[3380] = 19;
    exp_41_ram[3381] = 239;
    exp_41_ram[3382] = 147;
    exp_41_ram[3383] = 19;
    exp_41_ram[3384] = 131;
    exp_41_ram[3385] = 179;
    exp_41_ram[3386] = 35;
    exp_41_ram[3387] = 131;
    exp_41_ram[3388] = 131;
    exp_41_ram[3389] = 19;
    exp_41_ram[3390] = 239;
    exp_41_ram[3391] = 147;
    exp_41_ram[3392] = 19;
    exp_41_ram[3393] = 131;
    exp_41_ram[3394] = 179;
    exp_41_ram[3395] = 35;
    exp_41_ram[3396] = 131;
    exp_41_ram[3397] = 131;
    exp_41_ram[3398] = 19;
    exp_41_ram[3399] = 239;
    exp_41_ram[3400] = 147;
    exp_41_ram[3401] = 19;
    exp_41_ram[3402] = 131;
    exp_41_ram[3403] = 179;
    exp_41_ram[3404] = 35;
    exp_41_ram[3405] = 131;
    exp_41_ram[3406] = 147;
    exp_41_ram[3407] = 163;
    exp_41_ram[3408] = 3;
    exp_41_ram[3409] = 147;
    exp_41_ram[3410] = 227;
    exp_41_ram[3411] = 19;
    exp_41_ram[3412] = 19;
    exp_41_ram[3413] = 131;
    exp_41_ram[3414] = 3;
    exp_41_ram[3415] = 131;
    exp_41_ram[3416] = 19;
    exp_41_ram[3417] = 103;
    exp_41_ram[3418] = 19;
    exp_41_ram[3419] = 35;
    exp_41_ram[3420] = 35;
    exp_41_ram[3421] = 19;
    exp_41_ram[3422] = 35;
    exp_41_ram[3423] = 147;
    exp_41_ram[3424] = 163;
    exp_41_ram[3425] = 131;
    exp_41_ram[3426] = 3;
    exp_41_ram[3427] = 131;
    exp_41_ram[3428] = 131;
    exp_41_ram[3429] = 99;
    exp_41_ram[3430] = 131;
    exp_41_ram[3431] = 131;
    exp_41_ram[3432] = 147;
    exp_41_ram[3433] = 147;
    exp_41_ram[3434] = 19;
    exp_41_ram[3435] = 239;
    exp_41_ram[3436] = 147;
    exp_41_ram[3437] = 19;
    exp_41_ram[3438] = 131;
    exp_41_ram[3439] = 163;
    exp_41_ram[3440] = 131;
    exp_41_ram[3441] = 3;
    exp_41_ram[3442] = 131;
    exp_41_ram[3443] = 131;
    exp_41_ram[3444] = 99;
    exp_41_ram[3445] = 131;
    exp_41_ram[3446] = 131;
    exp_41_ram[3447] = 147;
    exp_41_ram[3448] = 147;
    exp_41_ram[3449] = 19;
    exp_41_ram[3450] = 239;
    exp_41_ram[3451] = 147;
    exp_41_ram[3452] = 19;
    exp_41_ram[3453] = 131;
    exp_41_ram[3454] = 35;
    exp_41_ram[3455] = 131;
    exp_41_ram[3456] = 131;
    exp_41_ram[3457] = 147;
    exp_41_ram[3458] = 147;
    exp_41_ram[3459] = 19;
    exp_41_ram[3460] = 239;
    exp_41_ram[3461] = 147;
    exp_41_ram[3462] = 19;
    exp_41_ram[3463] = 131;
    exp_41_ram[3464] = 163;
    exp_41_ram[3465] = 131;
    exp_41_ram[3466] = 147;
    exp_41_ram[3467] = 163;
    exp_41_ram[3468] = 131;
    exp_41_ram[3469] = 3;
    exp_41_ram[3470] = 131;
    exp_41_ram[3471] = 179;
    exp_41_ram[3472] = 19;
    exp_41_ram[3473] = 131;
    exp_41_ram[3474] = 131;
    exp_41_ram[3475] = 179;
    exp_41_ram[3476] = 147;
    exp_41_ram[3477] = 19;
    exp_41_ram[3478] = 239;
    exp_41_ram[3479] = 147;
    exp_41_ram[3480] = 19;
    exp_41_ram[3481] = 131;
    exp_41_ram[3482] = 179;
    exp_41_ram[3483] = 3;
    exp_41_ram[3484] = 131;
    exp_41_ram[3485] = 131;
    exp_41_ram[3486] = 179;
    exp_41_ram[3487] = 19;
    exp_41_ram[3488] = 131;
    exp_41_ram[3489] = 131;
    exp_41_ram[3490] = 179;
    exp_41_ram[3491] = 147;
    exp_41_ram[3492] = 19;
    exp_41_ram[3493] = 239;
    exp_41_ram[3494] = 147;
    exp_41_ram[3495] = 163;
    exp_41_ram[3496] = 131;
    exp_41_ram[3497] = 3;
    exp_41_ram[3498] = 131;
    exp_41_ram[3499] = 179;
    exp_41_ram[3500] = 19;
    exp_41_ram[3501] = 131;
    exp_41_ram[3502] = 131;
    exp_41_ram[3503] = 179;
    exp_41_ram[3504] = 147;
    exp_41_ram[3505] = 19;
    exp_41_ram[3506] = 239;
    exp_41_ram[3507] = 147;
    exp_41_ram[3508] = 19;
    exp_41_ram[3509] = 131;
    exp_41_ram[3510] = 179;
    exp_41_ram[3511] = 3;
    exp_41_ram[3512] = 131;
    exp_41_ram[3513] = 131;
    exp_41_ram[3514] = 179;
    exp_41_ram[3515] = 19;
    exp_41_ram[3516] = 131;
    exp_41_ram[3517] = 131;
    exp_41_ram[3518] = 179;
    exp_41_ram[3519] = 147;
    exp_41_ram[3520] = 19;
    exp_41_ram[3521] = 239;
    exp_41_ram[3522] = 147;
    exp_41_ram[3523] = 163;
    exp_41_ram[3524] = 131;
    exp_41_ram[3525] = 3;
    exp_41_ram[3526] = 131;
    exp_41_ram[3527] = 179;
    exp_41_ram[3528] = 19;
    exp_41_ram[3529] = 131;
    exp_41_ram[3530] = 131;
    exp_41_ram[3531] = 179;
    exp_41_ram[3532] = 147;
    exp_41_ram[3533] = 19;
    exp_41_ram[3534] = 239;
    exp_41_ram[3535] = 147;
    exp_41_ram[3536] = 19;
    exp_41_ram[3537] = 131;
    exp_41_ram[3538] = 179;
    exp_41_ram[3539] = 3;
    exp_41_ram[3540] = 131;
    exp_41_ram[3541] = 131;
    exp_41_ram[3542] = 179;
    exp_41_ram[3543] = 19;
    exp_41_ram[3544] = 131;
    exp_41_ram[3545] = 131;
    exp_41_ram[3546] = 179;
    exp_41_ram[3547] = 147;
    exp_41_ram[3548] = 19;
    exp_41_ram[3549] = 239;
    exp_41_ram[3550] = 147;
    exp_41_ram[3551] = 163;
    exp_41_ram[3552] = 131;
    exp_41_ram[3553] = 3;
    exp_41_ram[3554] = 179;
    exp_41_ram[3555] = 131;
    exp_41_ram[3556] = 163;
    exp_41_ram[3557] = 131;
    exp_41_ram[3558] = 3;
    exp_41_ram[3559] = 131;
    exp_41_ram[3560] = 179;
    exp_41_ram[3561] = 19;
    exp_41_ram[3562] = 131;
    exp_41_ram[3563] = 131;
    exp_41_ram[3564] = 179;
    exp_41_ram[3565] = 147;
    exp_41_ram[3566] = 19;
    exp_41_ram[3567] = 239;
    exp_41_ram[3568] = 147;
    exp_41_ram[3569] = 19;
    exp_41_ram[3570] = 131;
    exp_41_ram[3571] = 179;
    exp_41_ram[3572] = 3;
    exp_41_ram[3573] = 131;
    exp_41_ram[3574] = 131;
    exp_41_ram[3575] = 179;
    exp_41_ram[3576] = 19;
    exp_41_ram[3577] = 131;
    exp_41_ram[3578] = 131;
    exp_41_ram[3579] = 179;
    exp_41_ram[3580] = 147;
    exp_41_ram[3581] = 19;
    exp_41_ram[3582] = 239;
    exp_41_ram[3583] = 147;
    exp_41_ram[3584] = 163;
    exp_41_ram[3585] = 131;
    exp_41_ram[3586] = 3;
    exp_41_ram[3587] = 131;
    exp_41_ram[3588] = 179;
    exp_41_ram[3589] = 19;
    exp_41_ram[3590] = 131;
    exp_41_ram[3591] = 131;
    exp_41_ram[3592] = 179;
    exp_41_ram[3593] = 147;
    exp_41_ram[3594] = 19;
    exp_41_ram[3595] = 239;
    exp_41_ram[3596] = 147;
    exp_41_ram[3597] = 19;
    exp_41_ram[3598] = 131;
    exp_41_ram[3599] = 179;
    exp_41_ram[3600] = 3;
    exp_41_ram[3601] = 131;
    exp_41_ram[3602] = 131;
    exp_41_ram[3603] = 179;
    exp_41_ram[3604] = 19;
    exp_41_ram[3605] = 131;
    exp_41_ram[3606] = 131;
    exp_41_ram[3607] = 179;
    exp_41_ram[3608] = 147;
    exp_41_ram[3609] = 19;
    exp_41_ram[3610] = 239;
    exp_41_ram[3611] = 147;
    exp_41_ram[3612] = 163;
    exp_41_ram[3613] = 131;
    exp_41_ram[3614] = 3;
    exp_41_ram[3615] = 131;
    exp_41_ram[3616] = 179;
    exp_41_ram[3617] = 19;
    exp_41_ram[3618] = 131;
    exp_41_ram[3619] = 131;
    exp_41_ram[3620] = 179;
    exp_41_ram[3621] = 147;
    exp_41_ram[3622] = 19;
    exp_41_ram[3623] = 239;
    exp_41_ram[3624] = 147;
    exp_41_ram[3625] = 19;
    exp_41_ram[3626] = 131;
    exp_41_ram[3627] = 179;
    exp_41_ram[3628] = 3;
    exp_41_ram[3629] = 131;
    exp_41_ram[3630] = 131;
    exp_41_ram[3631] = 179;
    exp_41_ram[3632] = 19;
    exp_41_ram[3633] = 131;
    exp_41_ram[3634] = 131;
    exp_41_ram[3635] = 179;
    exp_41_ram[3636] = 147;
    exp_41_ram[3637] = 19;
    exp_41_ram[3638] = 239;
    exp_41_ram[3639] = 147;
    exp_41_ram[3640] = 163;
    exp_41_ram[3641] = 131;
    exp_41_ram[3642] = 147;
    exp_41_ram[3643] = 147;
    exp_41_ram[3644] = 19;
    exp_41_ram[3645] = 131;
    exp_41_ram[3646] = 3;
    exp_41_ram[3647] = 19;
    exp_41_ram[3648] = 103;
    exp_41_ram[3649] = 19;
    exp_41_ram[3650] = 35;
    exp_41_ram[3651] = 35;
    exp_41_ram[3652] = 19;
    exp_41_ram[3653] = 239;
    exp_41_ram[3654] = 147;
    exp_41_ram[3655] = 163;
    exp_41_ram[3656] = 3;
    exp_41_ram[3657] = 147;
    exp_41_ram[3658] = 99;
    exp_41_ram[3659] = 183;
    exp_41_ram[3660] = 147;
    exp_41_ram[3661] = 111;
    exp_41_ram[3662] = 3;
    exp_41_ram[3663] = 147;
    exp_41_ram[3664] = 99;
    exp_41_ram[3665] = 183;
    exp_41_ram[3666] = 147;
    exp_41_ram[3667] = 111;
    exp_41_ram[3668] = 3;
    exp_41_ram[3669] = 147;
    exp_41_ram[3670] = 99;
    exp_41_ram[3671] = 183;
    exp_41_ram[3672] = 147;
    exp_41_ram[3673] = 111;
    exp_41_ram[3674] = 3;
    exp_41_ram[3675] = 147;
    exp_41_ram[3676] = 99;
    exp_41_ram[3677] = 183;
    exp_41_ram[3678] = 147;
    exp_41_ram[3679] = 111;
    exp_41_ram[3680] = 3;
    exp_41_ram[3681] = 147;
    exp_41_ram[3682] = 227;
    exp_41_ram[3683] = 183;
    exp_41_ram[3684] = 147;
    exp_41_ram[3685] = 19;
    exp_41_ram[3686] = 131;
    exp_41_ram[3687] = 3;
    exp_41_ram[3688] = 19;
    exp_41_ram[3689] = 103;
    exp_41_ram[3690] = 19;
    exp_41_ram[3691] = 35;
    exp_41_ram[3692] = 35;
    exp_41_ram[3693] = 19;
    exp_41_ram[3694] = 239;
    exp_41_ram[3695] = 147;
    exp_41_ram[3696] = 163;
    exp_41_ram[3697] = 131;
    exp_41_ram[3698] = 19;
    exp_41_ram[3699] = 239;
    exp_41_ram[3700] = 19;
    exp_41_ram[3701] = 147;
    exp_41_ram[3702] = 99;
    exp_41_ram[3703] = 183;
    exp_41_ram[3704] = 147;
    exp_41_ram[3705] = 111;
    exp_41_ram[3706] = 131;
    exp_41_ram[3707] = 19;
    exp_41_ram[3708] = 239;
    exp_41_ram[3709] = 19;
    exp_41_ram[3710] = 147;
    exp_41_ram[3711] = 99;
    exp_41_ram[3712] = 183;
    exp_41_ram[3713] = 147;
    exp_41_ram[3714] = 111;
    exp_41_ram[3715] = 131;
    exp_41_ram[3716] = 19;
    exp_41_ram[3717] = 239;
    exp_41_ram[3718] = 19;
    exp_41_ram[3719] = 147;
    exp_41_ram[3720] = 227;
    exp_41_ram[3721] = 183;
    exp_41_ram[3722] = 147;
    exp_41_ram[3723] = 19;
    exp_41_ram[3724] = 131;
    exp_41_ram[3725] = 3;
    exp_41_ram[3726] = 19;
    exp_41_ram[3727] = 103;
    exp_41_ram[3728] = 19;
    exp_41_ram[3729] = 35;
    exp_41_ram[3730] = 35;
    exp_41_ram[3731] = 19;
    exp_41_ram[3732] = 239;
    exp_41_ram[3733] = 147;
    exp_41_ram[3734] = 163;
    exp_41_ram[3735] = 131;
    exp_41_ram[3736] = 19;
    exp_41_ram[3737] = 239;
    exp_41_ram[3738] = 147;
    exp_41_ram[3739] = 227;
    exp_41_ram[3740] = 131;
    exp_41_ram[3741] = 19;
    exp_41_ram[3742] = 239;
    exp_41_ram[3743] = 147;
    exp_41_ram[3744] = 147;
    exp_41_ram[3745] = 19;
    exp_41_ram[3746] = 131;
    exp_41_ram[3747] = 3;
    exp_41_ram[3748] = 19;
    exp_41_ram[3749] = 103;
    exp_41_ram[3750] = 19;
    exp_41_ram[3751] = 35;
    exp_41_ram[3752] = 35;
    exp_41_ram[3753] = 19;
    exp_41_ram[3754] = 183;
    exp_41_ram[3755] = 131;
    exp_41_ram[3756] = 183;
    exp_41_ram[3757] = 3;
    exp_41_ram[3758] = 183;
    exp_41_ram[3759] = 3;
    exp_41_ram[3760] = 183;
    exp_41_ram[3761] = 3;
    exp_41_ram[3762] = 183;
    exp_41_ram[3763] = 3;
    exp_41_ram[3764] = 183;
    exp_41_ram[3765] = 3;
    exp_41_ram[3766] = 183;
    exp_41_ram[3767] = 131;
    exp_41_ram[3768] = 183;
    exp_41_ram[3769] = 131;
    exp_41_ram[3770] = 55;
    exp_41_ram[3771] = 3;
    exp_41_ram[3772] = 183;
    exp_41_ram[3773] = 131;
    exp_41_ram[3774] = 35;
    exp_41_ram[3775] = 35;
    exp_41_ram[3776] = 35;
    exp_41_ram[3777] = 147;
    exp_41_ram[3778] = 19;
    exp_41_ram[3779] = 147;
    exp_41_ram[3780] = 55;
    exp_41_ram[3781] = 19;
    exp_41_ram[3782] = 239;
    exp_41_ram[3783] = 183;
    exp_41_ram[3784] = 19;
    exp_41_ram[3785] = 239;
    exp_41_ram[3786] = 183;
    exp_41_ram[3787] = 131;
    exp_41_ram[3788] = 19;
    exp_41_ram[3789] = 239;
    exp_41_ram[3790] = 183;
    exp_41_ram[3791] = 131;
    exp_41_ram[3792] = 19;
    exp_41_ram[3793] = 239;
    exp_41_ram[3794] = 183;
    exp_41_ram[3795] = 131;
    exp_41_ram[3796] = 19;
    exp_41_ram[3797] = 239;
    exp_41_ram[3798] = 183;
    exp_41_ram[3799] = 19;
    exp_41_ram[3800] = 239;
    exp_41_ram[3801] = 19;
    exp_41_ram[3802] = 131;
    exp_41_ram[3803] = 3;
    exp_41_ram[3804] = 19;
    exp_41_ram[3805] = 103;
    exp_41_ram[3806] = 19;
    exp_41_ram[3807] = 35;
    exp_41_ram[3808] = 35;
    exp_41_ram[3809] = 19;
    exp_41_ram[3810] = 183;
    exp_41_ram[3811] = 55;
    exp_41_ram[3812] = 19;
    exp_41_ram[3813] = 35;
    exp_41_ram[3814] = 183;
    exp_41_ram[3815] = 55;
    exp_41_ram[3816] = 19;
    exp_41_ram[3817] = 35;
    exp_41_ram[3818] = 183;
    exp_41_ram[3819] = 55;
    exp_41_ram[3820] = 19;
    exp_41_ram[3821] = 35;
    exp_41_ram[3822] = 183;
    exp_41_ram[3823] = 55;
    exp_41_ram[3824] = 19;
    exp_41_ram[3825] = 35;
    exp_41_ram[3826] = 183;
    exp_41_ram[3827] = 19;
    exp_41_ram[3828] = 35;
    exp_41_ram[3829] = 183;
    exp_41_ram[3830] = 19;
    exp_41_ram[3831] = 163;
    exp_41_ram[3832] = 183;
    exp_41_ram[3833] = 19;
    exp_41_ram[3834] = 35;
    exp_41_ram[3835] = 183;
    exp_41_ram[3836] = 19;
    exp_41_ram[3837] = 163;
    exp_41_ram[3838] = 183;
    exp_41_ram[3839] = 19;
    exp_41_ram[3840] = 35;
    exp_41_ram[3841] = 183;
    exp_41_ram[3842] = 19;
    exp_41_ram[3843] = 163;
    exp_41_ram[3844] = 239;
    exp_41_ram[3845] = 183;
    exp_41_ram[3846] = 19;
    exp_41_ram[3847] = 239;
    exp_41_ram[3848] = 183;
    exp_41_ram[3849] = 19;
    exp_41_ram[3850] = 239;
    exp_41_ram[3851] = 183;
    exp_41_ram[3852] = 19;
    exp_41_ram[3853] = 239;
    exp_41_ram[3854] = 183;
    exp_41_ram[3855] = 19;
    exp_41_ram[3856] = 239;
    exp_41_ram[3857] = 183;
    exp_41_ram[3858] = 19;
    exp_41_ram[3859] = 239;
    exp_41_ram[3860] = 183;
    exp_41_ram[3861] = 19;
    exp_41_ram[3862] = 239;
    exp_41_ram[3863] = 183;
    exp_41_ram[3864] = 19;
    exp_41_ram[3865] = 239;
    exp_41_ram[3866] = 35;
    exp_41_ram[3867] = 239;
    exp_41_ram[3868] = 147;
    exp_41_ram[3869] = 163;
    exp_41_ram[3870] = 131;
    exp_41_ram[3871] = 19;
    exp_41_ram[3872] = 239;
    exp_41_ram[3873] = 147;
    exp_41_ram[3874] = 99;
    exp_41_ram[3875] = 131;
    exp_41_ram[3876] = 99;
    exp_41_ram[3877] = 183;
    exp_41_ram[3878] = 147;
    exp_41_ram[3879] = 131;
    exp_41_ram[3880] = 147;
    exp_41_ram[3881] = 19;
    exp_41_ram[3882] = 239;
    exp_41_ram[3883] = 183;
    exp_41_ram[3884] = 147;
    exp_41_ram[3885] = 131;
    exp_41_ram[3886] = 147;
    exp_41_ram[3887] = 19;
    exp_41_ram[3888] = 239;
    exp_41_ram[3889] = 183;
    exp_41_ram[3890] = 147;
    exp_41_ram[3891] = 131;
    exp_41_ram[3892] = 147;
    exp_41_ram[3893] = 19;
    exp_41_ram[3894] = 239;
    exp_41_ram[3895] = 183;
    exp_41_ram[3896] = 19;
    exp_41_ram[3897] = 239;
    exp_41_ram[3898] = 131;
    exp_41_ram[3899] = 19;
    exp_41_ram[3900] = 239;
    exp_41_ram[3901] = 147;
    exp_41_ram[3902] = 147;
    exp_41_ram[3903] = 147;
    exp_41_ram[3904] = 183;
    exp_41_ram[3905] = 19;
    exp_41_ram[3906] = 239;
    exp_41_ram[3907] = 147;
    exp_41_ram[3908] = 19;
    exp_41_ram[3909] = 239;
    exp_41_ram[3910] = 3;
    exp_41_ram[3911] = 147;
    exp_41_ram[3912] = 99;
    exp_41_ram[3913] = 35;
    exp_41_ram[3914] = 19;
    exp_41_ram[3915] = 239;
    exp_41_ram[3916] = 111;
    exp_41_ram[3917] = 131;
    exp_41_ram[3918] = 147;
    exp_41_ram[3919] = 35;
    exp_41_ram[3920] = 111;
    exp_41_ram[3921] = 131;
    exp_41_ram[3922] = 19;
    exp_41_ram[3923] = 147;
    exp_41_ram[3924] = 227;
    exp_41_ram[3925] = 3;
    exp_41_ram[3926] = 147;
    exp_41_ram[3927] = 99;
    exp_41_ram[3928] = 183;
    exp_41_ram[3929] = 19;
    exp_41_ram[3930] = 239;
    exp_41_ram[3931] = 239;
    exp_41_ram[3932] = 19;
    exp_41_ram[3933] = 183;
    exp_41_ram[3934] = 35;
    exp_41_ram[3935] = 239;
    exp_41_ram[3936] = 19;
    exp_41_ram[3937] = 183;
    exp_41_ram[3938] = 35;
    exp_41_ram[3939] = 239;
    exp_41_ram[3940] = 19;
    exp_41_ram[3941] = 183;
    exp_41_ram[3942] = 35;
    exp_41_ram[3943] = 239;
    exp_41_ram[3944] = 35;
    exp_41_ram[3945] = 111;
    exp_41_ram[3946] = 3;
    exp_41_ram[3947] = 147;
    exp_41_ram[3948] = 99;
    exp_41_ram[3949] = 183;
    exp_41_ram[3950] = 19;
    exp_41_ram[3951] = 239;
    exp_41_ram[3952] = 239;
    exp_41_ram[3953] = 19;
    exp_41_ram[3954] = 183;
    exp_41_ram[3955] = 35;
    exp_41_ram[3956] = 239;
    exp_41_ram[3957] = 35;
    exp_41_ram[3958] = 111;
    exp_41_ram[3959] = 3;
    exp_41_ram[3960] = 147;
    exp_41_ram[3961] = 99;
    exp_41_ram[3962] = 183;
    exp_41_ram[3963] = 19;
    exp_41_ram[3964] = 239;
    exp_41_ram[3965] = 239;
    exp_41_ram[3966] = 147;
    exp_41_ram[3967] = 19;
    exp_41_ram[3968] = 183;
    exp_41_ram[3969] = 35;
    exp_41_ram[3970] = 239;
    exp_41_ram[3971] = 147;
    exp_41_ram[3972] = 19;
    exp_41_ram[3973] = 183;
    exp_41_ram[3974] = 163;
    exp_41_ram[3975] = 239;
    exp_41_ram[3976] = 147;
    exp_41_ram[3977] = 19;
    exp_41_ram[3978] = 183;
    exp_41_ram[3979] = 35;
    exp_41_ram[3980] = 239;
    exp_41_ram[3981] = 35;
    exp_41_ram[3982] = 111;
    exp_41_ram[3983] = 3;
    exp_41_ram[3984] = 147;
    exp_41_ram[3985] = 227;
    exp_41_ram[3986] = 183;
    exp_41_ram[3987] = 19;
    exp_41_ram[3988] = 239;
    exp_41_ram[3989] = 239;
    exp_41_ram[3990] = 147;
    exp_41_ram[3991] = 19;
    exp_41_ram[3992] = 183;
    exp_41_ram[3993] = 163;
    exp_41_ram[3994] = 239;
    exp_41_ram[3995] = 147;
    exp_41_ram[3996] = 19;
    exp_41_ram[3997] = 183;
    exp_41_ram[3998] = 35;
    exp_41_ram[3999] = 239;
    exp_41_ram[4000] = 147;
    exp_41_ram[4001] = 19;
    exp_41_ram[4002] = 183;
    exp_41_ram[4003] = 163;
    exp_41_ram[4004] = 239;
    exp_41_ram[4005] = 35;
    exp_41_ram[4006] = 111;
    exp_41_ram[4007] = 19;
    exp_41_ram[4008] = 147;
    exp_41_ram[4009] = 51;
    exp_41_ram[4010] = 19;
    exp_41_ram[4011] = 179;
    exp_41_ram[4012] = 99;
    exp_41_ram[4013] = 99;
    exp_41_ram[4014] = 19;
    exp_41_ram[4015] = 179;
    exp_41_ram[4016] = 19;
    exp_41_ram[4017] = 103;
    exp_41_ram[4018] = 227;
    exp_41_ram[4019] = 19;
    exp_41_ram[4020] = 179;
    exp_41_ram[4021] = 111;
    exp_41_ram[4022] = 128;
    exp_41_ram[4023] = 0;
    exp_41_ram[4024] = 0;
    exp_41_ram[4025] = 0;
    exp_41_ram[4026] = 0;
    exp_41_ram[4027] = 128;
    exp_41_ram[4028] = 136;
    exp_41_ram[4029] = 144;
    exp_41_ram[4030] = 152;
    exp_41_ram[4031] = 160;
    exp_41_ram[4032] = 168;
    exp_41_ram[4033] = 69;
    exp_41_ram[4034] = 76;
    exp_41_ram[4035] = 86;
    exp_41_ram[4036] = 79;
    exp_41_ram[4037] = 88;
    exp_41_ram[4038] = 65;
    exp_41_ram[4039] = 67;
    exp_41_ram[4040] = 65;
    exp_41_ram[4041] = 83;
    exp_41_ram[4042] = 88;
    exp_41_ram[4043] = 87;
    exp_41_ram[4044] = 81;
    exp_41_ram[4045] = 80;
    exp_41_ram[4046] = 79;
    exp_41_ram[4047] = 66;
    exp_41_ram[4048] = 74;
    exp_41_ram[4049] = 82;
    exp_41_ram[4050] = 90;
    exp_41_ram[4051] = 73;
    exp_41_ram[4052] = 75;
    exp_41_ram[4053] = 81;
    exp_41_ram[4054] = 69;
    exp_41_ram[4055] = 80;
    exp_41_ram[4056] = 89;
    exp_41_ram[4057] = 82;
    exp_41_ram[4058] = 78;
    exp_41_ram[4059] = 75;
    exp_41_ram[4060] = 87;
    exp_41_ram[4061] = 86;
    exp_41_ram[4062] = 71;
    exp_41_ram[4063] = 85;
    exp_41_ram[4064] = 78;
    exp_41_ram[4065] = 65;
    exp_41_ram[4066] = 81;
    exp_41_ram[4067] = 67;
    exp_41_ram[4068] = 69;
    exp_41_ram[4069] = 65;
    exp_41_ram[4070] = 86;
    exp_41_ram[4071] = 67;
    exp_41_ram[4072] = 79;
    exp_41_ram[4073] = 80;
    exp_41_ram[4074] = 71;
    exp_41_ram[4075] = 89;
    exp_41_ram[4076] = 81;
    exp_41_ram[4077] = 80;
    exp_41_ram[4078] = 79;
    exp_41_ram[4079] = 69;
    exp_41_ram[4080] = 67;
    exp_41_ram[4081] = 65;
    exp_41_ram[4082] = 70;
    exp_41_ram[4083] = 73;
    exp_41_ram[4084] = 69;
    exp_41_ram[4085] = 88;
    exp_41_ram[4086] = 84;
    exp_41_ram[4087] = 83;
    exp_41_ram[4088] = 72;
  end

  //Implement RAM port (Asynchronous)
  always@(posedge clk) begin
    if (exp_39) begin
      exp_41_ram[exp_35] <= exp_37;
    end
  end
  assign exp_41 = exp_41_ram[exp_36];


  //Additional RAM port (asynchronous)
  always@(posedge clk) begin
    if (exp_67) begin
        exp_41_ram[exp_63] <= exp_65;
    end
  end
  assign exp_69 = exp_41_ram[exp_64];
  assign exp_68 = exp_100;
  assign exp_100 = 1;
  assign exp_64 = exp_99;
  assign exp_99 = exp_16[31:2];
  assign exp_67 = exp_92;
  assign exp_63 = exp_91;
  assign exp_65 = exp_91;
  assign exp_40 = exp_135;
  assign exp_135 = 1;
  assign exp_36 = exp_134;
  assign exp_134 = exp_18[31:2];
  assign exp_39 = exp_109;
  assign exp_109 = exp_107 & exp_108;
  assign exp_107 = exp_22 & exp_23;
  assign exp_108 = exp_24[0:0];
  assign exp_35 = exp_105;
  assign exp_105 = exp_18[31:2];
  assign exp_37 = exp_106;
  assign exp_106 = exp_19[7:0];
  assign exp_126 = 1;

  reg [31:0] exp_160_reg;
  always@(*) begin
    case (exp_156)
      0:exp_160_reg <= exp_158;
      1:exp_160_reg <= exp_149;
      default:exp_160_reg <= exp_159;
    endcase
  end
  assign exp_160 = exp_160_reg;
  assign exp_159 = 0;
  assign exp_158 = 0;
  assign exp_149 = exp_187;

  reg [31:0] exp_187_reg;
  always@(*) begin
    case (exp_185)
      0:exp_187_reg <= exp_165;
      1:exp_187_reg <= exp_175;
      default:exp_187_reg <= exp_186;
    endcase
  end
  assign exp_187 = exp_187_reg;
  assign exp_185 = exp_147[2:2];
  assign exp_147 = exp_9;
  assign exp_186 = 0;

      reg [31:0] exp_165_reg = 0;
      always@(posedge clk) begin
        if (exp_164) begin
          exp_165_reg <= exp_172;
        end
      end
      assign exp_165 = exp_165_reg;
    
  reg [31:0] exp_172_reg;
  always@(*) begin
    case (exp_167)
      0:exp_172_reg <= exp_169;
      1:exp_172_reg <= exp_170;
      default:exp_172_reg <= exp_171;
    endcase
  end
  assign exp_172 = exp_172_reg;
  assign exp_167 = exp_165 == exp_166;
  assign exp_166 = 4294967295;
  assign exp_171 = 0;
  assign exp_169 = exp_165 + exp_168;
  assign exp_168 = 1;
  assign exp_170 = 0;
  assign exp_164 = 1;

      reg [31:0] exp_175_reg = 0;
      always@(posedge clk) begin
        if (exp_174) begin
          exp_175_reg <= exp_182;
        end
      end
      assign exp_175 = exp_175_reg;
    
  reg [31:0] exp_182_reg;
  always@(*) begin
    case (exp_177)
      0:exp_182_reg <= exp_179;
      1:exp_182_reg <= exp_180;
      default:exp_182_reg <= exp_181;
    endcase
  end
  assign exp_182 = exp_182_reg;
  assign exp_177 = exp_175 == exp_176;
  assign exp_176 = 4294967295;
  assign exp_181 = 0;
  assign exp_179 = exp_175 + exp_178;
  assign exp_178 = 1;
  assign exp_180 = 0;
  assign exp_174 = exp_167 & exp_173;
  assign exp_173 = 1;

  reg [31:0] exp_201_reg;
  always@(*) begin
    case (exp_197)
      0:exp_201_reg <= exp_199;
      1:exp_201_reg <= exp_190;
      default:exp_201_reg <= exp_200;
    endcase
  end
  assign exp_201 = exp_201_reg;
  assign exp_200 = 0;
  assign exp_199 = 0;
  assign exp_190 = exp_304;
  assign exp_304 = exp_218;

      reg [7:0] exp_218_reg = 0;
      always@(posedge clk) begin
        if (exp_217) begin
          exp_218_reg <= exp_264;
        end
      end
      assign exp_218 = exp_218_reg;
    
  reg [7:0] exp_264_reg;
  always@(*) begin
    case (exp_262)
      0:exp_264_reg <= exp_218;
      1:exp_264_reg <= exp_230;
      default:exp_264_reg <= exp_263;
    endcase
  end
  assign exp_264 = exp_264_reg;
  assign exp_262 = exp_261 & exp_228;
  assign exp_263 = 0;
  assign exp_230 = {exp_212, exp_229};  assign exp_229 = exp_218[7:1];
  assign exp_217 = 1;

  reg [31:0] exp_318_reg;
  always@(*) begin
    case (exp_314)
      0:exp_318_reg <= exp_316;
      1:exp_318_reg <= exp_307;
      default:exp_318_reg <= exp_317;
    endcase
  end
  assign exp_318 = exp_318_reg;
  assign exp_317 = 0;
  assign exp_316 = 0;
  assign exp_307 = exp_456;
  assign exp_456 = 0;

  reg [31:0] exp_470_reg;
  always@(*) begin
    case (exp_466)
      0:exp_470_reg <= exp_468;
      1:exp_470_reg <= exp_459;
      default:exp_470_reg <= exp_469;
    endcase
  end
  assign exp_470 = exp_470_reg;
  assign exp_469 = 0;
  assign exp_468 = 0;
  assign exp_459 = exp_476;
  assign exp_476 = 0;

  reg [31:0] exp_491_reg;
  always@(*) begin
    case (exp_487)
      0:exp_491_reg <= exp_489;
      1:exp_491_reg <= exp_480;
      default:exp_491_reg <= exp_490;
    endcase
  end
  assign exp_491 = exp_491_reg;
  assign exp_490 = 0;
  assign exp_489 = 0;
  assign exp_480 = exp_519;
  assign exp_519 = 0;
  assign exp_746 = exp_523[15:8];
  assign exp_747 = exp_523[23:16];
  assign exp_748 = exp_523[31:24];
  assign exp_760 = $signed(exp_759);
  assign exp_759 = exp_758 + exp_754;
  assign exp_758 = 0;

  reg [15:0] exp_754_reg;
  always@(*) begin
    case (exp_744)
      0:exp_754_reg <= exp_751;
      1:exp_754_reg <= exp_752;
      default:exp_754_reg <= exp_753;
    endcase
  end
  assign exp_754 = exp_754_reg;
  assign exp_753 = 0;
  assign exp_751 = exp_523[15:0];
  assign exp_752 = exp_523[31:16];
  assign exp_761 = 0;
  assign exp_762 = exp_750;
  assign exp_763 = exp_754;
  assign exp_764 = 0;
  assign exp_765 = 0;

  reg [31:0] exp_1124_reg;
  always@(*) begin
    case (exp_914)
      0:exp_1124_reg <= exp_1120;
      1:exp_1124_reg <= exp_1122;
      default:exp_1124_reg <= exp_1123;
    endcase
  end
  assign exp_1124 = exp_1124_reg;
  assign exp_1123 = 0;

  reg [31:0] exp_1120_reg;
  always@(*) begin
    case (exp_891)
      0:exp_1120_reg <= exp_1115;
      1:exp_1120_reg <= exp_1116;
      default:exp_1120_reg <= exp_1119;
    endcase
  end
  assign exp_1120 = exp_1120_reg;
  assign exp_891 = exp_890 & exp_888;
  assign exp_890 = exp_883 == exp_889;
  assign exp_889 = 0;
  assign exp_1119 = 0;
  assign exp_1115 = exp_1114[63:32];

  reg [63:0] exp_1114_reg;
  always@(*) begin
    case (exp_1111)
      0:exp_1114_reg <= exp_1110;
      1:exp_1114_reg <= exp_1112;
      default:exp_1114_reg <= exp_1113;
    endcase
  end
  assign exp_1114 = exp_1114_reg;

      reg [0:0] exp_1111_reg = 0;
      always@(posedge clk) begin
        if (exp_1096) begin
          exp_1111_reg <= exp_1094;
        end
      end
      assign exp_1111 = exp_1111_reg;
    
      reg [0:0] exp_1094_reg = 0;
      always@(posedge clk) begin
        if (exp_1073) begin
          exp_1094_reg <= exp_1071;
        end
      end
      assign exp_1094 = exp_1094_reg;
    
      reg [0:0] exp_1071_reg = 0;
      always@(posedge clk) begin
        if (exp_1053) begin
          exp_1071_reg <= exp_1068;
        end
      end
      assign exp_1071 = exp_1071_reg;
      assign exp_1068 = exp_1066 ^ exp_1067;
  assign exp_1066 = exp_1048 & exp_1031;
  assign exp_1048 = exp_1047 + exp_1046;
  assign exp_1047 = 0;
  assign exp_1046 = exp_1044[31:31];

      reg [31:0] exp_1044_reg = 0;
      always@(posedge clk) begin
        if (exp_1043) begin
          exp_1044_reg <= exp_661;
        end
      end
      assign exp_1044 = exp_1044_reg;
      assign exp_1043 = exp_1033 == exp_1042;
  assign exp_1042 = 0;
  assign exp_1031 = exp_1030 | exp_897;
  assign exp_1030 = exp_891 | exp_894;
  assign exp_894 = exp_893 & exp_888;
  assign exp_893 = exp_883 == exp_892;
  assign exp_892 = 1;
  assign exp_897 = exp_896 & exp_888;
  assign exp_896 = exp_883 == exp_895;
  assign exp_895 = 2;
  assign exp_1067 = exp_1051 & exp_1032;
  assign exp_1051 = exp_1050 + exp_1049;
  assign exp_1050 = 0;
  assign exp_1049 = exp_1045[31:31];

      reg [31:0] exp_1045_reg = 0;
      always@(posedge clk) begin
        if (exp_1043) begin
          exp_1045_reg <= exp_662;
        end
      end
      assign exp_1045 = exp_1045_reg;
      assign exp_1032 = exp_891 | exp_894;
  assign exp_1053 = exp_1033 == exp_1052;
  assign exp_1052 = 1;
  assign exp_1073 = exp_1033 == exp_1072;
  assign exp_1072 = 2;
  assign exp_1096 = exp_1033 == exp_1095;
  assign exp_1095 = 3;
  assign exp_1113 = 0;

      reg [63:0] exp_1110_reg = 0;
      always@(posedge clk) begin
        if (exp_1096) begin
          exp_1110_reg <= exp_1109;
        end
      end
      assign exp_1110 = exp_1110_reg;
      assign exp_1109 = exp_1105 + exp_1108;
  assign exp_1105 = exp_1101 + exp_1104;
  assign exp_1101 = exp_1097 + exp_1100;
  assign exp_1097 = exp_1090;

      reg [31:0] exp_1090_reg = 0;
      always@(posedge clk) begin
        if (exp_1073) begin
          exp_1090_reg <= exp_1077;
        end
      end
      assign exp_1090 = exp_1090_reg;
      assign exp_1077 = exp_1075 * exp_1076;
  assign exp_1075 = exp_1074;
  assign exp_1074 = exp_1069[15:0];

      reg [31:0] exp_1069_reg = 0;
      always@(posedge clk) begin
        if (exp_1053) begin
          exp_1069_reg <= exp_1059;
        end
      end
      assign exp_1069 = exp_1069_reg;
      assign exp_1059 = exp_1058 + exp_1057;
  assign exp_1058 = 0;

  reg [31:0] exp_1057_reg;
  always@(*) begin
    case (exp_1054)
      0:exp_1057_reg <= exp_1044;
      1:exp_1057_reg <= exp_1055;
      default:exp_1057_reg <= exp_1056;
    endcase
  end
  assign exp_1057 = exp_1057_reg;
  assign exp_1054 = exp_1048 & exp_1031;
  assign exp_1056 = 0;
  assign exp_1055 = -exp_1044;
  assign exp_1076 = exp_1070[15:0];

      reg [31:0] exp_1070_reg = 0;
      always@(posedge clk) begin
        if (exp_1053) begin
          exp_1070_reg <= exp_1065;
        end
      end
      assign exp_1070 = exp_1070_reg;
      assign exp_1065 = exp_1064 + exp_1063;
  assign exp_1064 = 0;

  reg [31:0] exp_1063_reg;
  always@(*) begin
    case (exp_1060)
      0:exp_1063_reg <= exp_1045;
      1:exp_1063_reg <= exp_1061;
      default:exp_1063_reg <= exp_1062;
    endcase
  end
  assign exp_1063 = exp_1063_reg;
  assign exp_1060 = exp_1051 & exp_1032;
  assign exp_1062 = 0;
  assign exp_1061 = -exp_1045;
  assign exp_1100 = exp_1098 << exp_1099;
  assign exp_1098 = exp_1091;

      reg [31:0] exp_1091_reg = 0;
      always@(posedge clk) begin
        if (exp_1073) begin
          exp_1091_reg <= exp_1081;
        end
      end
      assign exp_1091 = exp_1091_reg;
      assign exp_1081 = exp_1079 * exp_1080;
  assign exp_1079 = exp_1078;
  assign exp_1078 = exp_1069[15:0];
  assign exp_1080 = exp_1070[31:16];
  assign exp_1099 = 16;
  assign exp_1104 = exp_1102 << exp_1103;
  assign exp_1102 = exp_1092;

      reg [31:0] exp_1092_reg = 0;
      always@(posedge clk) begin
        if (exp_1073) begin
          exp_1092_reg <= exp_1085;
        end
      end
      assign exp_1092 = exp_1092_reg;
      assign exp_1085 = exp_1083 * exp_1084;
  assign exp_1083 = exp_1082;
  assign exp_1082 = exp_1069[31:16];
  assign exp_1084 = exp_1070[15:0];
  assign exp_1103 = 16;
  assign exp_1108 = exp_1106 << exp_1107;
  assign exp_1106 = exp_1093;

      reg [31:0] exp_1093_reg = 0;
      always@(posedge clk) begin
        if (exp_1073) begin
          exp_1093_reg <= exp_1089;
        end
      end
      assign exp_1093 = exp_1093_reg;
      assign exp_1089 = exp_1087 * exp_1088;
  assign exp_1087 = exp_1086;
  assign exp_1086 = exp_1069[31:16];
  assign exp_1088 = exp_1070[31:16];
  assign exp_1107 = 32;
  assign exp_1112 = -exp_1110;
  assign exp_1116 = exp_1114[31:0];

  reg [31:0] exp_1122_reg;
  always@(*) begin
    case (exp_915)
      0:exp_1122_reg <= exp_1025;
      1:exp_1122_reg <= exp_1026;
      default:exp_1122_reg <= exp_1121;
    endcase
  end
  assign exp_1122 = exp_1122_reg;
  assign exp_915 = exp_883[1:1];
  assign exp_1121 = 0;

      reg [31:0] exp_1025_reg = 0;
      always@(posedge clk) begin
        if (exp_934) begin
          exp_1025_reg <= exp_1019;
        end
      end
      assign exp_1025 = exp_1025_reg;
    
  reg [31:0] exp_1019_reg;
  always@(*) begin
    case (exp_1015)
      0:exp_1019_reg <= exp_1006;
      1:exp_1019_reg <= exp_1017;
      default:exp_1019_reg <= exp_1018;
    endcase
  end
  assign exp_1019 = exp_1019_reg;
  assign exp_1015 = exp_1014 & exp_917;
  assign exp_1014 = exp_963 == exp_1013;

      reg [31:0] exp_963_reg = 0;
      always@(posedge clk) begin
        if (exp_948) begin
          exp_963_reg <= exp_960;
        end
      end
      assign exp_963 = exp_963_reg;
      assign exp_960 = exp_959 + exp_958;
  assign exp_959 = 0;

  reg [31:0] exp_958_reg;
  always@(*) begin
    case (exp_955)
      0:exp_958_reg <= exp_940;
      1:exp_958_reg <= exp_956;
      default:exp_958_reg <= exp_957;
    endcase
  end
  assign exp_958 = exp_958_reg;
  assign exp_955 = exp_946 & exp_917;
  assign exp_946 = exp_945 + exp_944;
  assign exp_945 = 0;
  assign exp_944 = exp_940[31:31];

      reg [31:0] exp_940_reg = 0;
      always@(posedge clk) begin
        if (exp_938) begin
          exp_940_reg <= exp_662;
        end
      end
      assign exp_940 = exp_940_reg;
      assign exp_938 = exp_920 == exp_937;
  assign exp_937 = 0;
  assign exp_917 = ~exp_916;
  assign exp_916 = exp_883[0:0];
  assign exp_957 = 0;
  assign exp_956 = -exp_940;
  assign exp_948 = exp_920 == exp_947;
  assign exp_947 = 1;
  assign exp_1013 = 0;
  assign exp_1018 = 0;
  assign exp_1006 = exp_1005 + exp_1004;
  assign exp_1005 = 0;

  reg [31:0] exp_1004_reg;
  always@(*) begin
    case (exp_1001)
      0:exp_1004_reg <= exp_999;
      1:exp_1004_reg <= exp_1002;
      default:exp_1004_reg <= exp_1003;
    endcase
  end
  assign exp_1004 = exp_1004_reg;
  assign exp_1001 = exp_965 & exp_917;

      reg [0:0] exp_965_reg = 0;
      always@(posedge clk) begin
        if (exp_948) begin
          exp_965_reg <= exp_961;
        end
      end
      assign exp_965 = exp_965_reg;
      assign exp_961 = exp_943 ^ exp_946;
  assign exp_943 = exp_942 + exp_941;
  assign exp_942 = 0;
  assign exp_941 = exp_939[31:31];

      reg [31:0] exp_939_reg = 0;
      always@(posedge clk) begin
        if (exp_938) begin
          exp_939_reg <= exp_661;
        end
      end
      assign exp_939 = exp_939_reg;
      assign exp_1003 = 0;

      reg [31:0] exp_999_reg = 0;
      always@(posedge clk) begin
        if (exp_932) begin
          exp_999_reg <= exp_969;
        end
      end
      assign exp_999 = exp_999_reg;
    
      reg [31:0] exp_969_reg = 0;
      always@(posedge clk) begin
        if (exp_968) begin
          exp_969_reg <= exp_996;
        end
      end
      assign exp_969 = exp_969_reg;
    
  reg [31:0] exp_996_reg;
  always@(*) begin
    case (exp_930)
      0:exp_996_reg <= exp_988;
      1:exp_996_reg <= exp_994;
      default:exp_996_reg <= exp_995;
    endcase
  end
  assign exp_996 = exp_996_reg;
  assign exp_930 = exp_920 == exp_929;
  assign exp_929 = 2;
  assign exp_995 = 0;

  reg [31:0] exp_988_reg;
  always@(*) begin
    case (exp_978)
      0:exp_988_reg <= exp_982;
      1:exp_988_reg <= exp_986;
      default:exp_988_reg <= exp_987;
    endcase
  end
  assign exp_988 = exp_988_reg;
  assign exp_978 = ~exp_977;
  assign exp_977 = exp_976[32:32];
  assign exp_976 = exp_975 - exp_963;
  assign exp_975 = exp_974;
  assign exp_974 = {exp_972, exp_973};  assign exp_972 = exp_967[31:0];

      reg [31:0] exp_967_reg = 0;
      always@(posedge clk) begin
        if (exp_966) begin
          exp_967_reg <= exp_993;
        end
      end
      assign exp_967 = exp_967_reg;
    
  reg [32:0] exp_993_reg;
  always@(*) begin
    case (exp_930)
      0:exp_993_reg <= exp_980;
      1:exp_993_reg <= exp_991;
      default:exp_993_reg <= exp_992;
    endcase
  end
  assign exp_993 = exp_993_reg;
  assign exp_992 = 0;

  reg [32:0] exp_980_reg;
  always@(*) begin
    case (exp_978)
      0:exp_980_reg <= exp_974;
      1:exp_980_reg <= exp_976;
      default:exp_980_reg <= exp_979;
    endcase
  end
  assign exp_980 = exp_980_reg;
  assign exp_979 = 0;
  assign exp_991 = 0;
  assign exp_966 = 1;
  assign exp_973 = exp_971[31:31];

      reg [31:0] exp_971_reg = 0;
      always@(posedge clk) begin
        if (exp_970) begin
          exp_971_reg <= exp_998;
        end
      end
      assign exp_971 = exp_971_reg;
    
  reg [31:0] exp_998_reg;
  always@(*) begin
    case (exp_930)
      0:exp_998_reg <= exp_990;
      1:exp_998_reg <= exp_962;
      default:exp_998_reg <= exp_997;
    endcase
  end
  assign exp_998 = exp_998_reg;
  assign exp_997 = 0;
  assign exp_990 = exp_971 << exp_989;
  assign exp_989 = 1;

      reg [31:0] exp_962_reg = 0;
      always@(posedge clk) begin
        if (exp_948) begin
          exp_962_reg <= exp_954;
        end
      end
      assign exp_962 = exp_962_reg;
      assign exp_954 = exp_953 + exp_952;
  assign exp_953 = 0;

  reg [31:0] exp_952_reg;
  always@(*) begin
    case (exp_949)
      0:exp_952_reg <= exp_939;
      1:exp_952_reg <= exp_950;
      default:exp_952_reg <= exp_951;
    endcase
  end
  assign exp_952 = exp_952_reg;
  assign exp_949 = exp_943 & exp_917;
  assign exp_951 = 0;
  assign exp_950 = -exp_939;
  assign exp_970 = 1;
  assign exp_987 = 0;
  assign exp_982 = exp_969 << exp_981;
  assign exp_981 = 1;
  assign exp_986 = exp_984 | exp_985;
  assign exp_984 = exp_969 << exp_983;
  assign exp_983 = 1;
  assign exp_985 = 1;
  assign exp_994 = 0;
  assign exp_968 = 1;
  assign exp_932 = exp_920 == exp_931;
  assign exp_931 = 35;
  assign exp_1002 = -exp_999;
  assign exp_1017 = $signed(exp_1016);
  assign exp_1016 = -1;
  assign exp_934 = exp_920 == exp_933;
  assign exp_933 = 36;

      reg [31:0] exp_1026_reg = 0;
      always@(posedge clk) begin
        if (exp_934) begin
          exp_1026_reg <= exp_1024;
        end
      end
      assign exp_1026 = exp_1026_reg;
    
  reg [31:0] exp_1024_reg;
  always@(*) begin
    case (exp_1022)
      0:exp_1024_reg <= exp_1012;
      1:exp_1024_reg <= exp_939;
      default:exp_1024_reg <= exp_1023;
    endcase
  end
  assign exp_1024 = exp_1024_reg;
  assign exp_1022 = exp_1021 & exp_917;
  assign exp_1021 = exp_963 == exp_1020;
  assign exp_1020 = 0;
  assign exp_1023 = 0;
  assign exp_1012 = exp_1011 + exp_1010;
  assign exp_1011 = 0;

  reg [31:0] exp_1010_reg;
  always@(*) begin
    case (exp_1007)
      0:exp_1010_reg <= exp_1000;
      1:exp_1010_reg <= exp_1008;
      default:exp_1010_reg <= exp_1009;
    endcase
  end
  assign exp_1010 = exp_1010_reg;
  assign exp_1007 = exp_964 & exp_917;

      reg [0:0] exp_964_reg = 0;
      always@(posedge clk) begin
        if (exp_948) begin
          exp_964_reg <= exp_943;
        end
      end
      assign exp_964 = exp_964_reg;
      assign exp_1009 = 0;

      reg [31:0] exp_1000_reg = 0;
      always@(posedge clk) begin
        if (exp_932) begin
          exp_1000_reg <= exp_967;
        end
      end
      assign exp_1000 = exp_1000_reg;
      assign exp_1008 = -exp_1000;
  assign exp_595 = $signed(exp_594);
  assign exp_594 = 0;
  assign exp_824 = exp_659 != exp_660;
  assign exp_837 = 0;
  assign exp_838 = 0;
  assign exp_825 = $signed(exp_659) < $signed(exp_660);
  assign exp_826 = $signed(exp_659) >= $signed(exp_660);
  assign exp_831 = exp_828 < exp_830;
  assign exp_828 = exp_827 + exp_659;
  assign exp_827 = 0;
  assign exp_830 = exp_829 + exp_660;
  assign exp_829 = 0;
  assign exp_836 = exp_833 >= exp_835;
  assign exp_833 = exp_832 + exp_659;
  assign exp_832 = 0;
  assign exp_835 = exp_834 + exp_660;
  assign exp_834 = 0;
  assign exp_1151 = 0;
  assign exp_1150 = exp_549 + exp_1149;
  assign exp_1149 = 4;

  reg [32:0] exp_881_reg;
  always@(*) begin
    case (exp_682)
      0:exp_881_reg <= exp_871;
      1:exp_881_reg <= exp_879;
      default:exp_881_reg <= exp_880;
    endcase
  end
  assign exp_881 = exp_881_reg;
  assign exp_880 = 0;
  assign exp_871 = exp_870 + exp_668;

  reg [31:0] exp_870_reg;
  always@(*) begin
    case (exp_680)
      0:exp_870_reg <= exp_856;
      1:exp_870_reg <= exp_868;
      default:exp_870_reg <= exp_869;
    endcase
  end
  assign exp_870 = exp_870_reg;
  assign exp_869 = 0;
  assign exp_856 = $signed(exp_855);
  assign exp_855 = exp_854 + exp_853;
  assign exp_854 = 0;
  assign exp_853 = {exp_852, exp_849};  assign exp_852 = {exp_851, exp_848};  assign exp_851 = {exp_850, exp_847};  assign exp_850 = {exp_845, exp_846};  assign exp_845 = exp_667[31:31];
  assign exp_846 = exp_667[7:7];
  assign exp_847 = exp_667[30:25];
  assign exp_848 = exp_667[11:8];
  assign exp_849 = 0;
  assign exp_868 = $signed(exp_867);
  assign exp_867 = exp_866 + exp_865;
  assign exp_866 = 0;
  assign exp_865 = {exp_864, exp_861};  assign exp_864 = {exp_863, exp_860};  assign exp_863 = {exp_862, exp_859};  assign exp_862 = {exp_857, exp_858};  assign exp_857 = exp_667[31:31];
  assign exp_858 = exp_667[19:12];
  assign exp_859 = exp_667[20:20];
  assign exp_860 = exp_667[30:21];
  assign exp_861 = 0;

      reg [31:0] exp_668_reg = 0;
      always@(posedge clk) begin
        if (exp_658) begin
          exp_668_reg <= exp_551;
        end
      end
      assign exp_668 = exp_668_reg;
      assign exp_879 = exp_878 & exp_877;
  assign exp_878 = $signed(exp_876);
  assign exp_876 = exp_659 + exp_875;
  assign exp_875 = $signed(exp_874);
  assign exp_874 = exp_873 + exp_872;
  assign exp_873 = 0;
  assign exp_872 = exp_667[31:20];
  assign exp_877 = 4294967294;
  assign exp_548 = exp_541 & exp_539;
  assign exp_88 = exp_92;
  assign exp_84 = exp_91;
  assign exp_86 = exp_91;
  assign exp_17 = exp_550;
  assign exp_683 = 3;
  assign exp_530 = ~exp_528;
  assign exp_310 = exp_12;
  assign exp_382 = 0;
  assign exp_337 = 433;
  assign exp_343 = 433;
  assign exp_349 = exp_335 - exp_348;
  assign exp_348 = 1;
  assign exp_355 = 433;
  assign exp_363 = exp_335 - exp_362;
  assign exp_362 = 1;
  assign exp_369 = exp_335 - exp_368;
  assign exp_368 = 1;
  assign exp_334 = 1;
  assign exp_364 = 0;
  assign exp_446 = 0;

  reg [2:0] exp_432_reg;
  always@(*) begin
    case (exp_430)
      0:exp_432_reg <= exp_396;
      1:exp_432_reg <= exp_359;
      default:exp_432_reg <= exp_431;
    endcase
  end
  assign exp_432 = exp_432_reg;
  assign exp_430 = exp_426 & exp_357;
  assign exp_357 = exp_327 == exp_356;

      reg [2:0] exp_327_reg = 0;
      always@(posedge clk) begin
        if (exp_326) begin
          exp_327_reg <= exp_436;
        end
      end
      assign exp_327 = exp_327_reg;
    
  reg [2:0] exp_436_reg;
  always@(*) begin
    case (exp_434)
      0:exp_436_reg <= exp_402;
      1:exp_436_reg <= exp_361;
      default:exp_436_reg <= exp_435;
    endcase
  end
  assign exp_436 = exp_436_reg;
  assign exp_434 = exp_426 & exp_433;
  assign exp_433 = ~exp_357;
  assign exp_435 = 0;

  reg [2:0] exp_402_reg;
  always@(*) begin
    case (exp_400)
      0:exp_402_reg <= exp_327;
      1:exp_402_reg <= exp_344;
      default:exp_402_reg <= exp_401;
    endcase
  end
  assign exp_402 = exp_402_reg;
  assign exp_400 = exp_393 & exp_341;
  assign exp_401 = 0;
  assign exp_344 = 0;
  assign exp_361 = exp_327 + exp_360;
  assign exp_360 = 1;
  assign exp_326 = 1;
  assign exp_356 = 7;
  assign exp_431 = 0;

  reg [2:0] exp_396_reg;
  always@(*) begin
    case (exp_394)
      0:exp_396_reg <= exp_380;
      1:exp_396_reg <= exp_342;
      default:exp_396_reg <= exp_395;
    endcase
  end
  assign exp_396 = exp_396_reg;
  assign exp_394 = exp_393 & exp_341;
  assign exp_395 = 0;

  reg [2:0] exp_380_reg;
  always@(*) begin
    case (exp_378)
      0:exp_380_reg <= exp_325;
      1:exp_380_reg <= exp_336;
      default:exp_380_reg <= exp_379;
    endcase
  end
  assign exp_380 = exp_380_reg;
  assign exp_378 = exp_374 & exp_323;
  assign exp_379 = 0;
  assign exp_336 = 1;
  assign exp_342 = 2;
  assign exp_359 = 4;
  assign exp_366 = 0;
  assign exp_324 = 1;
  assign exp_414 = 2;
  assign exp_428 = 0;

  reg [0:0] exp_422_reg;
  always@(*) begin
    case (exp_420)
      0:exp_422_reg <= exp_405;
      1:exp_422_reg <= exp_354;
      default:exp_422_reg <= exp_421;
    endcase
  end
  assign exp_422 = exp_422_reg;
  assign exp_420 = exp_416 & exp_351;
  assign exp_421 = 0;

  reg [0:0] exp_405_reg;
  always@(*) begin
    case (exp_403)
      0:exp_405_reg <= exp_389;
      1:exp_405_reg <= exp_345;
      default:exp_405_reg <= exp_404;
    endcase
  end
  assign exp_405 = exp_405_reg;
  assign exp_403 = exp_393 & exp_341;
  assign exp_404 = 0;

  reg [0:0] exp_389_reg;
  always@(*) begin
    case (exp_387)
      0:exp_389_reg <= exp_333;
      1:exp_389_reg <= exp_339;
      default:exp_389_reg <= exp_388;
    endcase
  end
  assign exp_389 = exp_389_reg;
  assign exp_387 = exp_374 & exp_323;
  assign exp_388 = 0;
  assign exp_339 = 0;
  assign exp_345 = exp_329[0:0];

      reg [7:0] exp_329_reg = 0;
      always@(posedge clk) begin
        if (exp_328) begin
          exp_329_reg <= exp_419;
        end
      end
      assign exp_329 = exp_329_reg;
    
  reg [7:0] exp_419_reg;
  always@(*) begin
    case (exp_417)
      0:exp_419_reg <= exp_408;
      1:exp_419_reg <= exp_353;
      default:exp_419_reg <= exp_418;
    endcase
  end
  assign exp_419 = exp_419_reg;
  assign exp_417 = exp_416 & exp_351;
  assign exp_418 = 0;

  reg [7:0] exp_408_reg;
  always@(*) begin
    case (exp_406)
      0:exp_408_reg <= exp_377;
      1:exp_408_reg <= exp_347;
      default:exp_408_reg <= exp_407;
    endcase
  end
  assign exp_408 = exp_408_reg;
  assign exp_406 = exp_393 & exp_341;
  assign exp_407 = 0;

  reg [7:0] exp_377_reg;
  always@(*) begin
    case (exp_375)
      0:exp_377_reg <= exp_329;
      1:exp_377_reg <= exp_322;
      default:exp_377_reg <= exp_376;
    endcase
  end
  assign exp_377 = exp_377_reg;
  assign exp_375 = exp_374 & exp_323;
  assign exp_376 = 0;
  assign exp_322 = exp_306[7:0];
  assign exp_306 = exp_10;
  assign exp_347 = exp_329 >> exp_346;
  assign exp_346 = 1;
  assign exp_353 = exp_329 >> exp_352;
  assign exp_352 = 1;
  assign exp_328 = 1;
  assign exp_354 = exp_329[0:0];
  assign exp_358 = 1;
  assign exp_332 = 1;

      reg [31:0] exp_475_reg = 0;
      always@(posedge clk) begin
        if (exp_474) begin
          exp_475_reg <= exp_458;
        end
      end
      assign exp_475 = exp_475_reg;
      assign exp_458 = exp_10;
  assign exp_474 = exp_461 & exp_462;
  assign exp_461 = exp_467;
  assign exp_467 = exp_11 & exp_466;
  assign exp_462 = exp_12;
  assign exp_518 = exp_517 > exp_507;

      reg [10:0] exp_517_reg = 0;
      always@(posedge clk) begin
        if (exp_495) begin
          exp_517_reg <= exp_479;
        end
      end
      assign exp_517 = exp_517_reg;
      assign exp_479 = exp_10;
  assign exp_495 = exp_482 & exp_483;
  assign exp_482 = exp_488;
  assign exp_488 = exp_11 & exp_487;
  assign exp_483 = exp_12;

      reg [9:0] exp_507_reg = 0;
      always@(posedge clk) begin
        if (exp_506) begin
          exp_507_reg <= exp_514;
        end
      end
      assign exp_507 = exp_507_reg;
    
  reg [9:0] exp_514_reg;
  always@(*) begin
    case (exp_509)
      0:exp_514_reg <= exp_511;
      1:exp_514_reg <= exp_512;
      default:exp_514_reg <= exp_513;
    endcase
  end
  assign exp_514 = exp_514_reg;
  assign exp_509 = exp_507 == exp_508;
  assign exp_508 = 1023;
  assign exp_513 = 0;
  assign exp_511 = exp_507 + exp_510;
  assign exp_510 = 1;
  assign exp_512 = 0;
  assign exp_506 = exp_499 & exp_505;
  assign exp_499 = exp_497 == exp_498;

      reg [1:0] exp_497_reg = 0;
      always@(posedge clk) begin
        if (exp_496) begin
          exp_497_reg <= exp_504;
        end
      end
      assign exp_497 = exp_497_reg;
    
  reg [1:0] exp_504_reg;
  always@(*) begin
    case (exp_499)
      0:exp_504_reg <= exp_501;
      1:exp_504_reg <= exp_502;
      default:exp_504_reg <= exp_503;
    endcase
  end
  assign exp_504 = exp_504_reg;
  assign exp_503 = 0;
  assign exp_501 = exp_497 + exp_500;
  assign exp_500 = 1;
  assign exp_502 = 0;
  assign exp_496 = 1;
  assign exp_498 = 4;
  assign exp_505 = 1;
  assign stdout_tx = exp_333;
  assign leds_out = exp_475;
  assign pwm_pwm_out = exp_518;

endmodule